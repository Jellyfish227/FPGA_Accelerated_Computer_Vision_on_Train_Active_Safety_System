/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 430784)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnCLakmLX1fY5c7qjlPfHMwwhbJ3U6Jewr1Idxd+R9GBSPuYH/CstJgmT
7ETmyswtbH9av7VRbTASgEDQAcv/cn2QfhiuH1DAz4FQk0fX1cN/fCHukNpMY3yqdxzjYtVi+jyK
667FD5U1jees0xujNZKqCxSoacVDeF1rVBdFO9CdrFGwB3JeCuKM+auhCf8YIwIt/jo66+kwjN28
WBb69J6CGhOonL+jJkBquBRtQzBvMl0KygZQvhnO7ukmdub1F06lS6oaZUnggserxWm4RdzPozzl
NsDcjUjoU4BmmfN6rzCiNdPTFRnKKvG+y3b4DIhjhe3qxnzQaGNf3duXxEwHWgemeRyXGlydbtDT
x1/qRynDJs/cdMlThEekez9PVW2mWV37lz5BlkWs/RmkhBp/q5ZH/WDaTS5pP9/sR8ZrKpNyrQrr
Vr57SjJqoBSJ8Br+PDL4E3gD4MidwsARpcTm9FbS7rMnPZ6ZnFkloYXpsAIvCsCzT7fbLJlbI8qm
6j3IiNQ2/VIBelGxUl0ZyCHGSNkYoCeVFvsI9rq2kIEqtPP9U+JhGzcFjmiFlojXqI9+BB3uYEjx
6b95FfWnGpJ/wRegpdz/BSuaXn3JIihClIt/j0Qll5NgaK6ivXr8jma7u3bmh7Kplv459Bfki+m+
EjJ+EX4ONMpI/olXDM2uSGByJnP60CMfiBG11nkGJJYUw2kl57cQ9bWDXtaWmbduXaZbuC5BwxG7
DxvEjC2G0r65f22GiCleDMngu/RKEKa30t4w8cmiDXEK1PIIdwr4388dNPnDeRUt/kPMH8ewctSL
Ugdyk0te8gMkAH3d4OCONNvMmPqJGb5GBw2cl12N7TFsshcq2JXWFsskWWkR3/FYVBgRiLPvkHIZ
EodQCDmvrjd3mBU9BGI5duroTHLaQarVE+WzJOfBkricHguyJ7kDIKloxc2wpJODmuUc+93zTZzK
2HBn7Pvnb8t3I6tIASmGep+TD2KmkkWICaorlrZmYAMuk3voA5dT8Ca3GYoF47kSuSd0LzPxNVhe
sKQ368FYtlwaKlcfrgnKRtbVwFxYkw2jOh0D+eoMbgXGUQr36Mt6wz+SM9TLQRxmqBi9oZz5LP0C
2gTY2eq29vHeM05HuL3JZZKtEYptsZrzko3sviTmFWanuZDdP5fogNCIS31GzQfZwfsOsfjomZCQ
BcTCHTLVxKTdCrv2W1o7Rbau7cb9DvTxTxTZNo9mNGr0njzcUBqM7QtzilRYe23MbyfPn0QvCGgH
mh+bht354+9ZwrCrbP9mmXNwJCU2DV4vpU/E/sxQgYxqEnyJnAkJwdGwDP73c9RgKyvI1mcuGzGg
jNW306hxdPbE7H5bGlP/WuUzUN6nVnWsnp2Gf2GPGWoa+/sWuEd8ErKNEbo61xlV8tXg8aQXn7aH
CJSWkWv9UrwFujX3UoMjSE90OE5ewr4/kUuiDysUdWdlhZrKKxnAPDtO669DVHGz4KGtHjh76X70
Td0j9muziw95eQDyNs/UoxQYnTHaTydq0BywDbXqqQbnMlzC/RxE04IuY5NRUqmoksi/aJ8447bG
91M+U/qyRF8O9a1guFY3tImDeb4dtoxaXmUiT6qlkTD38n+Ik/D4wpp1mp7NOeZDBraKq+kiIQiQ
dVAp8yOjhgbH4AD+2wC9XN+b0fZ0Jhhk+qaxaQ5qCXtDlmFIqEHl2RYFUC7Qo7svG4xdlD8NiSke
q+cpJ0HseE72TDTfqPM+3z9XINOAjh/Gh4CJtvc8j4tXrZR/tz20CEHZWh82YoR8uKZYVIWxkxum
HfM0w1jAg9ZjchaY+Ic+8DsSqpPsWSmLQWvAXMs83YWA7AnH4wSBzD0oKiGvIQ3qPqcEoICRwh7R
zCYnE8tp88l/uqLPkHlW3Bz9ae8Eo+EN8yGMWnJ1Vhb1VT5wyhYbLKBZ8TBT62gMA10Uo9k9ta9/
b3qySONrR7WpHXKhB5+bLAfQ/o4wDl9VjyhuMHieDYSjJWDfiOt2ZhYK/kXhV5bLo2Sxnb13KS7l
8CI5S+sxCHTxaJHzs69tYFMomKbSCLU+7/hEjyZw1ceZHZ6jf5HXUeJXVu4707i7BUVzfNX/yvN3
tHHJAs5vU7egTDkUsOsfjlCDhebWutau39knVMqPu1thBINA2uedYGKYBE5ScdChwaQ4Quq+IpyO
oMSW7RJHeOdlSOa04FxaIBpsWH4l1WEol+fCFnZJvbSFvZn7zkI1aamKmSyBXsxBQXu6EEuQU7ah
fY6B2ceoBcqjREMm3AHcRPPQwWdFi5B9CbTTLLw6h9EF93Zqe/XLhfMiqxs6oNGHR0FsM8pm6t5T
FfCLxuMRWxA43mkG0lDky8raOBvah7wj+biEXpb+tqahfHWBlP4FEv9Qef4Cy6oVxI/OP+PCxMkH
zTaEpdwrWrYiAxJkC6xckCTfz6TSff0F3UiXuuNjnvO4Ry3KZz0aCZC87royqymHT2JiQgLNulVS
4oAxpsMjghccweF2+tS1MxBcl1EfBTz6NB1L/iCm2zrpAXibqL2oamDGGg2gpJ0Sp9y/u98XdUT7
zwyUXew3Gm2QGPKgyvn/j88DNzbvZ8h+rzwi+Nw55k5bp25P6DAjTRogTmzsbZQPtcbPrI+X9rwQ
50bfd8KSaD6KK7ztc6nZQyM9tH9NsGbjWCqtNISpElT9sIo0FztAHHspTGehAAdvNf9aumyr6Ceb
I0f/nAasPUfu7678FIzwfmefDZ3eyeKatZCXav+MydQLUWGMAZ0mI3bSj4+ReLQZvax0K8qeiN9c
0POTbaF1AcQLSgwStHUvbB5auj+WjSriW5N29VnmllJJl4vnQH1AvwwXS6q5mPiRegVJxUvy4r6I
JETjbXUib9/Anr6w25emxwTYKY6vMcHOE9VNBV/u3usf1PR6ZI0/BtMZjwAjoVK4EdXmscWh+6H3
fC3zMREd2w5yBaM1PGeMBo4costuOpL9EL+tn5HGx/VCNM9K9ToXqCzScVt5J9lkwfbVOAN0KRLb
5pxRyxwlNKatN5GvQZCDct8NRC4sx5uqQKKFo1/5D598fnqWv8gmW9DpbJAW6AxUBCEP8Gzr1drl
hjz7vL8F3L1d6TRXuvLDYt/sVuR+mxmkfaWpBqXssvpAE0XCkz41T7pyIV2DoLYJNx+y+roVnXlF
lddZI2f1Wrsxz11U9bU0OoXtEZXThGCv//lkthc5DHaLLfZlx1NG+zWjpJsGqtu2H3gmaiLG369h
qXYFipdRwvgf0ODiQo3wYOldjU8bmyBTWXFkM7G/SxR7s5CH8W2YAr+iSBeMajF6uf+LC0yEqxq/
0K8JP4xbhETcVUqDNXLYKZk6wrLxaCa6ymBOA6Cwb1X/Qk6O8mwNFEJ9LmNBPrJ19uy3cxI3bgRU
o3l/1Hiz642osMPWx6rvViUfX8beBNAUc1prDfh5mc2yqoi18iHr4IG8PDwl6cBXzzX+hOTs+Q8G
0y6MbeYYV7/qTmAueHopl8f2Y2T1VNdScSKLUvlsJcHifILxWbPcEk+GsVhDnz1RRj4E/4UfLNwJ
lUCPZYXa20bvLl575pt2tj1kLElV0DyqN+Rfslf2qQTL6Vm55LRdYxysnn41zbh2P4F1Xj1C3lRU
LXgmBgxoh6+42FMbuAiBHAyVe1Pe3hS0ETw4LgNM1gcwMYedzwJmjjsEffetPrLX8JWiROQdhlSU
fp6v4/1EH8EjWV8Ik9Q/V2+Z6PxAwY2XwdIrWV7wPJvrXw06VOistLnq8Uc0sjBXrE0qhPsLmR4L
GOmkKckakxqZW9MBJueA4H6CV5TpViZ/BaE/8Fd6tuARBI65qEe/JcuC/7NFAQbXy+yLpN6t5W2P
sy5aLoxM7wyobvPgLrQBD9pQmPCdcnp8AwTvHx4PkwZ2itliNjukvYx7auT0QyrBbyFe4Pms3KWn
NgYn8vGIiZKOhtNy62UlfggUiZJhAtM2aoJUAtnRuvIzqFYApJb1wUiw8DRhuZ0aziW4HK96Tt4b
bP5jIdyU5GGUgdbI65ELYxzubspEfZlW7kGahoOCH7j3J2T970aNLHQgyWBaelNwPx8BwgU+UJ2B
1W4Yjma3VAmhAkMyS2AZ6R39PgnVD8k82fnQou7nZNegg0LUh5YwXYmsy8cLzblP/ylbDHD1Vlkw
6YNo5q44u9vI9eGedTkooZKxSW9x81ZPtX7PyMpdN4o9XnbQ9rHsMunZFibVWxLNwxP7HXRmXhoV
3bn09E+Peb+ypaAnWpRQ7uItRKqiEW/QVBf5JKKC9CHMLYlT2b1D9cM5LE6pqv0LFS4bMrHcyHnR
dZb0S8+N9HVn+mZGaz6msV/xOZz5Rvz3rLJ2ZlKOgT4aK/Nz5O1KFSJqFhJi0POjc1oN30rHDBYb
/tmTYN/AU0qmJF3yxY2wD6wnCx6tlK+DV3eS01LZkNCuok+/xrB6EBo7OhBwf5gMM4m2jD2Ec8yH
5Xo5zrbNcvlvR7g8I2CQepE4sxcfcVjtb43MSxjAI4rARTZDRx3XyNuU9M18orRB8Um33YcI67Sg
cVFqW/gr4E/2uB0VoHq8smlu3bevQ1/2VRzxMv7wd2ETzHLWuVZ6GgqZhq4zWii8c8KqkA+/95G/
9ofKGqqqk7BmO8N66fKbUKucBCn/cN4TEFJDHy7qUnTiz1b50Da7w/yIN3TqNg3o3Uchwh7gE8ri
yEqBc97b0nw/QZpz3xqenLlPaOMmWb99vX7YCd+IvQNBgnZQGZGwzn5fjQ0Fb1dwJWKDan1eEIUD
NeD1RHvyOb1BKVl2dL0y9LnAeUNSp4dQb/J3PF46GaM6EVDPv3pYeq68g5jwdAzRHyGw6c8HtGi4
ah+OdJNXGjj7nFPn7ROS1nxqfi1Thg6L2sucemM5pnVXPXA0YOoouvFyqIWLG4DdvM6fGvFHTbR2
Gb36LyFUR7LpLzdKlzzul1SRBt99hAcgsZqICGkjAYg+kucsflbL9qLb7a84QZZBG3ub/sR3bSLe
fsHHecO77wyadyZK5cyFmXPaMOJX/LG7H+AQdUX7oC9xuKvc74Q7xszfmOTQwYJmBL+bK8IFOt+u
vLprjKjyG/C5zh2oefAwJFUU5f4yPeSsE9Wvo+w7OboCxEk/l/8kBEOYsmWGcpXBgfAm5peZkcwk
zf2pRP37GhOgLxzQx9Qv8KWT77PSWFo8zPrIO7kgvFeUruZph8Kz7CQzwspTFt3ky+OdcO6FdpRH
+EI4bu+YAaJFEZn0qkMCL4qIBjr/wywOFt/+uztOmrdUbBGB4VfTe5+jukbXLDzMPzq0OTdqKUuE
3kgtC13OLbOnd+oaphTo14fHzmQ/z3mUpn0DGPQd4Y5rf9HH3g0B8ZnCy0LwOyxegwm9btMHmRpI
CYnb8ksvbcnV0EMgzCsa2BZqEmV4BsoLpPCWifeciS8UV57Y4rEwrMW5yGojEW3sV3QAd78Bhop8
WMcF9bmSj0QFL0Y360WrN+Ait6tjM+jnvLmIUp2Wx+LwGR4eFkhIeEQb5234xclZkksnUatvWfeQ
UQ2UdviYdFToOvGDoVcH8QlrXYWnyd1qjoKc30YdzGLTiLALgHnC3S93Fa5uPA2EokIm5p1zc1I7
yJ88TMOgbWcL42HCIeHKWwxJH5Gi0a1DXTIDtNs8rftd0pS5Gx58LVqLmHfzhJBcebb0MYSt4qP1
gwjVGLSn8l/awf+3Nt5dDP+Jz5FUqa1ixlu+MTaBxkW+jNjj1eF8GHpwV3Bak6uaF/+5dWymVXWS
h+KASYMmY+pkDpsm8GvZL8G7m8eY1ZzwsnfTYdM8TzXOQHkwXilS2CPYD+4oWF/ttxMNsuQPrZ5L
H1NqU0U9sWG41sozdsf7Ox+gS3+0CpWUrdzeXkjTR/HtC2urbsS9+0Ik6KZcKr6EDCwMarAOfZoo
qAHKitiTrXYN1AEbWuFFQ4vznwhHv9IktoCiA+rsejA8U+G1W+gHEwniZUyFhg05czCBk7y0k5i2
W9ba3qVYTV+sEPFoz1JgcDdx4EJ6kFs92kbTjYbKk3V8zaMEldsDJp9FxzUlNODyO6GPs/FoNbPy
Y/WhUnehv7GUbjtCV0TIJbCF0hSAgpiAN0lmU2G+lDqeIyMLT2G6kXiTZF4edNI01ZlCDEFUEKLO
FWn8PeWhc0awk3ckU4knRuBoHSD5cYI7Z0Qg7R8R4Gyhb1izy3Qy7PcNLYqOamh+DyJPMBuOBdPo
18UbA5YhgY735tm5hiO+9AcWfVYhU18DnL6dY1TnyX5Key4pwWFXnMUkdyeU7SW1QCUl3ffNd7G5
iCAwBtwgJsXdPPJylIKCpdUg1TSHKwT+ytal0/xrvgxnMYQwXsdHeEI1IdtvJQ30V7O4XAuwU/4k
NlkpoRKiC/wtUJGythNTEfV53H8cQLH0zP4aFWs1MjmxgEn0iS3HaFL1kVZRzKq7x6f8ozpk/OS1
v3X6t/P9snaEXX5862ggkQIL399N5zUS/kJA6a4fCYUIFANUUb+oWzxyx/Vilr/DFqMPVXIjPn/D
yRhifUduIcsiuiYJNjTOk/iH/pj3iCVgZgPj4FQ4JuM77LGw4end5hKK+1hb1tlxE9XX3+xE8/zW
pCEwave2STP/rDZvpELOG4XXShZG+5HSm2jvUX6CIWmgEpBDxZgakKcfcERX/Zn0EUXz8NTyAlad
zPtB4CnHSU4fpcga/s4Xh994HiCQ3NNbS52p1WPY1vDc/DBo9YFolDXJCAf2NuJw0SdY3+2ktDcH
ES/CQ5SL2r14+3w7GYrw/hWRzELKl9VX3sqFpgwDVbxiAxIOlwGyvmdPrLCw5gYme8F2QszJrnye
aq+6nXfwKB8EV+X+eGySN6oZM8HJ3XXw58KwwjcmzwVt6H19+sy+YLGBUuxjl7zf35jL83cXwxST
sRtA2/XFgwiV4fT3hF5oLuPZL9k2OGw5te09IwZe0sCht/iooOoorIdn7jkdw+9mhAwgQENoFgxu
HgeI1DN39oO7jtGGgharrSfNKNjKzx/8EfFwO7C0+nulgHoNS30E/m8iPg97xebKuzDZf9FskkN4
K5po1UI3OjmmmLyj/Fu8hbqPYIEFwQf5MmqjEOI4i8KpOC3vTI43m84WC58ZTMX1Pl1LZbBFTwPu
+Yn/ckjz9qsdijm5cLM70Zol9UVs/5AWkoTaoN6lZWybz5n+Su9GOkvAJYRtw/uv0m/BjcnoIMtW
EZxn+I+DB6+pZJTSgl2B7PZmH2Uuua1q/QZE2ZMVGkWMmOSJkVCEpqmk9k/3LRUK0rcTtYXGnUFG
tJuSHfqQr9b3Ckv+XJbMkPVtdH5WS1fO0hfsHkbkRU8Bxrk2JhjL9sCyj/ot06XhCbl9mHxJUPE1
8P5DIqcVhb+1/ZiNmE4wJDvwig/vNqjk29xREqUt1noC1yUUn3rOj6nIQX1fPWTCweMES/SMzgii
PxCTjDQprwMFNfMO+wJaAR5Us8AFdBJK8wM9WaGgyhSrNqX40Q88PgxUN+zrStRBRJtaZS9mCUvv
mWV9luskI3LFFdC00XtMvvYvIuxKMAl0t84rvdMTB+LUZ1WG27jW4T5mnNiGmALREUE1EpnBZoIv
hxdIxrO5s3LE5XSPQBFlWJMYDv4OSajtjsAg+W2nZ8g85rFkTuuR1R87OkV+51d5c5ju/73JcOay
rXW1VpQurkitIgLFsmc6JOBPuM7ZgnGzbVXwqpm/3iomTLOnZ0GC3v4Dw+IdOB2MQT5sFDkFZG5z
74id0XEvXXA3Rjm49WbdyMDz8iSllW42Ad98s0wODJYsFNUsuKCN3/V5m4kd5ScdUrbUNu1eeYXL
4njj9yOTyyWv//J7bRaHbCrD2MfdjW3vMx+Y3SqCcKu2CMcm5kUjEWq4wFULFRQKkPhZHGBmYyGy
/wnolnJzhphIhnEiz4Z5NjqDuMQPzLEeKj8mVYwtzhe30VmNz9XJowLyM6tm5G4+SLTAfcG8PbSq
NHg2SEOgOrMALOVFdMZ3g85MB4bcBQnqUUIvzqDtvTul56PAbnAHCV9bh5TagEvnYYmfz79NMVjN
Y8czYRg4XOKma1ZwfTOIheTHmMVF+zh6KU3cvRWXWA47Ggnld5vRcwONpMGRgQinaY2D9RDqDoE+
K/1D8RsTMiHOBFK2MOQz8fBouI1i92bvh1BgGAoglOSatKgTjhyQzgXywYC7VrUT0RVmT2mznL7p
6zfHQBP4tpBG45vmcC59e+46DhUzTH7Wxk6XrVinCjbnsZIWT/x0rapIJO8reqD1DhZRALiMEzjt
PoG7G/uJyzkQA5L8pQoFiEP2MZ06Kts2X8H3OwTiKtqKfQ5Ig94RL8tgSviEjahH+heskvNuJ4ym
HSDdhojMff2tGDV2UX7OGdXAPNhS+ffs4Uvlfk33NsmR0zse7uBmfIe+mRB6v6dsMZmtDa0rIUCo
mP9oex4bZwWz/j8Rebqyr02CXNf5HOGw75J1qZsKKE9KsI+V6YbOAKErUUEFhkehVYmTXaowdP3W
M8VVrcT0iCd2Zp5BSdyKxhuvVTaywGjdbkcv4ZCDhAqkqRaENXOTUuJPobMF2HX940cPphikz/Hy
VDXu0HJ2fyUzLWN26fXiv5ZfbB7TtebTGn3x3u+/3Q/cr8m93b7QjSIJAExtH/iXLOr9uI/TjAV6
jq4j2xCtDU/wS3pWurozpnG4ubhkvX2M0qSpkiUgqqw56owHL1HmzrZ6bnLdrOKm1zUqt5Pgj5Vw
LKgRlU1Kw3WiQQZt++a6kw0edXPDOOSp1KHatgtnFikO1bnqtjpqpPrfmlBjLsx5Vyq+w9qfmHC5
I+IJ9SmMglwm0WvGjgqhppUIRbuxGZiYTp1wqJ1deKio0A/FGg8E+0Beoqo4JeyGMvjHd4tsglQr
voC/7p2QepnNphjnK13qtSSLN5JhsvDaBLkoBEoo/qlyRDfLb+5eK9aJwon7Omp+OnncDN2615j9
QbvwfAUyTeGdsK48/NnzRe5mZX+6JYSgCbfzw3j1GKYmCXlHgaJBA5eYwT8FcwsIUXT6os4U5wx5
mVnROBn1StN/9N2HL51CN8N5p+Hk8+10l24v9xbimpZ+XV+5UiRzXWJEIE+VtO4BuwcuEX2hvF5n
88Ra3+3yYqfku6yxGI/Tt7WSJM5D9jXwyNT/Bbo/HbeOj86/ar9TJ1vn0DDn5UmoAO59DASh/Cc6
2h6lNc8gSQ9PvUT31DIVNoWCsY2sDqP6+o8eB6t3QG0AUXVmv8raflFVCIoge34iY2mMeDQLsPCm
l7KVEb1/YuB04iveCuXVMueJAG5+smNYFo5CjtAWCk+M9x+iOgnj+8KJ9++E3VnvE4j3qQ+RCJPU
yeWy0/BRGHNCHBKpeyJlW4IGzJnmdpQkL7w2yGFBXD2cy76w2GPrCZMb6BRnPWwz0fceXQ5Mt8YC
PjhJCa/0tBVJvnXfWy8VSODj5B9JS/TeInmAGtwmFM/RijpcpFYfXHNFXbWaDg0RWlBKfvNovrRI
ZmyFQHcXJXmSbc5fYN4/R5Tyu1tSBJ/RncqaZmOO+nmgwzPoXdxDqM0hgZhsRRV7FmSJK3K/DCMS
8JkU03XXKrhcv4POZGS0wWRKwpbiVBBPOp7Ar4Dql/z5+5b0KGuzlJX03zxEgBfRhvgk1166pcLo
5Rsk2WW8Z+lujP7P88CiLVVhR3ph2f0Xypp304uVLLSe9u9dIXrDqg5YebbXZvvpbLBrIWV42mdh
AYe2hhCtAhLsQcM9uwhFqPzc55OPeF5uQ8BgQdUFPQJESaVZ7uPtu8xZY4iwL3eHIsBMuN7vu9iB
PnevmrHLQ3d8reU3NKyPPCDc/YCbXoR97FH0YGYEKVJ6sHfWGOlQTBajZNK5nPyFWd5wjQuF1NWE
VPRGomUg6uZ8MzEFQnCZCyOC2QXq4vZuUgRxnD4KEX16tAaKeP0n+e5W40LZ9pSuMT3jyhWK0IZi
AiJIXVJhlQdDZ7Y1tPvS5cpb1xUcfNJgK4y5gIcxdvBFCH0M12+ULRVq09MSlQ0nzxbLX8BYOQa5
VSbY2cBo5PuFIVz3ymAeMrKqf+IguRzEOjRhhuIUy4DxypPWJtdByOOD/Cr+1vjAkR/TB4eA3+aR
O6IoxY6TAQqoRwYTqYAfjq8gvUr5/aXXQ0UjV+f3/fBH9YHdoFDPi6wZg8jTxT6JIHbnRiX3E4Dl
V3vpojiRqQd6OiDu267oxyPuTzVYlrZ0MUCx39cdyggbCUtyBoRBEgRqJGv3bSDnhsBuDCVx8kT7
GXH+RLsilJe+lLTC7uA82S+gvf4CkOe/VEReoBqKycNPD/90uOq8zCr/xbf5Hr9ynhd2FvYp8xwo
WOVs9/b6pmxVwA9Do20YeD5md2OL6dGthnS8GHFLqOFcKLNf0vvhm61MGULP5NAdFinFMcTOc1+i
iATKy4cYPsuUxAhnlu/nQterigPFLx/6BNsTwbFGQmwT3ytQCQthjq0R8ntFuwKH2J+9es3bfAQB
JVeY91ofVvNhDMO2RL/lkEYMiShsIcsVw4hjzpj5URng/5loz731x5+IPapWgfOd3juZh5Ql6c4S
TCqR5R7St6u2TspmdH2FOVgNJKdoaDjLT4nfkkncYMr97+JNq5hKevi2mRUJl+gsnD8JJ4EtbuP9
0CeVVHAGrbNa2QajVUwtJEoq4PhimZB9UOc+pKPJQ5Eefz5APQ4OodL4SNWltsTaUgVcYAOgh1yE
1M6Pbrk/gAbT7BvrDayGnkGz0bpmvsxruNyL94lJDYbUU+bLPd679it5Th3qsukR0WishO1m2FN4
W6KtcXLu1B/LGPiZVFGMUT8iLpxdCdsPVaCBIuOniKL/aQJ2iTiDR85bEVB7dVwNeg8lO2AEo2xi
ST8wzf3+FC8GDfgGPCm9tJoQYf3ZZ3/ETEn1uR8z5kh3rwTvu7+LhcYunoJY38+rbk3PIXXijjQH
o/Qn7hRcZX16tDckHK8VexxqexOfD+4JXiKrfB2J9tuFr9l4qL0loPE4aXnXFp6Fq40ahX5W52If
xZQBPT3YNpLNEXG7KxvIBnc44V2oYzxbz3X89nwLShdwWVtxAwgJSLtFMbXW9zCHwoBsoTz4q2Ge
sMT7eMxEpz+56xRwVV0Lz8JtL9vYQMPKkDcaEf9I21FBpMNn9DE7HNdvJ+iuq80C2B58g8p6C/+k
uJhRrC2MAcMSiqdAV6T26tRjFdOWM1kX48zkAeQbWLOVOpMGdDM2lZW43hhd4AunBWu/Oa+3oFdN
iHixhNQONujg1THts90fbaXGl732Kc5Ff3XvudBT7ChBRaDojlJ9kur3fNn6MwdCEL/wshY6BMuM
nuNmT/T+xaU7p3B8EeAf09U5UR0jHWYDLy6124Ind7qn/JtUVn6DPa7c10+nBshSEO+sHQ0VuyCQ
ZklI+RrCayI+JTCch4SG7Z6Yd24MW1qRm7hKwKCsonaPV4hSM95TCtR62afqFhuZN6UNIfR4NURk
sUmLlVwUPmz+6iAJsQNDzc9iT3UHkYb0jX3doRd0WAAkl+pDLUANw9ZUC1b068ulXe8WlJ8At2Ko
ztd7/82/pMfJ2mXQE5w/7Jz5cLB0hyf8OtaX+Y59gffgDdchxWyyIXM6t770APEmVRjMVt2vHB4m
z2yjQ68h3/Mv0vq4Clr6XcYLSKFI5F6+hSE2jFkcPs4dEzYUkp2jc/BtXKeOcqYh/zLjTO5ZNDrN
i6U28eaCNcQz1q3J9a2sHZuKhbwhlSgvzkP/hPYN06s/I8VFCYOx2DFBY4bKLVQTUlDeoN/MZKFp
HzQWS/vcUJLXHb/ea1avpSO0Vc4SXnfuRwh6biQAcxRPVd45KlDQxTY+z6V9xJqdaQCCkBnoTCFM
wanpjEsaDwe9iN9lvaJpcpRmfthI3dDoMLLtAS1X3Xw8zF9bbM0hFPBP/WDVRv/FeH/XgdHfHklF
tMpRXaM841VLzYcTdRnT8R/JteWAYwNOhq0KnPhfVPVtLVL+rMub28NMvwWbnzrT56yB+vqUgyNb
OwGgPXZd5MJwvFC/7vi6FSxo2COjWoQDcJNC8lmwNLYqqRcnMP8RVsrQPDTs1eomaeU/gkbktO/i
IEdK3HHsfrE4wdfTCvs0ccRn3zfIvys1WJIM2L+MImL5J1ymWB8WuyyDkphnjfwWFZ28/JPi8YUO
8iLl5t2bJ8RUHotS6ixduicQde/hgfCDZHEo57I/mYZg4DEbS4ZkCgfCvEyWcgk5pSnh3+ovTegE
u4xFgZn5vT4TMwEnZkAcQWD2QSulhgU6dmxqCBFbG8PRX975rJKyXdQuZIISnl3DHHzuI87Srg/k
TW1TlEYE4pAimej3xt2IkbZkX9unMGzIkThhN5cGPuCor8wxUsHnoyx3ClYdNu1Bu4vD/SlkZg0t
Qehk39d5g4M3YmstHnVWn3whiFt++pVGlID6ZV7dx8gVCvHQROF9DE1oO/J5/BVknVks9fS0LX8N
qT1ITDqNA0pRZqNlCsG8KaT0Y1wPaXqlVu3+3RxI4VEpeNdDh5PltI6Vjk2QF0XIrOlAeKcqDfDE
JDxalOUrMH3fKTV4fkQI65sRZ5J944hr0Ear3ybOaSsCiIgBlZFqhf0X9wEDcAXJ/YZO7pl5EB5h
0XhvY7iSyjrLlfVxaHWdNBtg0qwTJiJ9m4d1gdC8T3PVaKNGdN3fW2BppickhOp7QRU6qodjXS+x
j/KiJwe3IYojLdpKClIttK8rYsDt4CdyWX2WBxKpm7uZ3WVtd1S1yldeg5hMVLypIOB4FyDKfgfG
SLgbLFfAx7tN/EzLQ58wEzHMt5jRQjpA/tHKR2vxAHOdvWd8wfqglZH/tnpFB/Qex+c6aGNNMOQw
Kl6mj5PdESXCTkxrouVO5/sQE8LGf23C7OtrhaKRVXkoOFn1fpxm5IN9caZkSJtLhky2WWzEfLdC
XsSLeU1sMdxX3d7vRqHiMKcyOuZPhU2YMKEFmr04O40VatVlbIjgw0CBmGPz28E3nMaDKBU/QBkq
EWVjEUGBCgwhw6p9S3i+A2z1KkGPoaYIWrqgxzrcIThoV6/9QFNP71Qd9kbUMZm+x9LYty8oC2nb
vmL7qpRQWo91MuGZl6Nq8B9HOG6Z6Ku4y6LRJhBhqxEYQwH7c8Dyyz8YwizBcLSMmne8tt4vzV+I
gnl1TvUpmViB6Jz2xMVCvPsINGhHrPYoDzGcZqxj9cBrjCHrVi6fxVTmzwzXT1JnMfFRRbNNlR2M
9JboCS85Vgjro2xaCg9PnuXYvOxNc6/Wdwn/i5DSLNtk8z4o9Cnqkv8YhC0X8dQAM+bHX58mkDVH
yUxQa3lBRVK/jlBw49IdYvUX6XKVIMB9NwcIFa5YXJ7/e40J6JOaLLDg2yF0jPhNfou5Pk17IJWA
SmA0O/8QubhS95y6VDbflizna/6/Qs3Kmjg42/aHWt0aPMIsjkRC6xZ2tFSUZ0Oiw6I867c5UGmC
wbGFl64csqcBIGhZSu2yWJuPw+5+SsPfS89m1piKRLlF0tCgeOjmWIxQcCznIIAZsVD5Q6HSGKxN
7NyYuXy83W+RWZ3DG44um7dN2ikoGE5w9z/3mcaQSSmJtGn9SuAW+EmOriY7Yn30wOtxP1GOu3NU
6rswcZYHUWrKWCdkw3NieP/GnzAZw/HMN+YQgcaH5zVfhkGyA5i1I2pH26qjHitOA+MeFLfFB3hJ
IUd/gGRIe7Pdktpe1mLz6Q+E46YD2/mNjDMq376YL/zUoTRvxX5n/KRvgqTSb8Oj0pqD0sWiorjj
1Pv1JXGZ7QtoBspTRCNjLAACrAfDGyjmU2hc53JRQDXKD2ORFyGMubqlEQa2dKfE0oUgEG1V9iAp
5E+THWQtNfN2Qe5/9+zppR8Liv+BaBAKsh1cf2fiKbqkjKzO8csVfnLNbpiz7kJNLfL+PISEZCT3
fN6TvrHp8wS62g5srg6B6Nh3eJJHw8hPc8UsDKoiDulASsJqLLZxH5gl4eWLe9RKZi7fq1KKvTu1
IKk6/JD4/NhRY9D2cimUktk3b5oTGtz5GwNQ9urBAkkgL3JFh53lVgFvUNa0ATHEg6AMaf7VfOCG
UZsf/dmb7bURvPded/mAImluJzKUnSnWYOqlT4MGec8BpVuJs0wrPFLBdfwZBhBErf65ok6r9i50
/PSRE4/GwiASzQF12nhu0SUvEH9O0OJPENPah6TRe2jYz13KkhjpNZD0082Phk9IcdEA2dsgWcWS
kepNMphs3jCRdow3KvxkZ8vBg0Ggk/mwsJ1HGIup0eXOhUUzt7f1XunfpkoU8bL77JoO61AvtYeL
0zFYrdnkJK1sYyZUfhY0qs9OMj46T8E0jwsMHCec5QSXi6rOzmmQKVVeObfOReS8h1B/82A7IN57
gXkED5T+rF9m6mnWK55dyWqRyWnvIlyDoLXKCzt/4SOe/dEOrrmBJm59bWjtwx1npwNod+WhElcc
y+xaddE7r6Qw3oEL7kzHSUtucEYSRUd0btpfbF0OOPe1oRH1QXksbhheCUFe4QZjd4V1PnMHh6rY
ALVP5XD7+nxWRuGkGCp4pPpa71hXbpurpUN1dQ5EUdFVRs8rqOlqw06yFYQLdtB+RjK+a/uUJJ/x
T7497UEm8qqgyOD1HzvM8ZmExabrLNFPmatOWiknXZ2Y8rzi6DcGcojHudVdqiBms67LEe1hYK5T
AGI8cFW8zdCNjWkYAIo7OVVu7MTdGP7QGSvkuUMBR5NM7BMYC4JR6ImdnszvzQZXBfbczmdkUBbf
ayAKrGQljAPdj6QKOgMnViy4M7a2jjgPT/WBWa1dWYYI8/9djdHz0yhBRV8JLlyU4SSSpW3tUoND
Svk2WwYkN82uyCRKbOml6KxHeBhP7Aiuj3237T+P7m/0PhwoJ9ODelki/lLfmOIt7YYF8iUb1l9H
d+AtfHbVTtU3OYJsuMLlSE/pvg/ft+yBUrN6yFGddiliLkzbsmBKOTlR8GyYtwQuUkkahat00MNC
6jjk2gLy7NGNgy1dTlbL3yqMpb+nqPlwg4RIo+Jb0jgLy6pc9B4npqSP7dySysMdLLQbONBUw421
Sxo88+rWmta8Gp8QBsNaaS1kadnNFkHhK0jGnVFXG+Zj6RqQ4F1KSAiU24Qwo/6czLNesN7yzSI4
Bgn+sfZAtM/j5wPIwLBFZRYoR36NgQfskKk6TbYoeXy9/BPWm+to6N1V772/1958PcDe79Z5fMvw
xZD6rs+bI6INAMYC+L8WupREdosiLL9FGk+sJehuW5XV4aVwErp7yG9oCNZwXdGDld7s/lM6ls1C
GoB8u+7fa1Mn05BNEy4UwkdvdUiJFifBtXc5YrGedFdbIH0bewpa62KAQkaMeedgWVr6a/ZTQiar
g3CmBmVy2D+nYOR+nZXLgMjpQdsOELfmEPKCh2qb6uJXwkL1zsiexD1dUCOjOZeTkKZkFKUr2BN6
BbVxrJqJHLMK1MUeYZZLy7hV+dwHNJKum76ckcdRppOPwDLHc4VHH/e9hhHXv3+49T3Lx6ZeqRQx
Y6k+mDtLXRjdcABQWy8tOeokIhvWQuCpOW6iVxh+c6qN33AHhOqTOZS29dwgIO6jld/ihXyxRC+8
Cqx2VlA/fUR2qmnVaGhQASnubokbKo+al1+ER0a8FHbFK+450aW91JA1NRGS04OgBIxUww23AHHI
9ghMukMLGxlsm+IOzbkxLZiK5JdGCOWdrx2V03PyZWaMok5yN52PmAgiMfYhazg5etxx5V/CGB7B
cb6EWtZ2HEe2UfjnmPMaBLsTOT4CNu+H468OCUvU+UiHOQl1ie6zGykS4EZW5YkG6tWh4tJ7sGlx
uLEtLMv+RzyfpTdSNOkCFvH1R0wrqOL950pdz3fdwD4+ONEEGi2VeJGfxOyK+skSw0+nH1nLnGtk
7sq7kNXMg5/SFvDqn9Q+64HMWaXa1+RUlaXasW2U7rw2wxYuhLofq/7WjaMkONQeRMtGuwk0pYst
JTCfN3xdKJC26PVYvYLsE9YqxOZvvghaKNIlyUkSu3EX+N/X1x8Jp0xVbojPKfiEI3MmX2qnwTvq
ZDJ7pkslAnkBzuYu4OQ1XwnybhjlOGNik6j40oNKSNVo7y8lESBtjMjMFN++Nv8WlYDm/YyIS23P
F4ujrpVEovz/spPdkinODC3VCNhcX4RiV4VXkD9lYJYOPKqxNrNUcgTvB0UMII1TFAyRLCp8CW8+
FQEodrmdU2uzBrz/3bM36l9Le0KAsQv1hSxUQgtpqzH3cmG1pog2WtIW5lu/WE1khHpu00vVQk8c
VX9ZC9WKaWPMOrV0VYi6Plu6zlqUoBi9/W91loknXxJkpGgb1nKOmEvPiNfuf0IX0oJPGUtR/Ca9
DqIeyd9q23XKKJVzf5YGgGxYDmu1J9hf71qndijA3AztKzpcIqeLp5LVUPA6J/jlUWg3q+e+fQxw
WV5zF9GseMsmrGkP/cdYWIvqy7K8UCKDX+c4lbwgXLoqBOBOjmyYPW7I02wb46ksYKIrXECR0Ilo
FK4n3mbFkPVYXtQdbPbto4qFnKEFI5d2DryLc7PQnr9OzP/inr72vhWg1nxFSz64KJ3L21UVfoEN
NTHi+lJVTX1Lk5vEX9ypPnUyOdsyXEsTOJi793hAZEC40Yvvpw/HA0pk3trWwUv/5VRicqOyVZgN
LYz+ThKCysZgObVIWDNdLcH9DLDtJfD20WEB1goEeCk9pxxZvHCO1izTIH0rvGFqq2LihyhtnxH/
yBy4SZt/DZ6eUdiTjpk/LSJlQqDT3Ey874SC3fFRStuCiuDqTWlbq8am7rzL75r367pPS8DvpxDk
uc/1e02Xw5GYN8OuWuFwoyWsFFWsHZq+C/MiHvkTPHwesSPQRuUVeR084Z5dw+Gv81W3H5HcrPAD
6ErcfwY94H2aZNe6gUFFEkhCc9uc2UhLpHEGIpGXv3Sq2jsRTUp1vo6T4ZJHa/riOW2r2ZnxWG+W
HLH+m19Wv2+diQagICOMaeWPEg3Jhho3HBUnbbZOXFZIeFd88YehxDFBN4JAmeE0gk6O92ThRI3f
7OlG/mARci6UxDY4pA67lmDy/QVpjKf6axGKMNvMJdqEnMY/CPOIUmu1lBPGcltiSgLHdV0aAdCP
wzJAIOUWsXKh6ZA9gL8LkPg/36EaQkHPyGmzsnkov7LaXteYvZVtfBj6oIw3B0UcnQc6+UF71kE+
xFCrwAdwqIkJJjZTIbIFYexMXS7ODIwbTND4HKtGjL4Y7nai6NKnfX9Qc0vePwQiJW/jRPlDFhUX
7m8si2hEldG4juGUC3NVjIqV+R0Ahsh7GH7dHZDLTNiXn8/q8dU0rFiFtTlU0l6DDb/KhdiGnqFQ
PdT3Vu8te7vi017zNWvJXcJxtojc66p4iJD7K1MLAdN+xvOb5VS+2SNZX2JJu2NgDt9jtTRqY492
Vo7OpIJbqEe/ekywyAWeQ7QxNw/5MvzeB9apTp70dEfJGkrzuXvE7+78EVdZZENx8yS6ozhG88uU
cT3TLeqK4Kq25iJ9XBX47By8ratDbdJEuKYuXU9sKg8LbggEeotodzJbjSj59i+LDtJso3ihgUp6
DKr6bFSi0rqofGvSSIJOcZj4nO53fZhZqXqGvKOlw0PClZYnV9EI0/GvNrsy3n4pA96izlQai4gi
S4ZQhXuA40LQ13ISMoY13TlavHOffEDkwpLejklfRCKgaj+7FrdbHGZ/N9T9BP0Y9BEchCjm1Kc7
tObr+gGw9Lolaf8JSvShgmShThQczJCkWsqETUrMw5I/0NOvjs4DB8BjQaGN0+tTkUu0rehvY1S/
ZNRTIK8h0s+pc0lNS8WXg/EjTMv3PTi12qLIIFDsYfoQh6znipbvsOxsM9nLXoOB8QBPHeVdH/YZ
3IxpmOeC8Qkf8fq+ba+MtBUzYBEdiBp8oX4rgVmzmSfqevxqX90XkfdWyTNhTSpwIfy+Bxf1oV56
rXaxiD3eMSrcdEOn+CqwcYmCXNMvTsp6Pzj717w0CX4SztqDxYxk+rgJ7eeaDakrH2lWns6Dodto
Qdtb++IZuw5zKzyXLMVxipfBr6Z8gIjaiatV1VrMP38tilkPBsDpKtNAw/2k8bYLELAGRQjVOjbP
hhC47so8VEDma4POLA36shVa/bTGzD0CI+hbvlMmbnq4pmW3LazBnlqtz2G/UNuuOq1SE6xvNEqk
ZADLSGiNNMeuysG18ISOVBaCYP74dU+PTdB8ZClXBKOo5gOcgGfFifkqskPndOUUztLrTiwT9bbt
xmpzq3jeTRJDtLVrTMDe+ZmSo2wOEh+KAUhYpomEd1g8eRSvYPQ2+QlxzUSG6SMThNjrDAsqZJho
hONN6fl1vHgsfqfoOzBs65ELIwZCKxV13SiNL0QPmu0F3XDEQgJQU5gbh2xyaAwq+p5UvywFIb8R
cNmNZtArzASzxQMxAPTrpJ37uDQq2TksdE9AjUHbIMzvXZyYKqd8vwNc3tbOgfH4kACim+g8ly0B
W4R2J2vzCx80hLblMhLTubOx86uDgaSP91PZZ9Y9lRje3zPs+6sEwMxtvnrPqVyYqBQqVnsg3w68
vqkjQpHY37QfyeE/L2fVv5XD6m081KO8VTmgPQ3A513Cpp4lUOI9wQ+bn9wK7OuAIK8Ji81ZFfOT
7H9IGYlRntnGvJTkdnkDlLG3cCrxxeE6neSnwW9syKJxB2SEg/CBydA/XsjyzuSgJEZ8kWxP/KW0
Rz1bSQq1TBueKH3uLEJufTHQdFYaov7tJZRUsicrpRUyRNmg2PaQe5rID4n4wp8brcoUfrDHhK6t
gXBkuU6pdD5ZBql+Q6NDnsXJMTi7a9cF3+J4656JUOCEotYkH+HemYJIX6J61h7Vh+rCE93GeM0N
9dpcRgNy1ZtFANPVbsrd8MZPf2ew2SIG/d6KPSimwmecwvSiaEg/wfXkob2YmsaFw48AEz31L5DN
JXjwpScN1BfHhaSjR26xoaYSSrcdcpHz5Hr9fJODVYR9vKAvfQTkMd+075qOMzQLloqEbOwHz9ea
mvpIUserqZ1Zv6XY4XtVYAZg1krRwrtZdutHVCisLGvhFilgNBPEKI9oXMKeKxS8J4YnCZC/6hHr
B9NaCJIbOMQmY562Hw2jVq8JLOkyJnjpWDcn0SMJzGIl3UanFt6stf7Vbf0Vaxj74voXsFwvPCew
G9DTkn1dJsh0sPQVSJF8aP9HZ+qJ2/eVtL5JVAn0bCkU1sfRsVeBlKD+W2is07sIiIo9tB8EVl1y
glHj3H6JMbCeZk/a+Mq+1d4zd+DvSHftv6RUOLeDF8SIMovsfWgzjSvWX70YSX2001TvhPBKdMcG
ZAhOMmyiDjOKpTKepzU5vgv5Y56Ix/ypoqzmpxyQqx6cFj3PBbn8bhBwadg0xXaB0EnvJB6cbt/x
IHMWYwLd0nB7lwBqf6mG1PysLTzQiLEa1xJYOtqwyhdc4OUS1lV+ZWEJdrDpywYe6sKqRMjUevlr
Xhr75v4+DFqgwGF1cJb4YJ1T9iSTigUE2S4jlU8MYmccOFXZEN3QeqO7duDdlQHMQ5FXcEV2mtBd
aYqdQKuOgSw9Qf1mX9M7hxGhe80IG2taWGNJ0XdJwCLbUlB/Ug7Jo1ruIw7UQwn5+gIwagOXJzMw
c4vdI/VLxoqnRuFc7KtsWseym7GchFBvnZFFZ2tAG2QYsytRiRCMsGDiwKptpNomqy0LLBSEjO4C
9YuAuhzVg+2IYCMYAeRrdUeUKMOjB03fbxvay6tI0qU6WCf8/Vm2JBgMIGoxZkaiMViqeCFBd5Sa
FlMJijmhzU3RVrJyCHrpXqVvtWWEu+2gDAx6G0qfNOUrBYQKhEUgbxLGkzua/OMYxsKZfVsiVoJS
qpvtebr3f869EIQHQ2wYXtSM0cJdif3swwDswDSOKu5uP6wqXR/8rbk88QnzPkNnYRZU/awLWduy
Pnye+cUMvRA19+Q6ZpNjVD7ACbTK7+PyUlwcNfh1QbOl5POMX6aKHQkiQZjonueCrlNX0AMgpiBK
ynit+w+64BMryIValMYj0Le+cmnTzIirTlXg1eYfhQs+wQOx23t1CQnyHZLUJv1olFF6wKBQvrVx
y1pUgXgsaGuAA7yDH1eGWiqWfq5Cl69pnf9d9yqVudDhP5kP+TxjInajjqKp612Zyd9Wdkgaq6s2
Il8y7mMUZp1GxWYOtavaxMTCXcgd9ZHee/PoMpRhs3LOCNeLH5iXxpzQoirU7/ndhz57T5LqpW3Z
lNfhkBOgXh4idLLQn5ruE1HkH3GDIbfRK7VOgtynwkl4E3PEhbbmGsiRlDmaE8FmajlaNuvch1+A
pKHcj11RMVKcGU8iNpB9gRq1rzIt4ySQjgJQrj2lg3qW6DlKn1XO7JyN4MQhipRZ56SyIzFBhRlz
POyNxwxqaqYfXn/hGYryRMIb9dt6vdO5vl2MAm8Y0Hsld6VwCRx4DsIqVuj8qxqmGJ17bpApS26h
G81iaAo/nmIICXetBpgSgvHSL7UTtcqhGyVj4cVQTzhuqCf7Dj7iaIgQglyyq0yNVBquapn8ej/C
JoH/ShUgxNE42wgeKvMnEQAmGf6rk7kmDWRTcxgWVsw8FsLM4wjYCvthV2Dduco6i5gpp1ohiwvO
eoIkFcm6+I6AJbAyJEK3ZQwL5ebFFrWXHAyDsq4uhM3/vbVmRNbcmwatbxk0blLM1XzrrnxWMdxX
GGvbNhbLq7GdujTSmAqtlExgm0wZjFFeQzw/HYtaaPZCXqwTO/WzEkvYfKxgqYhRpPOvevzFkScn
tSgfImvHNIWox2vkH2Q4jue8GURRYC00uWbYJPkH1+NU/6E8jgQ+g0p6Bfx7gbVvr6nxkzCsfCew
Rck+zyslkwyx3jit8rcp79nar4qgIl1po4NhO4V7aQ0QQUEyo1zQQ+2ZXxVE8vZReRNIXpdNeVq2
uRTir1TZejzN1xcnJDQ5gNYBH53l5wnqZFSbjES+21pxmGHUVhFh92+OVQYOEAPbG4WK9M5S8Ob1
YxnHSVwvzuYF9JFR8kqhAbMAqm+fUWW/dJRef125/nVAlXRLPEL0VEipiTxSNN7jx3EWUbkqB9V2
KS35L3yyImrCYWGFAjxvcoWWXYhNYvDte/R+ZlUHUWw81XpRRghZk8Z2s0nUFZMeG3np3zLe5puH
hG89n39rgzf03Ywq7xQ+y3X8CZGmW2BZYdkia7h9QLw6kq+grCMOyPq9jxLTsS53AYY0IAtn6NjF
+CpAL+WMaV+fw//6eDJLCnToar3heeNkUyT+tsGQesBOAI4LnSLymFmPpoW5jxLZdY6fC4qsb2jO
MxFhIQvhz3h4cQs5FXiK3SSKMOwTNgMVh84wJRO6aXRcWohsSD2JY44Na9fMvmqr6ipFd8AKL+Sz
Q9hF/bMwbPMsM/SpDTNMGApOpQ6ku4dtFa2JIqkpk+OOznPIHWutDlAgVFSW3GncLAlIfCwzqN9q
sPfWm+zhfIHdD+qoPYXdNj9kInJ8UwVRC3iTfGFFMqJ8xNQE8rJ68ludko4CALvxAvkaVws7ypnt
SJPWX1T8kuWUI9m9oKtv350PvqYfBccx8MgDoqXO2ZxenMlUSvynGt1ZqfCWf9oY8bqPIgLlIoSr
6YquG4m2jHdIqCyVin+WZuIDV2yxqP7hiw2uwq/8uHt+MTnfSS2Ivuu7qUkE8m2J/0bBW3QmUibG
yHHbGhpczbjlo5xgxEMz5ZcPY0qzrW1YbXIJweigZR9TJKg3SoTBA7dM1mvlb7yxb+v4mIwOUauk
t/Abx2PBObIzbw7jESJVT2fj2PCU+KEovZ/vFS2BQU8KS7OjjwWSIe/ID1GA1rNjI2aPg+scAIk9
EJveGghJMolosXVZv56Ap5Kir+5t787DhSK0v2v9j+pwO54NHqpFnwGP7nZDpKQG9Xoe5XdW2bxN
i/AcRvAhH0rqtmVICSA+KnDte1NRCUAHvbj9wx6aXj/13D2UoiKCoPEb7BkZEJcTRmp7Ek6y8OOC
z3Un0N7eMaiST62bBEdajIOV7lgD46p8BBAkIMH2lN7iajsOeT/bMORWYY8t35HxmcP7qqjDCpXW
NajxY5R8c4yHlf88aFBWiBmb2pmDyBDhuXisl173TKFLfVPgYjOUu2jpBx0MtjAOe6TuQClokdxf
F5koUpYJe2QGXQ9DeRBHM18VjBWf7o9NZD+agr8t8rO9ch1KpQRkxCJWIUXYxjswtBThhLBP1IOU
6d7gBcmqqtSx8ByEyoyPSnzaGcbnD5DaFeDj4eHUZWugLOMTKJs4a6NmZ/NrQYFfE8W7IvJvmeWD
DfzQIpuVVynQRLvFR/7ZK43l4tX/3yljGPG64pTUU/NFx8pAZHz0HloN5zRhMJEydiDR/9ScNKP6
gw2oisw3xMeBk0t3mKBPIoM8/oST2UaduXzfTqyCGz3kQcJdJWovl2rF9tmIsMdhNXcqYLOK4TKI
J4TVFhcYvpJJMoyx8s9GG4eOkFb+4GC1lAHzstWAwLDoNKkNQIrcYIw8r9jfiF1xaS9PUeXnQxgp
JMlGr/pK838pk0nTDds6073uPC2RoZO584WOax6LABuuZ766/PYSU4bPXVO6BJeIop0N6SqfgHbt
eahhdcrG5VJ2Fp7plYE2bg9w0nfJsVfKKAp5NPcLv4fUmxZ+Lu+nrw1eXDiXdpI+yRT9ByNIQMr2
uZOdHjJqhY7WuZgnwD/AyDyS+JGbyC06EbS2PZb7UK7zd82RTz0N4u6PjsGZyZaXBvEH4HBIWInI
8vJGi5YKTuss3M8T5woQbewPUrpjLZEDcc0TnqfURZUMeOdYohvmypai9QPbNEJbXuh4sLXryakw
dLk84MeU8ElT3TlWd0lCN8Ls8j9IOOD30LCYymKn1haWC6M6dE82WMQsbtMCTzUaPLNKTFnFP1tW
vNNXjEElrGoew/jekepJbucuYfwoBcYr2irT0oKgjzE+T0JO0q+Zp9f7a6cmgPEKQzfB5ulkhMb8
fAa2iA1En52/1vYFbrSC7yh5ZcC3ecPd0YrI8WnDaKhIt64s+JrHpvC+8hhJZOQZaXO6hYTZC0qt
bifm1Ay+Zs58a29/vY+Xvg+VvzdHyGcx5P9ZOo5tixW7gbSKkG5174nm/6JW6cf+7OHMs6AHnEY6
rPak9751pHc0BX/hqdaxtS9tsPhotmORb3zOq7KCEedEduWVvlQ7vvlV0qDIV/6wDNpiPaoSAwLT
1yfb1MO4hspuHjsLqMNbc+qOzuVVzx8Rz8ipitg834aw/YffRPW8yHWupXD8UmSGdHTHPyTl94lx
ph48t2SkAxyv22lR+TZ7QNvaUC00a64Q/KWPP2LGEKln8qGUGdtUCHhHPBGbGKCYqzqGd+kexEIM
ffjV0qITfPXzpgWEZxWrADnTNTFKWEqlRiOF/FluTQJ20YNpkccPOVkqbniINwgiYCqIT/Fc3ZS4
Hc/nvz+WSLZSpHqwWmjbQ0PNzs9KYe2aHcJJQZ+5J5QAUpf5CHHQlVzhwK8OfGwztiH5TzSafiFL
D9Lv2gf12JRD3IrvVulaxijQ7sVFFfOd/sxbONGBFZZ8Lt3wh5EzEimfMlyR/6tGGf1CvjmQjZO2
ScQtdEu16cKj+hKxhsM8UL9p2QmbyFnuzGRmfW8j0PYgv3KLmKKiMqPxabFwJvSrdXdbyDEs0k80
W/SWTAYh4m37kg27jKVxpdcUa+dtUTq3LJIkuUPq65XoeWH54xlPsgyeejtXjjIshZkxxLYFqhgA
Rtbc+zgmslc3P8p5rb5LZUqgo5w4GXzXXytYBcs9/SNqhN56O8OMg6KhJcFay3PqktywE6qVZ1t5
0QaQiFm6r4BlYH5GkZXC0fJN7yAtff4obwcvU7T/MrP5aV47iBf47/3CIJIgd/e1yH7i2GGI+kt4
jNqKT+/XwuDtWRcRpKeOcJzSF1rAvnHgTczFm1yrVlo5zlwK1YjtMy+E6JB+AQzvARLFIZc+xnui
nKptNnCPLHC9rM9csKrVeqDQWkdncxvLxaFdXYzPYw2hQ/DXk89Yf1SiCZEZs9fYA3ULjWB6nd63
37mNLSUmkmjtJgBapOVnfrsslKazoaj1hywIep8gi5rv75CYCpWfc0Mvu37Fqd9HNhyM0B8p0Ym6
UsN9PpikSxnWn4lBYrHF0j1Lg3h5YuM55jJqU5ear4o/g5hXhZT1kARYQiyhqwnl0T7ZP5q/lDnw
4nZWh9i0xgVW+n9DsCsTKjxylOvjsd4uJ/m1psMjsINJZi6/p2i/TAhOvtJF4KT62wbda9mbZuiJ
XDcykwW/X0Yd537Ju131vNwbaJgRsXuHZrCWt2mnjeO61Wfx/hBW4xlJgmmHHEeWbky8lPK0ge76
W0uSM5pK9nJMSCTuQeFpOPVnjTo7zl3knR/oj+uJbpYqCrRsoYYZEWnLaqOwYbyHIRE9veltbGQ+
FiwLTGhXGwymwOp0xJkom9Ica7GebIZfEEPM7iOWHWNLVKLmyVOXIqK2PgL8a/i5ZaD6cUWWT112
QUJAeOtKlJ3bjtSdLhZ9xjvJrT+IODo64ETt/X2A+rdnHZt9ablVIh4WZdBncq3t3ocHiLVRmAvm
jzoOHhBz+ZI81kjhCQaF3HYYUDKSbCbKWMbOi7ALXiY8ezeqgZ/Mk0NJPBCLf2yNP2+R/EV5Ipoz
Tk8micnPqlq5iYvnEalOcuV1TsB/jmSr+vqwDM8TgWqVbV3dUYhh5ZKLDGsa91JHo1e9nk53Xq1l
qVerHKkl7mKplrHiBgUqt5vFmITzl/kCPF8TPgkWPPBEgYOQjm6i6yXe9n5Vjr3ElYiQOuQJSyeH
FhiJJ/3uPIVDzRGsHMlbMy9mi03i03BUQdkyPsdSi3Dc+Jhs2ZTn86jZWUatX0nPKg8tnVkj+t52
VcNeNTgi9hxYlT5Q3zVKFpVCZ7jnRACaSofvXimR57gOkVS3ccyBhZonCxKqHa7ubNm0nbXYqMre
+hHfFbZLobvdSTl6fV4KcqFDxgZikdBI9njRfa19uTsu1OXiqHGOoMjozmKBjIYaJh3djeVOujq8
Tqqi+qttyE2wlgzqV9kyQF/6Sp4X3iz6UiU606HY9Xmd1irgG2Ci4tH81QUgGuh66BT1JD0HOhD5
v5YoJhL7Cwm9JpOzc9Ot3GtJqisOfwmfNEaqDijrMu95QtWB4PSVxy+DV15rbCnh6rucylYHlaH9
aWjqr2DZnr6pnInGFg2sjF8RK5+PTl0KYi8XPqTP0wX24f/Q+SXPGqwcxh69ZoJnRO4FT8N4vhFc
fRAw318BPNIMqYmkqSHnsqjnabGJ83y4Kw/4i/BwctA1+B7OKrAXYxkg53Pq2HerOwrF5RA8YSib
lNRWaj2jWNu7mYMQ++L75q/vIojiuWCHvrqlU3qjOnKsjVL6Sx47h5lwnvheTi1coLDVaCYP6YYH
qUSumDw8KKQC4QnLGXuHxt2wAqbcjhjqAq3PDmtHe/7SC7magPL8Npta+SATVhCkpzeYTxDGlSCA
dNYs8Tb766GADlLWF7wmoPkN4fD+DrEk7iJJPQi/v7KmZZk7QgGPSE8sZ1MIa2bXWKHMZ52ROrvm
WatVY2nH3jCbo47BF2MC2UqM0prrdBj+Ur7VmmPukRkxEcwM2TC3//oYoHIrgaXhn13yWiE2AguX
VBy1L/Y8aR1AK9wAsFenNvIL7xc2vTcux2ujHTuVZMz2XqC/Uv9Gu9VhcllbEsagwhaBV2N84tsR
WmJCq8GS5D1158ArnaF+hIHJT08PsQQ7w+PAqmPkDXSHQPkTJftipC0L0pCxZT40RaW2y6mhgZTH
jKGE1N5qjC4Co9Z4k5fE46pT0UpuusiHQ5j3V4THlZNVUtYfC6zxjELuLAdo0HNNy+otcw34h7TI
JPmnbpS29+VGQXh/+Ws/sv3/Ju9aWChArYs1nTYQtYnKH85pVID1mekUHsGosQwqye21T0sL3KVG
fH1py7yEVzj1s/h8jSVlGIO+Puff8KnDM6/R6pz66aoOXjq3xoAHvCK/bqWmMSJEsKj9uUYSqg/J
G6oAR1WTUECaY9Z/NAFdGr2ni03i5+wNF3nSUfS1VkD6TNsPFwhtoHhntp0SovyjZjolinaAplYt
lSrvOMkoGlEjeItWIFICaGc9vaqud90ZgGIwB99/dRaGL4ShAf5iaLccW3zK9YpJFyoiZxRWUa4a
SR6qMpIeckIrBpve1bE4wCyyTgL4xX8ChbHnP9ZTf7NqUhfyh01lCyW9/QJReAfV6NaxFeD0CJA9
mVmJaC9gOfJTn8j2rmMLgNMxC82HJKtUJWlIVOoTO2Ri9qphNOn1uDDzPhns0g2c574w7vmMGI89
0Ba+k1y4XtCxecAPmLFmi99n5NpHf8QhWwR0j+FIqN1lD58zKsAg+zss8qT1vB+8ezXyCYWGFoKJ
XQzmnU3WPGteZD1omk9I4Pt2SFUtwtjbdBF35BQWtlAKVxNYd38rrVXKr7aOWQ1Q2Wd/8t996ZtX
SaRNojqClR2IaEyBHV2vkg/6A9Y9NSb+NBIrs761SFI7MpOhCn7QrO5WljIMVm1fCOuwxjIq2To4
jVS+NQYujFnCJU+/yZ0brAVZHFRPtSlsHirbw7TwOrzjiiGc7KHf0ORy9n5R5QCPfOyOXs1j5fuv
tLxdiB/RjHvyI+QJEz0S5d8ZyjTTgpS8B1JfS055cc+Sez88rG1OsNxoB/Gam5NO6BV63E32JUb9
gXmwLbTGYQAs0uHG4QU8piKh8kGklKzh/FVJctSWiatM/MWltS/KcpXYoAJzceflMKmdxvtS9ykQ
8CWGv8CX40hQVqlvmn44QIc/Wuug1b3sgJ4Q67fzfpFjv+cJeKqLBXMwpMjaxJCOjozA3dFfpJDa
9L5QFIdyojFBQCWOR16NAUzuTeQi85eQpObZ87I8i1Su3tVzr90+Fh6I1qfdNrX/wU4C92hafLIO
jP0w63IGi3iWUYvIVYTb1q16+5I7aqK+QGoyqpO/ABoZ+4ZMwMJLFn42R6f2YfcTA4mKfEjrFS48
D3FfkYUV3L7/R+Jc7ZwILpl+hMSZPubVzIHHTeC04U7y7h+ShQ/UyVw1+kpFBmLHYpQpcsi45DJ8
hfuAonkmTNn5EFXMB0LJ6qe52Mo9nTYiZixSozY4TdWVSD3KUi9zKh5AOVqJIj6cwqcktN03WXpd
re9fdd/49MiQlUD6pXIRWZFHexaon6uFa/Bbyhuq98wHjQjvb5kmXNAfs+4EZWAwyT71XbE3ZbFJ
uNnPNm6iPWzvq7OeurOf7eKkzhjiuUxEACVZj0y/zMj33kOWxYeae7FxkE4H6+jAbyGGz+BNjDzJ
Nkqp9hRtm3ldsL0bUfDtB5iNofb6PvU9s3FxKi3pbNNb2wgCZQGz2gTaxvJjengK8Em5dR5JQ9+P
WHJ8fts1UHwOtsXs2jRY8ePlWsRHpRkCF6CIvGcAyM/1ES4aIxgKz2stjjXjorTrmx+SSxGzLnn4
eQHCRbOuwjj178Y5IeaZjpd1rLdHwky55stoyEU3LxQ2nXhrWKQh7oQCwumRAJ8kcNxOUvUnbBF7
P6DTsplWlejv4KNgBLuMoJJwTCQ7sx1Q3cyxlcahumf/WBz455rE7DjIzVfWuoqE8whQdt2E4/N0
HhDADNLmx8L02oasAar9JQlvw1dcB3J7ubK04zddHzvDzUcWf2lDYDuaOldFO+n0vd5nRWDq1ZQn
pB4nLKRoM/smf9voZMmBWwqytFyXvhMiBNknuiq9IHa+yYCcsEaGtg+vT9tD7DwkRaSBhni++8c6
j3/UsqXxUp5RHl1JEZjVcgWaoTRcr/POA4eRg9xww48Aazj94dzoU/KOTg6TgL8RJmazQ31ukp0J
EOGb3InzqHGaF7S6OlzWzMKDh+sqczQzmNA72BQyVGoL2BndUJ55F1EexYXMqUzw0VwY9q/U+lfO
nIeK2mQb1adBFicQizbw9GP+sbK/TkTAxMzbWRY8rHvvN0WBj0SQCp/K6XGQXdL9yw+R/7Ml9vMA
Nf5P2UL+4ECAY89UMarjkMd1IXWtaXF6HvE3Ml1qXjnA2S2R8LtT8Uo6TkF5tkje3jSnFa67hBlU
roeNP+YOejZBk82gooXF47ipZIbNGmMvglaDLBeu5P8dsA3YBmuS0XtV/0L5CcBLSAXP8grio0MN
p4pc08rQ3rnn5228VhWYADs54iAtTD6b8/mjNU+kp1qbllDsm5w2S89iuQz0Bzkzq14NHKsipXYZ
EbDS9MyTWoFfMsKIJwAVX6norB9+09qDsAzTJ6Wz1bcIgJsJaelHQoKsQgPfHuppG2FztBoLtYu4
HMQPW24GZTnm2fLfgTHswupmcAWkZir/q031q/7WhyDfQLwX7BLx1rBwI+/DastkY5u8ao+GSOO3
4jTJ44POSuHZ+qam9yWjgwszYlG4FDGk4E0AACMtIeJ7VTE3zet+bdpdwhcLJqaK+5f6F08SJBRr
g4xJvFDOBtZ67C94CtXQE3mo5r4R1v6aBk56c/rt51A8ecFZdg7QdfmKe3stxaId1+NLmdqHQYtu
e+lqKmVoSBQpqLGnI2nFmgNjdBKdtpp3sVWeQ5hlgOIAz5RUgRsx6zFMBVAiewUOeXlWroCyyAt2
99N1MOqDuldhWkCl0LxgkQKgSLa/2KnjD+tE7IfJM+Nsn5SKnZ3ZOz8YK+XmPYlkL7W9tVED+Hao
ynoiXaV8Swg1PHe1qT6MWgcrqmx/1pSr+DCeYWKGIb0yqVGfvQAW3f2fxljK72Fr/KopSrnx6WTD
skChkTIvjlTrZlpdVUnPzGZ3lvYN3WbePXwDxe0W5f59QgvCyLvmf9PUDpckKJjNHxR+p0rycvGg
/JmcnIsdWvBkh45bC065Tn7wqdITvTIYz2wrzKInK6o5fpLi8cs7/Z5ahxRXdhTaKz/p2Aa0Exeu
TzlftlyC+vvHv9hpwF8ys8LG/vFeR2rah6VTyLuRxA8ELiQpEO49wBUYeuYaSRo3j5S3lYjY141k
Cv5bEfGWn9qtF4e8PkxmdHnN9Pm4RJrcKmzp7i3oQIFURwhcSkpivDdc1J5VWijUoZJ9xEbS1KXi
UAl8Nh4QfEwZhAX9ibbqnz2OKNuPzNSks6rDv5NLSunlxSmBSdhncMfZG7QflUNUWue4uUxr1N9Q
7X6S/udNECKGddWVqBlqQB2NfhC05g3tWRPuRsSs02Q0eYbDWTSWWyMaoE1XEyu5I3dnVZWPY4cS
W97QlJ0tjx7rACIfghcZ8c2xGRD+wtkRJbtyQmIKKrJtYb2g8J/wIlBnF8m3iEljgtG9wk0umsgS
/lyx6uvB3aw2M2l4ncbVQyS6Az52HWZNeN65WAClvc3nZh7lIfTRBGzz91Eyn5CLbV5WFAjA33en
XInLTZjkxxOIzYIKSNG9Kqy+dnMmPAjV4HGvxUapaFhBZKn8OleGe9tDWC4xHpObLYCrSmxet4wQ
PD+jQLHl1ey/62hCZWg4aQGRTWATr0jI/Mrz8TXDf1HH4Sfz3MppOXaBPjSF66jlOYseB1/M/tBj
mhms1mBBnrfDDKjUnOtq+w73QSqGPmDauzewvA67bSB2czC8T+B4Tc8rNNLaFIQnQioKuNOiWVie
/p/mWKffJc4uQAjdMOQP/wPjqi1QG1wTJIe5koNmA5oxW57tWf0FyZSKgMTHh8wz/ivELw5WqOi/
RqiLxR7kr/aCZ9KoMlIgueDsjW2UkvwCOJ4k/7Isbyzml/0Sg4umfhyd2KXq+wkmmK/ZqWlkDitM
cnYNeGuLjW6WRXIvQj8rGLFVGA2G/jAxitseVvfS8PjkqftFUp8mivLC6TnVCJ+NQQG8KtiS8Eia
sxyf0Xjl9/4/Wd/YD3X2jSHIH+/auHEqZpotHP4dfRXuJZZSNGqQgcrx5+zLhhKmbYz3QYLB+2Iz
pxW+RIQPsCCPC8jF8g8b2q2a2Z2nhFC8R853bO8WznnqK4pEVGU1n1INsUaWPbu9Y6rEatDWSubQ
rKabix6jbfNxseJtm6Wkk59WgNm6rB/fPzFZzbfqSIyArwbmqSORyrJ9X7EEqn50uExkEyxe7ocG
t/vPIQT48um7ptCL2Iqy6cT9hy9LYPdADvJfvdCxLEgqIQi2Le8sD4rXq5o/UW4IMaNA7v4vbfma
3af6UfnqFao4E3FxCbCRemBT3LNGL6/0dVWsIVvus2YjwwrcXYHw4j2RuE93mN3X52ETx0fss2ku
i+R12ka5PHLVh7Egecr+TXVeXwcQEeKqjM6W/bLaOQCa71zHwGS5AK3vN76nvQZmhI0vBazZ2Eab
UA+NzfTQtK2SLeOa8lHjAJNtY30zOZwgjemDfnnil1B8hBUX7rnOsZ2YdjpY3TDIq51b/UBqNoog
Wi8t9cCgZ+MEDI3GlzG2zh5RustwpqPjxaPERoQBJaBvqaUuurvgcZIvUheTFhaM/qslc44DCCE6
VLcurJa6tVoqgA1YnDcgE+BuXT1iaLQSrNd+i3MRWuZqx8Fy0lYuVT8Ibz4xHHbHxelapDlP90vd
g/3TALkaLyaaA4atknQNIvDaS+s3uVRru3B3D1X9mNN9Cb95rLabTPYSZ55PMTMOT8E2iUVkyGUw
qjkATGj9qEUT6VuvhRgv9tYrr628X/Dba479ucjJeulmAhoLZaKB1MonAJOVKHbNZVIirhFytzFZ
VjmGH81qWTzUOLdakzT0Bnv+EkoUFgIqV7jqywoGxWlYIyOTscnKSsmkg1uq4yI4uw7SrF89ufco
ujKuWqZQVFLyjRHYsb8lnM7CMyP6IAAVqdWgpBj8er24YVrUQZRsXt+eeKUZ4hrKiDx5ZCSAftrg
x1shMMe7gObHmtWFqu+c3NIGONZMtORbSwSJQQxedI91g7zcaGnRF3+mnciwGHWx4J5XBgRc3iIt
TpaqRmX8M7ZlsIuC2d5XzByYbFxlQxpMdqdxeI7la0wP1EqFbdkXNn7mvA09JTisMmRGD9y/tRT1
Fc4pu6cabEpQ/05YiNftGFegNC8tSk4n1S4kUz/yC8iqg/lG598xy5FmPlvIiP3zy5QuzmtKqWE6
tC/ykQvxqCF5mgoUxT3ijBZc6IxyArOQXmGOaxclrReEg3i0D2HM0Avkxzv83gVwqf+3+4CQlf5z
HS4TnaH46IlDE5WAp0XZ+gC4/GRihSI3S9g86J5RqifVampAceT0VBZ1rLXN0gaW5RJRaxaq6CgM
PXSrBzz/m+hQCn43ptu2IK1vVX8y5D0LolCRvjQ/MmmrJcjm0BsPxiSXUWJoxzFRfAWzt0/ayKH3
Eb2A8RZ6F49ZA2f1+6+EP/PC3Zv9ARQLPDlcjeElYy1iFkN7Vp454CJwGWob3q2B/STGZ9AUBOQ5
1Qgk5S7S2vxE6A7B0z6QmdnB/h08nYXdhpzmnUMKvgPQVvpTlJD2EBrCEg7bEAaKcDPVaIuVZWnG
Jls+wcUgbgiNhYLAp5bh5flIE/wNgE1w+v2qbBwQASFlgpSWp2WlW1eMdZcDVvWKDzwEv1AFumTU
0fMVOcUuxb5ebTjdYTRDelCdIb91sVgx/uGvqmaRfyaYVPovLqAwiaiKyrmwyV0NTDRdqLpbDtqc
qYsKU/R+N40d4orYhAcItIVZYZZBi704jaXASqOVq7tJZHKFbFX9BqnAtf5Vu3Tys6k2U9iz8giI
Btqj1TqDO9NKbUdrapiIoyu4ZVxsbVpt8nBemZHu8xdXxdDqHPKoj5O1VgAV2y0Og+Q5W3fub1tN
9E+v2Vk1rLJurVQ6Al66esvtM1HyuFdIbZYXkNuhmGwrD73pdP4jckKNc8rNsqFjjNWXhNzxrDMs
+m895sHdr0aVvip5tnz9DPyKBtgYsZtZGY6k9AGC1W4FSnKqzDBMkiH+xUfZHRxvP71FVBh1HOWx
iliA95EnOCBPAhfFi7ESzRpcgFeLvNvwaRm3TQMmriKefade6s+Pb9Xo5O70jKBeO+aqMMScUX/r
qbvKj7VCWg4EERrAeBdi9bbEjdqWDdHyCG4+4D/jf90MTMEf6it0tER3DD+Hc9MwEC2GYG83Bi12
X8eaXjaJxyR4vK8YaTKFJxv06GxQ13Couv7FJKg3zblhX2fJx9KrbuQ3ZxnFPJCw5RcGf6mJ1hkv
XMjfI6meQJM4JA3b8eUdsbbKFkzMo8wrW29hlW9DaeFsnHdXW6lBjaQ43yJ/XeMRso27k6ZhXBKd
X3uYbiPFJdhlkDAYEmwv4FlX65KSixmp9IsG8yE5Enhlh6J1k71HMVF54qnT9cpRVIEkqHFy0yQr
CyHiSK6Fe13KZ2jP+uaN0nbxetV4BtHqgeKUbjdcMFMCiPZ97gr4poUYcX3BXeQwVx4OU2KBXlCQ
Iq0fRnmh/e839YGUMRbhlIAg3LSTOKnQtrac4YNYpIGeiNIdxftKxqz5NE7CU8tt7x0ydn1VUvsM
W5LB/PDKud1vPVrF9FePBQo7uZ6JZESHqAODpVK/wEvTcKDIN+224KxgCfu3qkh2jyTrIuk9DJ4/
SC/SEFeITzS2BKzMT7kNpx0154EfY3ew+mGqTCypa8m9EEMQHcj6q5NJm4YSnQBW5uF62pLNtKcv
yY3C3DUi1+PunM7znaSq3awQrOhvZVI5trDsoTnGi1ZQpGXNC4WSkvHycVw1KI8T6d1ydOougq2x
X8ElWghWxWrK14gN2c8vHfAeC79UA9BCdeDCreGayKP4w2jIxx29jjTuCNp+U3EP2fioH00lzyWT
YCIPH4/LKVKQgDoeIC8CEtFGM5/dvT8uZVN9mkY+zLduWosi3KmI/WXImqAL1gq47e2yP1sE1Gi1
ggyRnKx8r2jP2WnQZ1NkU+fAp88xeuLk5d0FcoK1wxkvJRNan+uRB4/P04QKVHYzw1DuNWGqG9v5
YUlZYSGousyiGQBC+f6AyPgnxUqWSZuYb2UC36JJ86ce2olmKHRVblFnNJU6xM6Wvzflw7E96I0m
pqPiLEULX/Koet2RpIqem3fq8jyXBjYy8NqRbRXvkiEuOeUWKUV995VO2dptun08in+/Nb2s/jDU
rNfdyVgrjDDDu85tkvLv5s4eWnJRaeqn2N5rdsfskRa7sMkG4ljduG65CUs/RmXYotSGP/q1Ym5v
7GLFTnXmP9gHPWF2Erl6wqGvip6mfJIJ3JLGpofutVY4U6VY/ePl71izfdFugR/m8Az/Yt1fhrsP
eQBqs9z6ee9lLcrdBQVLbirgr7ADVazn91pUVFyXzH3NQcaIymcVHbDDftVRv7WljNtWZIrDDghp
STh0cEqiGLaBDin3r2b76p1kQNmkv9NmTWt36/iHtiVdDJ5zMKVb8OYYxh29He9nbp1qEi7tAxD/
z+SMD2zaPdqmnzL0Sx5tGq6nHfGcbhJOnfX6SWeqOZ3Wo5OVyaG+Xyx0RvKn1vaHRPpusiqgBbuV
YEo6vSclmCyl0NeiNoBozhhZnKVUB/JfONNLdfkq6YhF78CfqCdWOp//Ct5tVeJvVor9iQOmG3wR
WSEUtXVTPmK1Sza0sN57Z84CjK+zX+mCSvigc8fA7k05/EhU0yjzAq0CWHu+Ii+Egu/7rl7igxYT
F11i50uyAbwweCkClw8q+A4llO33OEvZU91Liq64LZw+qgA7GPlBCtgrvB0E2W7VJUptldfi+3pC
zE035/nTkLmIuFifHLia0N4OfReM/DEkPYhVJhE2IDhm+0VbU56zpilp+xih994oZCsFHqe4sp8h
rKpOwFxG4IYJijtyWMiQsZpl+I/Ypz1WvtkRY3LjKZhm9TGLR/0QHRxvgPmF1EVC2kgGBgNvpN4Y
YbPV7fco4nA+JBzcn2+IBBlycD1m1JTVFURnQOFhGjzBSEwURiEqKKlF4J/ged36RurlneDXcTQI
PjqICPsJELyt3pKDbVQzhjWaEkUbrdk4r8pmWzEa3YLnlSZ/dvPUr5DGlBgqtkoNc1eUVOwYJAJa
P8/NJylHm5hYc3zBWwvo+brH2TIlhWzerJkPYM/wMNjPdBQdJZtt7Hyi9DetR1AiEx01u5SyNnu7
Pa245c5rnyxZLXt1NM8tZTCidn1FwCy5VjpCIKvVFEARMoQ50D44Q8GoXERAY0x8y38p0xPd4pHa
my3Y/sgYfYIfInQ27LId6rlHYxRf0FmMW+/NfOXUDuiuwoLjc4uB7ZltDvot8pRwUbCw5FDRlLlF
6LwvFNZh94PyNnf7pLEWCsv3dZDszYVtMRasvVR8LIt7jaDY3y/yRq8ZY2eLzh6gBFUyzbt1bN4c
j29zsTQpHNiccw1ntoKKuTzsA4hSrONzOtw9J67o8P8KC999bVbcB1axQncWa1j0xuaj16LEM9cm
FRYMeJLmc93HH87XnAo7UHwUQ4XZ6JH4/q9px+q9kUjdZ9JOqtgRr+NELoNTnStEXmGsml4cik1I
CGnNPZBz/31psbgALjkxddhqnYH/sQmmLpaZeBkdrmc5qSSjSS88zUlL955yfP69pH3JQzsgWLW5
aIAIeyL+6q1j3/p16aW2LyR8VrwQxEnik4v4wnhYZ5iOSSRcwvZruDi/xcwWdftwp+v9lzH9fVSG
VujU2Im+dYMqt4HU00RaivQOvOQPoMZFz67g18eg7k72eIL4z/ePQRAkNLkjq9v+uBHV3vl5uJcW
SAn4zYgz4UAoTdsGgSF73XpDy8W3guwyoordpuDHd1sQnOvgQIlEV1FjUUr3B1MUVq7dwJL04H4I
e7bWDgirMedbxwoEMuDHLIVHbwmf7BoChuPChYL6krAkhjAlaOqT0+xAHFwMlE9xMmtMnJwnjK0C
6FuTIGiCa7FSfxq3+bsQgsVj5fe3EJYRsw2pEt5gB7j4Ruwt/rADp7SVqrgtpzF04H14hzzueNt8
oWXjAEScG2Xl4S0bo/Ftls96nOYubawQpyIzDEjf6hiBKzRIADzjhOtZaSF7NhAn3j3avYvobJ3m
6dDy37NXFxVO+l0MasSPcwoUzrmXG9spZcFhnkdvlqPr8Z6z0LTCs6KNAIIgrn8jwZQlr2v+HOZU
VF+uzO7KUdYTkXb6A4bMsadHloJmPDhHVNPDUqaaf9ndhc/MqTP4z2lKm+3VO2wv/w3SNZJmqyNw
NUTLmBbMlPHEMyn71iRFfvgaCfDqwcAwnTNrZlG7m+zDH5Tf1shTzshVgEyB8VMAZPJ7iz4w+xHB
eN7tfKvKcnimZ4N2RNRGF7/QrXFKMRvcLnIBC6f3xReVHYLFeQnheNHluxWxwhr9tKfhGu2l5KyP
pkZ7rRtdmHg0aPUnA7ov5xocSFvLsuA3S9kZkpKv9SgYTjCOETqSEithyu4dobtm3JeRZyt4yB9w
7ITiM1Nsrs3noRhXD/7UdJKbxiqjPaVkN4N0Fd4bvucRxJ28iegClHEfmROGSPoYMdlD6lQTrW3F
4s40Judb4EeDqssvhDonVv2PnLdPZEr5wWLzK6othLS1HcAeQ1x5QlW3sIus1KCDEgeSFVORUSjv
Embry9xvE6zsUKuB3nv3Twx90qJW+rQvTIhScvew6OcBeWbHbpD6SLRXuKUIkBra5vRXlsZHz/XT
HtzIkKY0j0jooG85Y122UP7tNUFglAaBUK+XrxxxP74a70W0X4z4HqeNOytptaPywk2OUfqe/SU1
X5NbC6BjZLfqaASUe9pO1hMgODn8bXGi6RNTSm7OSMi99eZrR9rXEg3eBnVqdZVLKGRqul95GbrX
YJb0pRqCLwUj2GotWW8LLPwiGLqDTISD2E/2lXFfs2JlhGfGFEOCk39nEAiZ664CTLf4etbnXJzF
7FRevVxOOsegYZo4zasZEc/um9JzK1qvnEYX6mcpFSu0FO2klZPGxocYzw4UFc43ngX+L4Dxzelw
xQYI1amMmB7XS1RdKAt5gkNntZVsyylD4L1PujLCt7vdIjWnBwzxSh3J8mJLt7wSf9nyQrge1JCl
d8HNBeWOtBIHFz8IAYhWfBjOeQbXuIsV+Z3bSH2iKm0N3SYLDTFMTaufiICaWDV327GT7qmUD+RU
3ulyw7riVUTpg5UzhWED7jeRc9ZxNX8gn+1GeL37Ip1J+p6XJ+sHpKiWq9LQkrshtGUvqKdPDhAf
45Grj1Quntwobqky60b48Unn+5hdinco/zGFygGFx0kvyO+QTeo/zVxULOGNCFJSF1fwQwZUt6fP
KZBeJzRgCXABxug6QQh4rJrgOJJMsfc+88rts2eeaPsT7C49vyvOaTiemxb8jtSY/opystGmELSu
xQOBnSrYS1BXxp9iyMy2hSBSmc06OyFV2t4zXs6DTYwDtOby180GxBvOe1+ivTKZY/V+CcV4gC71
WlUFaz05Oy44TYY2l2wBZ65eKZOts74USwrCYSQ9wIBVfti+uy5PriKNsrY0o+ozNJQcQhpL0/uc
o93RyhKI1mbWGVJyTm1tpSXilb56D1LK3HtzIDG7KNZkUCCnT2hIZIfrtDt+D6x0tTL/UfGVFz8Y
61eUhHza+n291WHjBj+7CuKlmHKAcPtQ853490GaBD20Xkt0q8SD3Cyh51lliKXBtpuqyowPK3yV
J4J4Xt0yKRWDWV9iK826FB3bGneh3KA7JRnMC57rdm98pFIud11sNSFhCARiXfD5K1nBjrVJFF3U
bOhNRYPhNN7uyUI6HLw7cwa2FvPji2bPl8QeTlBKS5PvEx2I08v/mefd1ge0wsHTzZl2yVStDXOQ
GOW8t4PQX1hhMTiSa6rocWdaE7FEYb+VwYWv16HRdrREdr/HpQz/4FeftLeGCdXw3TXgR44bGD2a
fq3Fx7bx7EFP2C4Yy7MlRTD5TeI21u2dq85myk3TCdh4Ra6rd3i0CNmNZc4C6oHiWgwE+SCZ2k24
k2OcPPsS8ZOFp6/xf9J0OMtnHBbV6KMcu4eYK8OMsH62E0Q4w28Yqn4dd4e6mfv8ANwHp9gf5mdg
p7UyDcQsOaHqiNNmV/LmZJ/uDS195WNnmiTSeNViZK5g9D5DhDsa1qz9hicU74U22AZhX/I3bHEG
4h0qlMZ4CKqJ+bMxNK9IydAGL8caYi0XbOr25NBbwd2pxIYI/ppEuzNiMnFuuzJNa3Nk2IIzbfgH
FjreIbUDJhIwZfL885a0MgwOxzHbUVWUdSLnfbKJkgU/g00OTGCrPgJAtnAavAwSBQZKvGQu94G8
1TXmOqDa3vssd9i4OXp7mS9XcMFakrQxKTqsdAu0Wmga0MekTL+GbjE04u5BAZzds/hYnN3GJOva
mvsEWdQe6IN3MVZ091DjIojQonDkbkBzu1LlJ1oHlwVfPKlh2nSioGV00ReYXfWX83cRxhANMVca
pmOU0EDZR7RPY4Ak1iGCYR1z8+xAvneZUFC+UsG3eODtksz2CQj55EFliRT1/n9SieWalszwTzGP
32PMRJOl7a8rzPU3P/r0h5LOw+2mm9r1Y2qbOHkD031tDu6Khgf6ATbxdfFXk+46hVdOzo+L8ets
3415QDtAw6PB2Ctgj/ZV003UAELFE3/5oQHqlijRY/8DqQ1vGlBw40eefwS71Ah3GldqrzQeYs8G
L1Ixi8I3d4vbajfk048qnJtQdKRk6XrJ2MnO16QJxjmWt+PqQSQ+RNB9uJTR9JxG+nS/YRnwNeVL
akAvthgMtOhRCC8t7Sp4o/ymmdliMr5NKNJUwJFQ+kUFFbDWHGHcahiqD0Ul+calMPrGFfipMKCC
K4pjIXGGhGyIJmUcxZYUMLzx+SAr6z8ra4U6IDMGKbEVGetj5lCAYaB5o7NTCb65sPKfy7vJ8bLK
ohgFtioaHcJmf8XJ1GdJTMSpIWt5zdjckFf0PwpwxF6mWcLKiERr8t0fpr0PwI94c7wXnmJlxzu5
B3PAY96O9sW2XVpYLo+9IJc7u0nQMkDUeYvXW7rEarDQg2ORKVqAEhFpfwSLEi7WLfduXrtlMhYn
YXwzlWNRPdBPx0R5C/vOwWYhEKCdI0jeP2bypbe/fNIe254l3POKvoJq/I8aM6RH29Kc9iE8aqhe
VcQz+T3KwdlkEo4t72dY4f+VDICnwy+y+EExsK/Eugq2pflyuEjHDpvcFmtZlq6wC6ODCKXKzV1p
GQbEPt8uubN60bgIVmLwGqFMW4SUiBYm0oVTVjB8YsDKpJ08CTYHWjy2RL9qaapFU717d8acb7sl
BpfDYgROv1wtHzuHv+2XNNUo13u/BH97NcK1Gh7MfJaktbpbTHqYyJZ0iRZAXhd7pOh2TE54zItd
1LfrUyM53JOIKueOJXQhu3eIYY3olQeoA+wIfRY0oPnEmf97GkLjNW+/GyyfrC6M/uqhCMgwqgFW
1iBp0jWBpOUatRDpxy5Lk8SWSX9nIIVuM/q1nXTFRiiGueAJWVufrYviDzJpIqZQgxpU3fnj/K+L
BEE0KZ2ueu/drsbv+kH4mzZM4nUG4iWxGpsECPt6ExP7A7+p1OzrTrMKmB3yUy1bgVy5fzWbNVmj
0136g9N2+vTNr0G1ALcO4rfSAI4/LNlx/OKKacn0TcawTueYEVKsSwl6VxXwhbhT9mqKPXW9RMqv
kOGMRQPpuq8J+ia+BdU+Ib9i60pqjnck5rNwYc6bGByMBVbsqVzKUljy7VSJQsxn4IwA2MoQBp+2
Nis1T2sloFtF6Xj3ysd3T/Lktl7o4lHGeeaTOVa0T60xN2SF3b+95NfUSvZavzb/hVr3/B2yufnJ
ZNG88tN7lH+Up4Bv45d9x67kGUlqq7zGyeAkc2w3Mq5tQZ+sJUNtXKv8CZVLLdc2cTKtGpWkADZw
hNmZS6UV9P5pDDdEC5NJNmsvjc2XdMBW7FHfjSRkBt2gQ8dz6bknnUD7riRc7+FUQb7mTjjNrBCV
skxIJ8Qq8VxmxqRQGKA1U0e9sdh7QmS0KQRTXXGyU/H9LqRs84Q+8Gd94VBs4Tu/ekCNORC2yS98
bcPa+vgi1NAK86lyEjnf7hZTQKN3BV6Paez0Wm9qX+bUsup4KGiU7q3w/mIUDloGBdcCWBDTmGDQ
Z1HRgexFoO2NdTjYhCE3Py5f6oIYw829zY4dbK06QvYvUZ+IJ+zkaPYBIbdw0xkERkazzre9o7J4
GVsJsgIyeu900YyUSZJ+vIUi730luveK1qGC+27q4DD+aMoi1G6d/A7VgYo31FZ7YD/3iB1YkCP5
nSUcXReypsS99BuVSjFM5j5yPpc92b0jEjypmweIOmUv2RP40pYW+mdZOkKuv3iIPrZELvftOQDF
eCgONnSOdI2M1EzRumt0mCmAI+yk6o3CDdIRa4u2sCgyTG6M3c2ro7g7OL7pEpkD+8Xw22cfG8OE
6Uxp+jFDgFA4Q3BBD2E3cDhwVV+fUp7GRp/8jDQynn/ihSWJq+VoJqXlRKI/TXcPAfjCsF3ZR5Ug
bimfDgvCzSEh8HhwklifRn/AIhR+btRaUaMj/R90bxfGKuRfQGIs4Yru1SkwWtnRLnhjyKZS46rE
keo9jnQNKuZk2M8X4vLyKJh1Y7CQCsQxLsTtRibunrqhhfLJuajVy13WzNc1rnnsPB6ZYnE3p9i7
vsQfSWgGkRjO6fphnZpOd1GxcJdicVwrHQ8smFf+pyQ1bQ++dVltpaeRCoFF5G7Ft+4XOR3xA1Ni
w0S/zdzaZrcgzrXuYeJFKvKZEhLydt8W9/13OdoPeGkjTmRt9DqoLDDwLDu9FFQduc1oNqp9E2vK
o7+NINnI9TxIq6HdItkhP5Zqh7nf9mYLwoJAkm8GqIjX3MoBHvQE/gowuYDckvKsBETWd7tJZnWh
9vjqQf76z2N90GbvSkgEVruhFsq+5xiAYtCXcL/v6bYlgAsmNS9eKomOHGFVWX8tfM1PlAq3nmkx
2xR+uWMG7P+W/AOwxhQH73ubqqDkeg8qzJ/uFpdZ9iZbfluL2tU931SslA0K8J7GYLxbHGpReBic
9J5itpCaWp3ktvHwpBr+ke3F6iV1OV+0mbK+wjIHkqGtoebdqK62LYNyadTB67IxeKE99Trc3vYT
HHw5p675ifE8dvlerZAWd13syBB3am/WZlEdFefYGhf6Ke+Pd2cksy8WEdAEiWzRdupYEIkQTka8
zhlb9P656dogOKhCVsZQLE796GerUevgVgcmVBJYHoh3WHhRhKVlkYIMyTEip2g1HezakjVcML9e
Uf2P+D2jWeeDjo9A+l+zTwGBkXF0UyWk/jc9xAsrbq66+zPD0ekcvBoUJDChWPh2fCO5gxdkr8Gu
4zLKeuklE+8bSJ8Fb7XwhNVRhrekFjRbO2qIyFNAsYY/AAJKXCHDrgyLFGd5QBXBkXr01eU95282
w8Qiwx4ebrwDLjD1UPAo95hbzPlBAO7bEH+KLaDG05z5fnu0lcKS4vIOSBK/q0JfO/FgFyyqALDV
azQPERJvEJS/i5PILOmUZekjZhf4DN1TKJc3Przf68Gd77KH2Rt0u366NlsrAlhZSxOiYgy+ZzaJ
nDCigaMcoOUvl66t3ZwRfQfV2g0/jD594mN/Fuvalxa2wAshT4+X63v1rU13LJ8QV4MWLnzSNaHG
lqwaqIdddoSFr07DDshhome/cLEGBmZcGkZQbC9vCeU1PI37wYOdkMIAVguhaM1l8Xg7swetOTa5
htnadR8Xv+yhl2SpK4JDyBxqt+bsBJDVq3y7UXq/JcrOCsgSUJn/g/mSOKn2ftUGOLCU3ZMIS6TI
mLqX5kJgYZR3U6l0nJEB4I6Oyr+0K7peadTgp/5IQIHlEZytAAK2Yc5/D1sYH6s0SCYbp+PN3G9c
+G7tVL2ENY6F9zriui4nB7AGmOJHRR2RY8b3lYLBLJ480lDljqX/87qXiNdEFBuRs6KOsoiD0pfH
ZA2fLHh+MkP7B1cwvbppzSXRHxGNMpDPloxckDWAG95RIclPtrSox3Iy6ttqGvWFn07ee1rc2tSv
q9BVXZGhOI1joA+6JwugVSxzDQlRFwPC5LgsmRAnXLenn2rQtb9eOlVXPSCQvDDDk2I5yIE7nkUE
yzF3J762shjWp+EGDElSeNf8I7+HTNmUP5kfUUnfKyIgJOUaPBxGYBsyTgJue6Ehr5r19iZzWAb+
p4oYjJRcBthPPA49jun06ecB2mkT9PYDgJGMn972kj7h0aMQw+15pBByWjYUddOgtd/tgOIVkQbp
bH+rzRHLA0Mf68z3T/dtS83OklMKC/zqEMQlL/zBfPiJ3uCt2iTYoQjQwz7poGqA7+Ij9jK31r63
U+p56qOovvxckGm4qwLPCm0XErTGK3GRbAqkYOmcE7OIe1P04YLEpn4s7yD78/HzR+X14UEKABc2
0v9C36koCveCzUOvDKlAd0f0fBfirfgA2hRvUu/epFlwoaUUXir4M8cgcwi5hwWsanvkjJmx2T41
MlvT0Uid42x+UySMkCtkYQy6slR0yNexuiVW9o0fuV0loBpsiQJnHuQRRs7X+DjarP7evoHI04st
Kc34Kg4dlf4r9fD/9CDjzox5E8K+FdgECPa3r0eXxrbhJKNGiG4XnrK2F/tFXAu/xEpzDbXYPYyv
Y1AY1rr13HZcOCmAUaiMr1TyUBJr0Fl3/C26d/9f0bG/a0wmLB2YTXoY7Qv5GZT6bzyFYVUXZn22
lsYqt8LQwb3oVFC7JcdsnD7WE7CHnSfntfUx0uQpX9dw/tkgB+Z388AitmmUvEeH/z5QWEj3aeMf
evT/2nA6ncitffS8pF9kX3K6GljLIE5GGLySg/a3WDIwpJ3ii4xcnrr6fUGEq0ad+vXVsFgZqAWa
9Qq3/KqFGuqsxz+v/bIDbMQ7oK1PXsXCcpLCBNOobSqs1YOKNdZQ0s45GT4MlMDZJIIvPiBmLFuk
kfO7Cw9ZlTHucJ70m+S1gY5oEHx0dBQTeCMzh9RKNSZspuJScpNZrEndqxJqfeV3WFkLc3nQNswH
vp3U3FTNz0Eg+U2f2Etyiee3VTHqm8u2h3mIZ2i4Giq1AGXGZv8F3evurm3rsV/HF4hks7UIrPX0
wh35/1UJF/ZjQilCvz/BE2FzFeJL/s+eAi5skUnxXanNVwhShpR+0TsPnR7RYRdEh06JBfg+NCRa
69mo++xYBgfEXl0R/WkNH63dLhlkjissbClbknX8NYN3nxwGVFJVU9fBUIIU/e4UtE1wSAj6F3o3
5Y60S5mUkMTSpc14EoqbiXwtE2aSKqbWe173RxqJlBFE25laUj4hsvCy3CSaex19Q7wN1RTgKK55
ljUOotzu+0MiwgDDYGSevLK2167G1TLLCzfn6LqcyC02ge9dWTw4i9WqIcDbZ8iCyRplzE58sVt/
j7tS3FvBPXsfoBBVR25FXLQ9rppmL9WvbI7ibMYjpYnkMKvgne6IgW+lpQBUC65isat/tAO95/j7
AgNkBCxzFpW/QCn/qhmO2vjzqKK8Oi0OUr1zH0caT8vrBKvdQgTEaiVDulyFrpxZBxA7kmPnwZZd
jlzJsHKp7IG0lZi4K8PdFl9Yez4kqbXp8TplgqbChFeHyS/97hzTSqnvlTrAtPnZEsIf8wZgqmrS
db2Cn5f4rWiQXYuYTbOWDvdlXrjFj0lTYlItgTFRXv0pB7b/1HXxqFeVJgbH0PubOQvqL8gHwS/f
7lMvH+VlhgTmJtPqlJlYuR7TIvnQALNYW/47xtF29Q2aHcPkzVJqyvA+1RxzxRPcQuo0uNlUivrG
lL8428Zv3JUdWaFLqu3au3b7mWgIalMH5i7hERpBIAMFRX2G6/9KicY1OdSXvs0uRlEA6sqBFtmB
sqmj3kTZt3oZjrm/xTW2GwZeMuLarwGieSjAGjSWuc6RnxU5XpnUEXTH6A/TqcCZzp5rNtgJY4Zl
h7UsjMfWyouVc1QCPC35OsggBS2NHZ6dDUe6914OdIn0mcB+zizhwMct4RhcOVnefEufWMctM5uD
/jPgFEab8RFM64DCY9T3SwC19ih2RBKgW8YzlgIsvVzThHYtOhPnyUAJD/n+vNg8aGmm86wUWGqf
U4NvBvkW0w60TxyUaJI/H/bdj3Ri2yOKrZXthe64rOuSrfGly8JGjJfSLsWwcSSf5/fmu6rxs80y
JYSw9FT2vsweGnpxAO2LNen1lizFmNxP+OIOGT9OmPLZLhsK/3baWDjpRsmoFR/V5q6s5Ye8pbn1
OtdEIUc454kGMOUYHCE9s8tAkbC5WIxplwNL6GE2jyzmAhjxUt9R/dduPyy9z1VjJ5tO3VdBAn5G
t9kUHdQ95o9yB5O+KWizNQoyWAzpqWOMxhBbhMQjRPxpWHxNbmTlIYcsl9Zb5T7A8c3xEZnDGmyJ
e/NnlTIiX7aAK+2k8Sc+nI01yeTxzmFDbM2K03eQ8SOUtH9D+zAUK6bfqTSuUwXFhBRX8NlXEqdh
8rzU0+83UBSleBp0+6FJVY12zKBZBBVXMvzwFyo2aLXy7BFjNAu5XEJtxGZq8h/tSKsAs8aTC7MD
2m+yxF9zD5Bh9h4fUfYCHPq5uaFRYdYwN0FCCrI3G5Awkp59qYMclTVp8oiseEesHq93oJqG83Wd
Pi7LDRoHAb/BHJFT6q72PVqbB5sy0M60BX0cTS7NXFHQkh+xbIOnOtSYgd3La17Gl7iQ9Nk4ZE0F
QrE8o0cn6XN+yyJakL6ztqOkXLuGYpQG/oX0xx8GC6mTQE8JUOR7z2hBSPZqvFaJ+RKvThdWfErm
/l+bfYzEo1sdoR/tT4TgrxNh6DqRooQZkNroin4DMs1igesIiD2ubLFch2z8+Fe0hGi3POYEeqOj
w64digKutwzsOSIH66ILp8FsvllXn3WCIoUE163nSneX+RW5kZcmhGpRIl7F17HJX17AZfCIwRPG
e1M2GZ93XH1iNn6w/qKRsbTYXtSt3gXVONk0Oe48zjbiVflktihuOkJh2lFr6Mwy1HDorBGVKPmk
U7ILg41AxSbehk2pXb4GjncGIAOch4lL9+hgj6ctwrJi1eEdkTcUOjF4AaH1hQDUIkdLB8RaXld5
HYfS/N5a3k4HtLHddNXOKUgLFnsO3otov459+OhOrIvsR9UHt9lxbs85d6NrP84wkvIrUTtiv7Le
y0+MMsb16ADKTwbV/1pDds5F2BThWxYs64c2QRgFbIhR1NLB1itvKboc/+7eKtEb1cNuMWUFOXUx
UdP7brrqOB5n6X0WJv0DHMJmQHG0ae/dRfmS6a57Za5cT9YBZymKLs/UezbGfpNcENX5jKUATQ9d
AcE0mah2WzTUqFZ3XowZRpP3a0eGw9V9IIJtK6be0OHfKiOTVKAdJvAvyUxODkJkC07sSZ+Nl7Fx
D7SZqiV0CsN4CBNbgNIM0EjTJFv1M0I5vqj6+tXd3VFRQOtnTv3dCZvxCnjnYNxNf9tlMUUibrpc
FTGBsFrZP4g9I1jejyYjHbqJwQGNq94EESmXBw1XmfTbvASc3I2R7wCycwVfL7oYOQAjHI6MY+jl
TeZMPkXnOPWQEAGdsqd2qDnHEpzdUXYeNC0plHF/iUU7vjOjmQR4Yo73a6Rs+CyWPXfwly2UsBLq
q4HOaq87Kw9cG5o6iIW7Utbce5DW3uz4V9oKMERf2+1L6SDNvmOtBk3bdWHBwPJh5ZfVn/Sc7WlX
s3rUIlNQHUjCduUu3VdKjY5KVV6+rmYFbvuHIUvtr0md6Lcri7pwf8g4O+QooNTmtGIr5JuQKh6o
jAeD2JSZ+HhhxSmCBx3ERdJ3wTg4P+E5rB4xj7VDrVu+kzK7tRdVo7JTWDLBMzV6BI/vCiUAr4X/
bhKYXDh+RKhM9jpc9X3TCUylGYi9U5ymbDaMkyR8rZJ+iviT1dChqpaRbWR62P+ILwE0do+OY9bX
6bmC5NXhncPXhqokaEow8PeNcv8AohBHyotsiIFK0e6bCF6vgCwrfGQfQx8u0w0ew337Z7htujL2
J0x+58duJPbss8Scav1BBscsAHaamVQs0mFxE9rbtPs+9ZBId7VfBPFT+ehfppkW3nCelm6t3/ar
gp6MF7V/PhYo9NDFQLdGzfjLBBNQkst0Mde+iF7KchstRl1gN8FXwfFgM9uQ+B5u5ZsN2up1kiQK
n3oyoYu108fsnb6SYYw7/GkxNmLKD5v72kPEmObl3KyUHuepuK8uxgDft9k6iCZvJm3vp/0/lye8
s+ZlAOGwJuDO7jLtj7g+u16DuLp+4dEZOHZz+oRrT1lKL/ZAd12czvoQPlQPJf+CwtrV4nh1VVdM
DR+5IRkyDn9uWtmxBvt+9niXb3hCCiXJJ98OcF8rartQvmhc1OZa0Kh26JkST1sA0ihmyJAFIixk
QETmrHxvviQqxy4rpqgeckgSzAvjO5I+kAHxumWbnT6FLy4YFamnLb59iNymaN8Af0EFRxbKwIAq
bBMXlHNB0T6MhzBwNRIT0gbVRB7EmtlSXgiOImmPGWsKfH4aE+IXlCrRF75jLKoOuEaq5Ro4Yy5q
KYulcdkroMEnoxEsm1bsM+EPv54M4xkvjq0VV403ehTnljD2mIlzG0yyLmvKpdYAcjFVF5SoWBP1
OcgRoPEG8KqpNAfykXgG07QKAENbR+o8fxPabVvMp/RIDtSyMbLRp1llgYAVHDD5vcs4DK752+PS
Ux8vj/MQSstKv5pySy69GqQ1+wHCIArKOP/+l5amrvW2Ojzft3n3l1QZXWhUzWyMWkAoTYkb+EyK
1m++33b5Qt2FXM4QY7eSoYH8oFQ4EiwiApR1bqt4X2V1qdHL6B7A8xnZTb5dIN9BAwGINSsTmIMm
CBdykmkI5X+29FK7uHdABpcktrALobhyv5GJPdTZzHbXYRGaA14PgGGrkzTmKD6OcHrJdnKQF4aK
3gDe4wZ+/JEt7ZLX+GbFxawkcEwWHGyAtVa3nt6d3/geCIFYLIt7VqAq6m00YiHIjzW66f1oAw7g
Hm2WmvBK6HmvC7VfWpeYBiEW1NKTsM8w/bDt899mRUJ9tIKB6q3g1aiwQoJ+eJYjtHy1rLk4p/8A
pLeRCzOxv86RpRrw3FBm9r+63M5L0OSH+SgezkqtxEYCKgFvOQazg0g+RF1fiNHuQNu8KwWRkw7m
l7mjRwNeVAPf0w5zkN+7rfR6EpMKhT44w3Y5GurYl9UfylhghLIG+GYJZxgqiA614QdNTGUSwaXJ
l0JRDunuwle2JaUzAvuQJJ3aJ8kLce+wZCMyuDuXr69QOn0lVmTkWxU/KVz49BB43c/fVhAWNWQU
EZ9UF8XQL8J+zodMFM8fj2+22atfzlTHkw1Ez4uInfkHS+SdqYxfuqqtBAgOMtCs0/H/fBcLTvYO
swFMT4Yu5CodXu9DTzM6YsWKxBUv6SKfOVowJjBZePgrv7U2JxwbkcBywtD+5MmPr7hUSwgXITKF
eWIqFtMKodD4AQoY0Ff5544cTNxI8Mb68d00XwVSveEoSrmDmSCR+jYL38GFChmd4QmhgW74sAuz
Ch2pzFg8TLmPU4QggoXwE+UNoW9EJprYLRCQ2xFJSs+LPH+VhO2Itnb+yzpJwbXLR7+zia6XQoFb
4ezP5ZDWFbMtQqj6owpaEO0bCAvqxU2v39tw75fZYP6G31djdGz/1s9jfLQE99yJPQFRLxwqSKxQ
QLjal8RLNGkKfIE3bWwJt9Ww5X8tGtOyW6bpddO64jfPKqo/05wchHKpczyW7nE3bo/31MwPGXZM
O5E5Y5iLjSSEufVbP9u6DljxcWNDhIPoBfBH9NikYXhKSnLzYTcK4gSlMNY2ZZ0QOCG93GabhuUB
WqJpJ83/yV2/LeXnXG2kKHGI+WXhwsOO5Nwn7HZVHzNuHOCAlQJS66cjEGTcRj8XS0gya6S58b0E
K6jzUhClmdWXAJGTkOVaq86etTTN+WRzkrKHaSEsDQxmWIB0jdt2Lfhjik5xCG2yRVXnQ3z/ZcDT
RyeUAt1HUo92rP9ZHznufExJ3RHcb7r8a2j4Il5hpDaej5iFjzTkF1Te7R875zA/SonJIp0++3oz
S05sbXq/thGtNXt3xk2+9WIIZ0vHPGUYeHgPPULZSD4inTFWXM1GF1xs4vnN6Ag3dfiuPXrnV23E
ypYtTo63EbtiQ8qryuBIgtnYFCca/asN+FtQsb1bRm73GRlul50oshyA1YYOgRYcTWP+U46ikL5o
pVsxP6sxigb6NqGw/gfxZEMT1KyNROz0mniCO/vKO/Z06oepFwgotrLn2rk9foshTVB0bg0zg6SB
3e4ANYsPXDIiVUmmPs4wvomeSG2xT5zV0wEVfoivlh9/app2pZbht6c66w2dyQ6rQf1bSSjS0fhJ
7W+K6WaSaiu3ul1TqC76c3rQSnZvPBbZO8oJ9ajvciUcpjehRvf5RaD0dMKQsz2Gvdgy+vk6zOqv
UkOH7BSSOI+sJ0QUXA1s30goXmZFICSiuwUGsyHsalzSeet3P5IZpYuxsCtnm6A710pYxUcBVRz8
R1JjRRvevgFbm+TQzaR/y1Zq7rYPN8vab8duoAb4hO5GAEbOXdaNnj4li09wcNi+lsgQvm5x5QtT
BPy2EaBkKYavwFxeeYkd1GUUi23nuSxdPdiBTMd5dQr/sStj/w6lkNwTHC9O3s2tWyPV5azsV/RC
xHqJw1olEs+ehJwtFyrzkA84H9YnqovDP1jVM731NspvpEU3JXlYqJvjn3Co0Zu4woikfaQL5GAx
QAt0+uR+9CfvIGVK9Nl7Q6hJa3ibgJvjGeZ1MPe7t8L+OIebKNJNzlJHXB/ItLF0MzOh/64VIEMu
oDLwVzOO3Lro5KumLEzHR0kKvGujFF2N3DOil+3iBH1Xe6+n3+XnMu7sLjQP7EwX++3cXLYHCVD8
zi5CHq4qRbPyHyctKJ7Dtf/UTj1lYPfS2x2qZJyWP11v5SBiRPNQjs+owKW32Fi2aII9MxuGBCs8
VUgVHHEhhOyezPNGHajePh09t6B2ou+sDdHTgnFS8Yd6cjyOBQMc78MJQ41cBrgC1IAraU65pkUa
eblfaCDKuymkxx+4dtfkuFr3hsOEE1DAIOGCHzJ7WErLgkMCt8jyavJ2Q1KojFMew4Sd/AdZXJuh
pYT0aSplQC+IZWe0OydLZL5N6gdGrbfjpDqd3luapBH7JR+HK0/lTWigyl7EBrzwbmkDy4T05Qj1
ArjSklezraN6tJsJteuQGtTdCCS1keh0z8349LvZNTpkCB9pUJjrlV8HGaj1VOv78IPEdPzv/T9/
ibxmf/xmVABnrD+MzEM4JSa9toAd8d+ohYP+1HuXMwoFeh3xhhXbN+zTTbKtXOZFSN5jFhtihAr1
gNPgVfl4CQ7S1f/158d6X/6PecY+GyC7uTc4vEmv6Vd2f4X99Polxr7Tp8SayGjVd/Y0N7jLv6Qw
qXngvXa32nm74LG9ZhOl6JWJ8wSRF5FcbTPCsYk4/Gq95jhgPy8iE+mZ1xciyuGTAe09j9Vj5/pN
4rPiR7LNzrue77culMmDua9HQFDNqKgMQekDfyZCKvcYDH6WUy6fAFRtN0xBu9/sfW+E4R4mzaWa
t6Zs7wC2h4BHeZCLCj6y44HwNcFvfV/Lm+HI+O2fW1HK9abtJG/FI/0PU9hCUfgWRj03v1HNuM8t
bzOhyXn3GbCxCpbKDwWa2UX8zOiSoXmvhpDiPGNRaEBdseH5xAYLFdNk1Bl2t77iCczT4yPmnnTZ
n29+zf9nQugAa+kZgvQ8Knu8t894Ged/N0Btuwnh8OWILuHarS/XidyLkTC5y5QP5hfjla9x0c8E
g6Hk3IwnmYC0tYWNkFkjwCHembTAKJDxoY/ngtFyPawRAk2qQDmX8VobmzdpyDSZHbcMOjmiEVwD
sAW75hbIHT66CZTcEgpVZCz3juStQmzPwfDEcW4Vuo+If11XEHBKJ9mVy0iUZoaqTPa8r9+kLevO
Ugq1HhmnE5AAgkWXhghTQzv+CzJPM0OxNG1pNOl5HiBzbZ11xti56M10j12PT1kmBLuXXeW/vzY2
Qai0xVQaiwUdji5WaBhQ6vnHw8QyPQGNk8kT8g2B/qgnpF9hjINPoTTrxBzXX0lL/7D/7U4B1AUD
d+NczRiO/annXi0oyjUc4avpU9nLwrjEZ519xTmmmwNZw7T8cOKfFab52BvzjoBgL+mwzU29EMW/
9CAKz1m6gfvepSDDN7tBjWf5nZxf5WOZVQ6wqUTVK6IteTgElg4z+ETaXC8xuHtHNMWcMbnMDmWC
Z2jl4B8jhTOv2MKZgcL+PBZ33O5OJOnQuToZfAi+C77FSnB4ttyeRlYab31ccDGgYWGichkwIfG6
ew0/fVusyXUgORLXUNoUF5FdmzDkLXWre5TrVec3BxaePr7/9PX1tSyu12vRontnO/TZXaMleFpi
8XIziDiH2BEUZKC4JIw3SBexxSv6DJt3pHov0xH8QwXNttudRDXwJ2V/qjat/bLy9YAm5acGC1Y2
c5JgzUF1hJ42+eAeHQSTyR7TR1Ah+/NACLxNvUdgXLOX33j6X6wOQxW6+1I40YuwOjnBe8104IKc
oM9Nbo1nbPRVJu0ozb7r11GAJmKMkeD6OzJkTbyQ1StRTKlaaIFHrksUF3fwad4tTG4xphHKFO3V
ZK2JQtRRTBp27Mh2t6T6py4MK7cKLzT4NT9nzgqHnx7UhLW9MSNxlk371Ps0rRXqNv91d9Y+tyjU
z1Q4drs+Q/DC1kGmb98+IUm5bl9SC2sZ+Ss2txit/qTWyiYj3ChVpju3EWMisOyIxn5PImCUK++B
JAs+97mUN73nl+U9whCTbEOgsXn5FWHtZMCPvITqPIbox05XzW0CxvJJ18/qRAcARqUMW7Gxz6V6
tBT18erZ8XswzlcAmmFXV4Ok80oVgGyaYUo891sP/ZcDIGsAVmBqZKVDwHpufrppmcr/8WDaWJMM
RS1Of2MRxmhs0TWgXqQzF6jjcIyRp3+Bs+DMfYluZIR+SMl0BvHPDLT5zn9B+zxFHRmZWtE8Aicy
p0zANNjKwgxTIFVteftfDm/iP5NVKDCTyuRlKWbs95KwQNsa9ZhONA1IkwvqW9sqlsp6doglhZ04
4R5Kb6ld/ucDhYu81C2CFLLjgHbfMpQz2lHcH1buWUQf0BmcQsOD1SNNRWpWYy25P0wGQjFEeY7j
YwKnU8946DWLOMwZuPqwv6tfNB2K2h3QuvanQTR1QJ+lymN6jVMEOLdGYJprEBpvFeVkKB0IYDV2
S4FW6agPZ0WMb/kQzGt8/5gysWIUbQdV0Pk87o5S7dJBskEF3CgOxkujQKx3DoPNEWSScbGXOUYm
H1GJflGeVaRLKyx2CwP4uw96jV5DAO23oEqagwCqlh079kU3Bq1fGD0MRayDENnJ0tmrbH8dfIpW
yBxM7k8X0Q2vGRlC1fp4ze/cMp7cphUECWaPxyfTzAkn/Iat4DThqG6vpkRNTOFeM7ldR5OhUJDy
y7G6US5vEm5U4LFS8mVmQsp05k9qVm4EzQaZuEI5tIwdyYwUHysYJuxVV061plKPkGNM8bYG34N4
MJOkw0QDSK0TKaYKvpT9s3D+FSj+Qn5XEmko7v1hoVqPSZyD1kP37A+qC/qevupgY3sJdYA7qBb2
hJWn/SkkOQOBV503ekxN1UJIq8aiwSbQvK4Vn3pvkISHso+Y+NB38qwOFMCPWm0QhIX59YJWV5b1
LKvGhMn+u307ajwxNBFSduiE+UQVkMvxUevdten/hJY5at2PK0JFlgyklfdJmtTN11vr1PLIe7o3
O0rHKzOzpo5llEpnMq/cT7TQUIFsz8d2tYUdPMKK7uOQ6uLjTqoN6U/yeWQxR7+Esl95/gsTc7yO
ieEl8MEDq2j41fD/9fIFQ+ZJ0r1JgotyIjiyJ0k1OYLValt4zJrBJyxS2u+baiZP13fZgEdEx+mm
7te6Vjocj3cOgWNpJ0dD7DAUhg31Yy/WWe2xb08mt38gPfd9DA1cdzbIylQA7aAzJx0kPbVdxNdN
rKyoWJhFwNP4oshcCXuiXXV3jG7yO6Pn8BMrZ/wvy4jNtD4zp06X7iPOpuzop8RKPRxX6FBflmEY
uIDK5ggi+9Oe+JaR27smPBjpDvu5+ze+kkt4MfUlfiE1h/pXke0vaHfFTU25QOiv/hQF3/4P8a7l
MZMW9L7R7DTIcL0kqioJyLtiZW8mwZuLM8YUiw7JsE9BWCPPPN5eHJcPcPY14++YnObIfzK5+ELS
SqmEi0ms2ccT2BPsx0U7mOkBh8h6obwX2OHYP1A1ZVQGzT4g7ZfYdwpYN+WYDUpUd3MO2DfDSo5x
XD9zRHadyRkEr78nb1k44CDXseyKu2TrYUloZVr//lxf72mrw5iVc7cG0/h9YheHG+etpiWV0NQ4
CMJbRg42Ur/gfYwbqCbcFRd6dBQfIZLFGGrUrttaSSrsXJLSBIBSzslLZrnNnojQS+PAa11dPadi
OvzMwi+y4OMz7pdLN/CHRvQhPePQrKPRMymFqqUvgkPboOvuvJEvnuyiWTmQPg4jb+8Cl7YgPEku
b3/Ajeu+yVMZ6pOVYpnmtft9taxurBB8yMqLQLH7ypoTbjYgoRVbteMhy5nUkO4QeFlWe2hHOpF5
eh8lpMR9ECTNiUwan3TxNUZT1MYzoUpZl2nGGCNjD1BXNmAPd+sFLoB6Wi8bdWLN5laCK6PWQ13f
xdTzMVXbcWGRfsYxYHMFNtuTuex7xPacdVo+g4TNenFxH+2uQ7vPBxlzQ2WEb7tpJCoxTpcKKsT1
UTZ8cKUCXwqJGwaaNv/Twq5nFLFqxNqgjgJ1eNB9Gzq2FvpKxoK6Tgg/zvp7xB+RaT/ktm4DkER/
K33u6c+6GgSvXnZSKUGeP6wCZ9JT/1ZDN8vEmXCavtPo6Nj+GKpFAhvQqwhIMoqV8NlYB+dlWDTA
CUFm2bfI2ZJwWXqmzGVVfztGdZQBRkQhGdLF2MPTEPZO7jYB/qIYSHpJf6TpAs12kXqbh0HukVw8
w9Jcnzq2BUuWzgKD+8F6wqV1tSZ9UwmQM5xfoM55Ouhza8hKeJJHifPzos+0LLGy47OL4d5QHp9/
oe2uQrQh1HIKUEwPkhZqlhEhSdswm/nhNI8WK9M0jHzKJI/w+LHdO7kygvLGM7IbTVrZpUuI3xdB
VHV37MImH7TLLlnhr/7X64vz3jw0Wn8X2Wh+1TywPVH325sOW2hdBTF2qN5N3yV0KdAJ1Uiyo91l
R7AveNCGMfJsokKXYntr+e7hEz8kAGVwvF/Gb60HekifoWQyChhYH5LkXRqR/EnP13RYJeIOC8AM
FrDisb8HMTITnxmzzSdv5iE5TR8st6BfOkWpgnEsOj4YnmZZPAMG8/qm0nzqLAhftCGIoQY2aBDa
VM9Afyg/K1C4UNM09jzTu4oHUFn6S/E2QKywDxw8k32xIbFyd5kvw1IayiUb5PKJrMa5ZyiK+zDg
+HVsUr0biSyCjGI2a/J8GHgFlhkeTkMFgOxGADygEeKioQPJbbFQ8Pk6zVe6nsnWatg4xXBaqM28
k2G+GzsLUuogB9G3XBhFC2Fpsa8iny9GdJ7aLYNv4OFB97SqCxrYq0HV/Sk0XK7rjRjUXsH0AyiE
t1Yex5C7s9P7gWO6NEdY0pNZmAcUFAr+5JSIgYlsIyDOuncDv41qeR6x9or9nVsTy5787M/vm735
bALd2dWMKRDo7kYkm2j0JBNauncKUR075zyMNjqOlvJbgjWn4yEuI5SbW6nycyt3/BCxaDUgsJlk
jgmmv9pKzh5AqYlncTX8SYu4prL87Zh9rXbcT0cvJfxm6NlXvtpRG/5iAGetWPpH0iB3kmsunSNz
1qc9SvRd0rUrxtZ5X1i3LKqM74nTu715hn190dKgDX4WN5jeQmy0olFV7uZz4LbpuFzazQZ4K8MQ
9mxJXR127tVrGRvFceG7qpLePb2i0GRMFJTU8Igs6rjqglowHe/mdziZ6VGYx028oIQdfqBKtRvH
OvbKjFg+Xls53cmSjPPYHlbBNFYgZb/EH0rxenDAkFsXi9Ied4/F3PE8WntVfNVBkikYt3Aqr+0p
QDNL25bcMN2WvIe8D2Qij094fcNdpwleu+Cp/vXyd3JVC8D/mx6Fe5ku2fJshY+/eYSHfRyMu7Lp
cm5W48XDOI8zptSQSFOUIhWKKMGbdAtgE5d69bPnyttijscA20vupo4t+4l3+LoS2Q2O8d9XEM96
TZ0kHHtlqhRBlawOjhBAUQOUytNdnOPYc+iZ4vmsuMlu/AFEPqaexy/QfzU3SeBU83scCCTjHQF9
qfxcf4VNRge394xz7zjbXtg/UVByzRA3J8f44TcikFgFlvait9YWCVO77xozHfop/dJ8/JZxAyEt
GOndnw49PQeMfjKooGJAHLiW+jd447FBRXG6efpa1znAXFOhLGCF6K4cvuDRgbEU2Ks4svwuCRhK
YfgoWARY+HeJG1W2hYUlEAJXwm1QcNtTeg0+L8USBXQ+BpM+vGtqY2umaYzYIb4VAymTxonE3IYu
66xcU/7vM0Yw1QpLvcYlERzdm4iLsCD6Jl9DDUgG/+oVQrA72NsvPsDFaZmJywzCINa0RUVyrSu4
Hkm4LHCTDZV6GUHZmBmY3TYPXDBMWeRT9VF1T/HxXKceGPIPlc5F0U28g5C+CH/PUARUl+qYDl9L
2xzbyjKQIyChUjKnIB4gQ8few/OQlq8BBu4zLPpRaYkx8fAka90inZzfIUfU9E63D8zhjV2nNzl2
89xWVvKu0xUEpRPqqz1YG1N0Emwm7rLWh66d7MVZqDnDmCCupbHpf/xa1J0FWxbwC6IocK07EOis
SBlREObzARi979j3nh1XVoPQ5Lvvh2jjL5vu+EDKexU6fKidATXGJ59wP4QhKPUFuOk2yC6VLysa
S7lfxyIF3T1cLEd11DKxuX0auVuzFXs8XuOK3CXV3l4GPSaujOrHoWW1alHOmtdh7yB6F/A0e8P8
0Lit36n5nINuDioLgVI241KPHbztfYxV4tIoKquFPSVsTAmnOcrhCaZo1vv3ko281IEYtGj+PP/3
bA6RuDZXwEuVVHqULVeVnQuwNn2EpWYSdDXE/+fzyQTH994au4ihorms8pZCWlGUhZGA456/wXZu
HIIiySMXrNpK9MM40Y/lUD1eX8hq94+9bvOI5O6DOB6xzrJ/nFfTGV/3z9bHAQ771BYz4XAfPSUf
sh9/U76Z8dfaEkyRi8GL7kXaVEwo3u8IJ//WG47eS07qkSbWE3fv3niqghMz05uMot12ljJ6+fuQ
Dn1XjaeeG1t1qYvd8T1AdtIO6+I19IkuYCONru5PcsWIFZL+EXyWzB/0cop/QCSemiYinn7o22m1
KtlyNqAgxLGzRztXI38ZwNUzmi1nzxICLsE21F8JI2TLikCGLSHmdLDZquMCjAaQ0HKX2TjYdv5q
BMUMauZ+PUU5inRRLyuHaPDP7Qy7EbVWyJHgPrb73WnliPnEe5FSidKgQaS3zjsrRgWtbT+3gHYy
rXSUBIHaS+TIK91ECda+BT5eLZ7aieg7Hn+MN9K/f6E5PVpBd5UNZitw9ZFd035hpwrozU1z42Tv
OxpjnOmD2w5dvtyyf+YkBQ3/CvUkslCcpl6PRxkDMo978/8LDO9kqm84CLGw1Fbd4eXNx8xi/nD1
vF/qRIydWFXljObMk8M4sZrBLiTB9voGB1/vcXG9tdJbNluOjLRBtRuNTnx04KfNZNb3sNx8IUhm
toCVny57pxXjR3c191QlPT1UPar8d/457R7K53t2U6SM/lGOiFhhWk1svcAZjHdyYpeSqUomg5Hh
m0h4KnzEUsoxdLoc1IJuCx68Ld0hdbvAu9uLEISsyfHtW9fKZ0GMz0FzOQRfovGm6DtvwfcQqLG1
pcrO2R14nRiYORXnaDyNMDBdrqngaiLjUQlfuSrZca+fnaFr97AHkzKqAz1f5RBdTckG00WHsaV/
42+Gew2KcDxsZ9hBbDb1E2s9hOOkSTx+bXqAIDmyaGAOVXBSM+OPhrfo0vHzWCXWE0LSP3Of3RFN
LfL1VzTaWRryrxxRIN7BTEWyL7c52IFchDaPeisVbZw0TToC6gYYXlFHHBKT6fUgp8Kb4Dt6yi8w
LMVuvAQtxxDgAIUA07Ktd6IQPq04+potbkSazlpq4aceKoQ6V4dK5BNQRvKXsmxnazejDkRAdql1
nGk3dLHwoyzMcmaZQay2vTExcCZNtLGJojdLmEtd188NfFs8wmLtsvueajW8GsrkEE9iDQVdzi9L
R+xMVgi+UG3dMX3/2r3SsBbk4ZgmMw3qaktV8bp/Bz1MOdljLUqrt0uODEQVuGgfVVmsDtt7t51+
HXztLzclIHvdtRTwkS9jpvPVlbhfv3cbCQLa1n1Cr4kkTFdvjnjG0fUKkGRcHDTOMGAslGVLknUM
/A/r2Fq5336BYiGiYqWNFF/K+ZirLIHFTFFYtLWb3XI41ngDusno3RV9lNXfV9dIZwfMlbUxfsoE
KPC9FxPVwgMzlIDMxk1I19dJlJCoYuBil2XVlhijqt7/a2kAajfAu5XwyaQQU9UzHC1Oj37JYNUn
Q+32TZ8OKnCoznb1dx339oqVO/9qmV286eIDgeADK04/+S+pbPNYSzz0TQ/Vx0UrQj3G9/YRIVLb
zT7iwlPcCyGLgIfOUeVoRceIE+t9Ps7kqgfPR2HwEO8ymRxKXitwk0yhS36f+H9i3stTbWi3c6XP
WUxZxoCS9iemuMlUVAbnAef3wT2JZMBdr5UxssBrGSXlsfxdL8lqIBtMw22tkat1Rzi2BKSmTw8N
QivAif1BMYE2T2OhC4Z2AWnmTKhlyRjvF/O9xmOvsNk2vO+H1Uu4p5cxWbeQKyGly+LUJwcUBnAk
PEm+xShY3p5Vsbw8QGcrqyqbWk7PduAbQZTFjG24oKsH09BYzQtTrsICNCOg1Myy46rrOK+KJVk6
tZqo4OXDTqmGZDCwz+OiNs3QEE9hktm6JY3scN70R9RzMf2Iq3NUa1JMT5+JWjHLsRwT9C5D31rU
s7kIqA3RCucbwi3Wj5AoqOSxDmsxDPF/E1dS6Kc0mz9YqogowSE1jQCNogxx0uz6Nu2EOGTSlVdx
GjWZ8QH8+mjoIiugqXmQXHFWjMN/tvngEKdz9wObpTj6aTGmZ5e9wSHTrVRyNSdPMRMOPHCKPUaf
m3lrkdBw5X0F8rcY+sERf+bHX/be4sNcx4hKLmGv5VpvWSHWVVB5WK2UmUR3AbrLSsLEexA9dLRo
bVVri7TqYjpXgb4dC0ITGi7S2Xe0SfYw69nyvDqP+VyjARarVmBAO2933jfxLUaz1bqxgJpvS7Cy
EIWBZBrLVDABDTpptvoC1puyfkasvrT/Qy2jZAhCthXchUQ/8wFaBaZ0dmCwiys5d7A9x62Q4g9u
Ak87hjOWj1Ak2K34SWwE2Ahvs2FRb3Dp5T3is8t8Ym5MOQId5sAIpMndSAK09O24eh6cF4JYvszy
4PjBn0LHSH+tKBP9vx9H+P+SkcVS7S4NpNn3JY7JJS4HWYpi/M/dd2N0HKEai5/1EMDBLgOb6rMT
JJIb0vKlpp08bvOz9cLhLY4bdfDKRtVgeasId6pPLoceeduC2ubtVbJhTN8jizowmX5oSTJU6m2o
GZxTYQys1H8S01W00thM4YWa9W/ca0ZXf0myEG1hsP1mt5rnqGesFnXxgVYLW/QV4O4Lpk7uR0Zu
WgG4FCdO+uxiVdnH3fk3idQIfKiLMeJgENnBQz3vXYYIC0a+LrRSkSjdWCHrA5wKdqIf1pkoGg/B
Y/lNzH3Xn+yiyiXCPEgrP7z/6DCZQdXre/x8gCC17WdkSzgUVmzBurWza/EY+hwE/3P8q0h7kt9p
cENKPDRCMN5IHCtvE2CgL6rhXcXBFju4iN+NBJn2G1KIdxmxeEcFeRIEO9li9emmkspkx8DOkoTS
BiqUhdtCX9TNnxJWFdrW40UxbeqpIFdDJaxh58aVIe9kL0foPjf8vHlVR3NUHN6J0fNBgJW4TFFi
+rzf/e78Q7XZ6+6DHcRsQHDQdFRWy68NM1vHoi1hNpkEC+TqFVL4Os0c76K9LOZo+roylNmPBbGB
tVU+ice0UID8cNT4SOrM9wWf6LhkR/li0uD9V9uFe04oNwMnP9Dwqu5ntOK9moez/i2K3SfHl8Aa
YDkguI1zxqeiQS78bF5eAnF6p1HrolJpDvet4XTetL4rTZIvIvfvNikxVpFtIJImtyXiOTj5VMY3
QKdrcWtOsO5L4oR/tEOVAeWcwIcYPq4zdiETkIwq4QfOhsjH2DpVnxHn9c9UL1ivpfd1elkSN+cD
9ceRK7+Xq+brqagW8rU4fROv7x2epAy0Ae5+jXDjdfdIU8Et0QksHjTf92WnEu5VdDTUPMKREF+z
oRqSCvrNi3LxdkmQSBpbkyh1Ck0XClQEB1IJ+V++Qsmvsy+8hbDkxMcxxaNt2quFdHhvZzIL9WJR
fNNtijBY2UL/I3P/vdXs8H/8HN02G9kp9d7V4EHD+v8cO0EMFTn9geCasXMfDgXWyubjokYaVNm2
2z4rZqgT6MR5Zp0guBf+b/RaF+tOVcglLKSnw8ZW0OBDu4Ifrh6Li0FlUvPsBtXoYJtoNHVGu8yw
iqU9auO1eiSWdqn7wWZiTsDXGDErM2rGhKGDRJv564RGY+2OphTHb6aXqvuPXM1QO7xkqQ0uoBH0
AcH7DuXl5TgPoF+ugPIEE2fE8cxyQKYX/pQYLga4caYBtVHc09Qpeq5d8kn7mGxn7m4BHwVPclFB
mI5+hz/jbwUp2qoNASQRuaNJWr+IMxRRgNwYgKD8GamGv6bJmdpZhG1sb2BIjTYR91N9K5taSbsF
VuESg1X31WQRQqZD02+Lv2F/qJAeugn2CTAaJrU9P+D/9mFC4ll2SImzRqePDH+NQRtrvdDZC2ae
nUyNPBWTfXsZwqg4wJXwhwjPRsCMOkXH7LZVPt/mWM1DvqgY2Pf8BZ1oYW+Mh1WiS/g88hWQ/ACH
VWmNnilr3VU/RDZxeiflYROOVByMdR42J/7kQ/+JTQvGyh+eD5blWeLKbWIz7hrTYTvpsXeY0P9z
C88trJiYW1ryzkjVDNqZsBz3QNdw3nreg9opW+ZKQS8D/oDAdWuuMp8ajNjnPOKeNglWwuw6w8Wy
LH/9ROso/rPj8KcFwsv3L5xuA+UdOklShbToHy2L0uEoKORKvbwZRReiaCVWnaMqE3Lm/sUXmQ7W
YOazz8NGGfKzROvnDpcQthE2F54CkJtaaB7oB78sI3HIYjne5VAgupaO12USseWsmFKPeIOYAykt
p0HKO6mnwXDnoNKHs+u+0F1mWmKJBrhYfg7h+rM/WbgrTLoVZiktCc1Z/+JL/eovE1f1Dphaecmx
nakXhNLsozGaDiErky93VfEEYFRMYXGChcq8w6fFSmejXAGXLccv2Kf9uskmXyKsUlh0xJLY2oEJ
maJdkt8eRojfUirP7M18UReCnhWyEh5GQFoNrBlZ3ukfDeryZ/7g9gBgweSvW67OZkWuRPT1pCDz
+w7NQHy0s3uJfGthUAPszj5PU/0L0uPjgRmgmJTM445JTJQeEg4quKh217hLI9N2pLO4fldThPgv
g2wi4UCf5R8HZwDG1MP7OONC+9fg8TwP1hZwbx8B3ld1y09mU2cB3Tq+UHjEurcNaucm+celQc5U
eZB621LYSWXAKBX7mJzx8FJEm0O4sOTmOzK/q/gl7VhXmH4l8lOKqXBmsaa3qzERkNWmc4Ie+idA
AdzAffAyNYXXqR360vIzfVGdGDXCZcG7DrPI6Nv6DlVivVtOk011KbxK5f0U7+p5HiJBLASEB/zS
TyglbVufV5JyDRND7B8lzMvhpqHh9vzrKi1NSFzjJp4rAAUGoNoscydN/XR9siGtCFSkN8lHul1s
kgGv18lizstb2M+mHhBGL9/eU/+pJbwkmMs40NgGxvLrl0V4898n4EuUtaYM7cIz7+aMce5ZVfo4
HIsl/U0Zbd0v0pS9LhEO9CYgtRDHzXsfmLZQojY4jsluGJ0e0e+rrIxH0VOw8M0zb9oW+7QL8X4J
/i+/8G33cHCkrAdttDma2l9UMQDFGDq5/AOp/e3SRoTLg8rlb4kT12g8O61hCZPx4E8f3a/hZh60
YBy1eT2RiWxQi8o/WtOispvC96XG4sLOThjuUTWbEZGAXersFg4WomC3vlo5t15fku7/CHSYNhSp
iaUzmSP9vwwBbnRhEmfQqhlhBCXEArYeyAMILVZigquA2mS6nhcc/XfW6s7VEyz9wyQv6xla1fgT
5uu3dIfEhw8HFjgiwKmgKsVFc4rvQqnzpUt3WAv8yM3CtAC/ZSHAvPwvxNeN0JpyhSZQLKU3atkF
vyFSDplZb05jyTZmD25JqgdC8hw6al/0zEI8WXt0K1VPxh0T8DXfqyAI/PRVKC/hTBz0LLuhh29m
SDunbY+cju9sC4CVVWrgLvaZdHz80N838Y4zsN1qX8v92Vdm9sPy32Qx+FwwTqvee9VDPsW/iHQh
2M867GLW527FuiGGqhbVy67vEQk8Cqemtnp5yuUxN8C1YxH1Q1ASP5BRP4XDBADOhhIYbp2oVt16
lzT4E8voer6jOnVrhupnf4OSm11s+5Xa59t3J5rTxgTAbPL1pYU8TKmpf+Gp6/EFHkz843bpIiZV
I78Ma5OT7kRYvV+ZVSNHBm6qT3tr8GwcXMuqgCkGftZIfScN+wGI/8ZtpdUAvo7vhDyqvaCXRh68
nL38UldB77qSTJ87NDGPpx8AydfpKt5CdCjzK7hBkCd7kddVgkJI/EQkAs9kj9emGoV4DejvEp5a
4cIojV6A8jITJt694eXnOqTAK9N9bgPihs+DD1PLK3PR/1I6z4E47EvyY9hOUhutjoN+7ieeoxIa
x98gYS9k2dncV7lK7Q+poDnqa6mrmwCe17Pm919uZm55Uv8XclC4mvKKE9/CTcYRbbtzVRarxPvG
mIpyYpulR1eeUbpAne9YeyBp27pKtdggd36pzYnF+jDkCmqnaRPTDgmLTRTacdlqIj0kDp3a7c3C
gZ6H90AVV8ryr+IRWgyQKBAD6ySKj3fZiOKItl5vJ879KAJPCn82Vp9YQw0oY+SiZU4ERJNsX8li
G7PoS6HqMpwSTRel8BGxezRI+MvjG1IoBBQl9mCIojhdgQ4C02ajEr9pGgKIuXag9nVCE4vHJ1Cb
yQhejOuXNkVVCcE7kK5gdpXnmPz+G6rI3kDMMUjcfydmRn4sZa68/itIi5UhtjZvbwP4VSNlFNYE
szqV7UFfkFcOdb0t1nii5174IKSy6vr/3rfy7+EJ7/Qra+3rG/3DmISc7IQs2QfXmwLwxSKpFUUl
/RKwqfX1gaFU2AOhh7p/NMU1j/xvvXHewRizNJ0dghUQRWUqYABVQXJ++xzNFe8CpyJvLDl1x7T+
GTEeFEyklo6bHKkifQNyhrYoBsFUk07Ub9ZJoi0iIv/3Fr+tOyrg4LOwlgmSzfFV/H/EU54kS79F
edC7rH51QVpqa6p8pJVkj08gfx4J5EM+bVI+H3ImxU+2NpYP6jsr0bqfqv8jdG/V9Qwykn/2o7Rv
mYWqgW9UMXhATnpIxOdYqQuU4VyX929gbImivzfTiBH/xUVtUNrtsls/F1QzluStuCEe3q+bc3m0
SnFNQSt9C6pGm9WX2IpNrHpDGUIX8ixaU+UJLmukWPZUU59cs1gtu8I0yQloIjAlPD2DSnEEsd9H
tOeEKewacVh7xX/YeNG+bY9PrUqDMwHWzNJlr08oJe7H4w+z4Nr/VimX4vy8415sli+uIZ+DYWWF
zIRnsF/WfTuzuACswQ/PMB3YgU5tvnUB5sJrLKrX7pOuB2NjQj13Lv+SXFkksSDbvelm4pipn/ZZ
iTHaP2OZembgfuxZJPX+fVQCyKP7PeCyNesi0V3BdXNVeA5wAYbe2wb/mpNl/5pXwZ4Fo4+VRTQB
PNsJC+gq78wCeo/TWWYg2ayLknomSryHkm3BpYd82U06oJww1+gmFp8Vbk+MITkUn0Bu/ymUSh9r
jcsT3plzdd/t7k8xwJzdZq3xDikM+XOLdh5rer/8Z/tEtkh7TftOemBLGYcmwyEQ4VklMJ6DTm2f
mVNK1JaGXwjTSKM8XFNG9acFMk6pG0/tSAN3sYHNJFMeSpQpU0D/He1MkPRBMSUgJGrwSprX368Y
a4/iqKJuSvxtEplX7fdc7md4Gru8QGqLlC9NMI1ZA3nUd1moAqIjGHQ8kh95pYGPzrHmkFa6lgXO
pTnx2jsowYvxLosj/0GDac8e4agk1iwsmwb77BvWgJl/jDlJFcfSgdH1b0rtDmdUOLjXCqr6e4ap
2wjg8vIx2TKcAT+AFGfcD35VP93HYQr8A4RsOcWtoYh8vDWTFcpYKNN52OI7lYk9cCbdwYL1z9XM
OZiJ7KNX0wkEgKmCgpHIieu5b8KSolm65BtZbR7P0ty8gFGoDB7VOSp7WkZM5j817FAvggGNUOQ/
prlsA+o5oWCYLVYmMOiZdMRM1DFo3imA7j3K5mI/S4qrXL21mHbRQymhIyHbwmJXo8c6OXsz4/xU
poHVWuckUax7WbhaSnzzoOHtoUZ/Z+rFJBbCS6IxThUeHYoLkOsn/8VqhNsFTiZo3RROKedgRjE4
0DgBmLGldqpQZE/3nXEPryR5OBYDkRcBlFSrdG2wPFJaV2tAzy3cwqzlGQV0INZr2/jYaZMdOyDN
px3Gd9n+O6OMl1zBNeQeIoAHrWGwrKE0VgT3v/P8LK4dCdO0XbuSXCqFTFAVeUFObSGPjLyAOaZ3
u6O45bcVkodlQVTGeBCf66evcePH7JmU3tDb6rL2+icrxxyAhQFURD7CZM+/6U3aGdLWbZ4X+rlH
Ig032SfyrBYNSbggoq0/MbU90pKk4qjsGpE014TNeHyBob/MdyYYdUlKWbsHfmGLIte82ByOwNBY
d6+C2BmMH/7aHb47lQuvCMNqAUW+/jNiJz0bZeiGXShFj5Fo5YwB3TJksSvQRT5AVSfx+Aj/rPbq
Sk1OgADhXCMzltkRkbsBOLnuorlsQWarOY4cnwpWURSk0T3RrMf5KMHTT5PDT/guzmUIlT3DwZhP
HKVqdnYjGwbPB6nv/3VVMtqosQoETr/Wmj39pZJBmhsOdo3/rkhfbLfikUi2oNrzrkTiO2147nkm
xoHcclJEAqlY6mBOm/vnl9+9aU1p6gR2pFJC2N3QgKl2lBSO/EEr3bIYXRuaFtQWtXf+48sWX7xt
Gmie6n6LXkXmiu9DgaZujomoVPRMeJv/i2kdLVlTBR1AbQN8jlVivWSvThP0tZV/QLbBlTrk494N
J3hN2ejfqJHvRjR2Ao3++DGm6rBu8NxMJT0qQxy8IpCzs58oID3fNGL2gK0EOeCdBGD+bSndSlVk
PXuPe+g0oYpEE7LP5tIUfh+2Da6oExUsccxZqPK6yYNGGYKryhfKCDKK9uydvbEYmrhDYgIwdg3k
ViZEjri4bIAt5x1dHQCuHjVXYEkXJA9V0vwJOCigtQCLGDSiEGlUQuTUMofnSP37Tx27ueH0kxCR
iAew0zz4Cn3Je58YzFe65RfFc7wcAJ7JsSkPVykEabYDeoPmpQrKKSNoGkRoDJmCcTEFmPJJsDCI
TnSE9jn+lLA5R/+aujhWrRynxTukjc5OKYzTaRPwQQ7Z/sVMWMhLOBp6CVkSZjUxaGJuavN63Wtu
nOUPBiGjEDvjFa0iCOZ23J6vvaFLLS+VTOrMvsSQiFYV0q6OauOkYbTyeyIfK7AzgTpcAYSGdsz2
VxpeM/BNXpACLn2RlsTFHXZtCdmSBJLcFETr3iRfPmw9YHX9+Sob6TMDFY6xk3CfOOckgyNl7ajt
Ezqot0XXYqpGuZBKgBYKAY4hE4mOJjw4nZEYI30CI9/rCqOKkJ15X9ZQtaPycnQyt1D+vBGna4c3
mzmWhG7p0bdBa2KbjBSZMq6LRF8siljjdmPpaxLx2gwPhgv7capRca2tjzF1C7MPDGYUZIxnlwL/
TMSm0Xu8uKjLbHnmM8twh16af+ew8L+B68GFoRDcr/5no+PDnpPsPPzr+JZ6umH0fAnzGQGCX8gd
qppLYBw6CNqFvzgDQUDUMOW/F6Xj9tj9aBk2Hi+TQrWeS4NhK2BO15x0SgncKB8iHHdUGbSZzcbq
1KQ8zxp9OcJ+v0KPnQol0gCL2Nt4n6yYaTdMcY/kJyg08GqXKED/4g3QZoCea4azYnbzhOiT3uK4
rq5hz0lac+/in3PkIfmTWQj/laRKmOcNEJIUsuMukeOxtOEvIj/SkR7UMKL/2ui57VPG5z5I3OsT
3tYRM4BhQg5xyJkk+jwcgewQq27iSaU0Y7E4x+WaTADrmhX2MDsOxOn3mknKrD5Bh9rqM+Zwo1h8
A0sOIc3b3trSvcBJaVm9Wd85X9I7Eh9avC1538ZSuGiPrC3wHFmGGeKhGEVNn+TaGPY2/3gB7Vzi
tQvWMO+EIdZR+/8Wq9fN7K80576092VtrDldxcPhJm8I0XjaAYsgb+xBSwJ+xmQ7dEe0mW72OikY
7ZG3AQ50lySKURKK9mvxPqUZYZg2eJ5eSB7/OpL6T91bz7QyuGJtpeoR2/grwbayti1xJ6rCgrue
gFScavy40aF2IYMrb0aeSM22HNAHimh1h8XAMKsAGLJ0+DBtZ790yb2n2xKPlWSaddV1u4xGIJJ7
9a8z+MOJMmi9RQzpXhJn4pwsn6NSn+5soMoyDxLJRxsnl9ptqXsCqT0yY5jdS5Lwk8w5u/8qpg7i
BWlneULX7O1Do7KhkCfXZNAQjv6xkZQk1w2SVTWwsUIil2W8K1C3EE5P/eOsQEoFlz3Cx6JSw7nF
lY+Cd1knR5jvR7byKs2X2qZzQrgD9IIfIMrAqhVFsin6AmQvG2WJ/oeCO9n+41LSSAOM3PY4eNX1
4J5dKF96ZDruOf+4IP3jTmgjFZSyg6NOYL/Q7k1ZBtBgJKrYKJOD+3fxMcaCElQzn+UHLvdPZia9
AhgmT+RRctp7aevoCktfHMg8Q62NhRlgOE6J5d7cVC6C5QcECNsnd8MED0RoUD40pxDgYOdnRgjG
Ksqc0MWTNUwQ5tQzVAVvjvh+dWVJwggcnzJ97eRj6D3QoAEufldqm8wKOwEpcSfdtvijvQMpredG
zmDOokYmL2rWM3PPOESE4Q3TKJaZwRb02Ee+mDFAvPkG3PuMHu4j4gTBe0nkDoKrgJXLTVrkzORl
cVwI3yZTw5+M6mia0ZuCBZQ14JMdx6COzB+jKEbAFKNUH9N4i4+Blfnr9CLqeWLAzkRZnnSmJ9s1
hO18QWJbr3UIEzcA/JYHfi3Rc7FDZUu9nk4BPleC+4L7ozaFPeCE+SV7e95oRPFU6yyEt2He/IbO
kAjfQjSC9BfVPoVvzJgHj1+vzTkyZORFSbPamxu4qkHz144Eis355mNKuF+77SnBK3k7gv78PHlJ
7aQYp5D924EMMshAICog5QYGZ5HGMI5vP4moScB5cTueLOwX3S+KojYCY/hFpuaHDX3J/rz3Rpvj
JQYz+Uqb4kq/6tdSQjnYDfsUZip4uf4Lvf/LZVyK6XpGycHKkD7tNJsYIym/ehEttRcsqcskJ4/W
lx53FiBAWhsTf7tNqXFzX38cxQ8aWA3vugMr5piuh6WmDd+Mxdg38YW/lwSJX52lNDxn9RsUneez
50SolmBkry8CsMByL4YvLil13z562/SlQlJq3ttf8cOhE/0Iv4zsdvxbsUSrWE/rbZek+4/WyxYf
Lr47d2hBqeoRcE/mnQCZA3uohJBW7HhBvxvJV6BSearFjeUQ6uGbE1sbsj3cRsbtntE0dau2S3ac
w3xsWdZnMx4tHsjFNs2IVpib6N8Tx44DVi84tMPTez/PyHnyMkiHuYFm+ejI6nIDrM2Npj4PC0mg
qOnVQvprTVibOnkZnvIX6i6ogqBGqdLqDtIsX6n4dLQ2AYKX78B0vBvGWreWe5QZJA82GGEQRHBZ
GEs03nhogdKVDBfzdJeo2h/ZVKoarg5HpLeLDNfYglOCS1hx6KrXa2rKsADXGoWvkbUO6RmjGohO
v47rdd7bLf6bkFkCpIceI9usoCtTYFsPvvQ223y4ht2yF3i2IxYskKsU4+fCtCJ/iKcKLvLUuUy/
LzmZogES7Ow+QFFLgo9y3Rn5b4ICLYvqvPfLWYFtpBHWlQdBF2v0MnSW3Xiga4g01nJKcpBauvmx
JtEfr+fZ0EEK+bzpWTmMYkxyxpidD0Y3/pPg3JOJvZDR39P9dKOhCFhKbZZ0yFatDh81NpABZX1C
ojZysLCYqXawai4JjdOZSQTS7b3z7c0PuWxUlE+sEib4IvuREh2kUhj0n/AWqrDvFqAuEiuNubNj
5TNx73OT4d/dpDYFHpRtyyzSRex589eqZ5zfLfgBNccD0Drdvqo3WE5b8PH2wk+MEuhIXObOQYCH
58hsyDDZM5JxJO1L6R17385xmRsgCEveY27YVeYZlRXbhxYfZ7WSzG1AgVBZByWqydHvUgOzCA9T
tm/KHflEfoeRKsAcV5C4YG6K1Loiv9+skCDIxYGSbTskaUalxiq04PF9Ml+ZnbL/mKnbJJ4kYekQ
LlFRXAmhouP9hp6n53PxP/8PBmtYdiQZqrwf81aRSFu40QSvN5xdchUlw3VbtGqJfyQk1Rik6qm+
lUV2MgXMOmgMzgm0YnPkOB1GyqJduUlzINRfJvkCyTTbwg3AXz9HTD4l9q/z4rOynCM0n0oLILPj
YHN1/7q4rXhZYjUiXXOYyqZUZScNnL2ClB6caL9PQ1Iz47VZZx3nDEOy/fodYmb1NsryaSr6xX4S
gCKWAE3nCrFIOlkyBotixNvODN5n+epUjFe1KuT6k1lQVAk9p4hF1c9vXgaCE8aWAQQ9oAPYoEhk
Zc050rnlKXNn6rX5dhdMNsZ36xPcIIT3cD5HlcL1iMNfIu1BNpM/ka9wnVJ34tagYuLI+h5J/aBp
XOOnVwkThr6fYyuw180j17oNt7tc76X1rfMz3pTPXGONgEHcd4yaWC943pUl2n7s6diexfO1gNKL
glOK6zbGuftiOoNzKrq+6vVkwBev4r+3Fhmg3IELuSlcYlpsfKAz6vrlBuj//wigXvfvmNgrBV3G
gsnIOKCOiYcxHSiRfwU1bHqPPe74nKy+0ctYDM66VyrTW+uWNQpx3GUqIWDR9geto3Zxea6u5W2A
IDOjrCa+QOuCkMawjeiM4OI1JyFh2OJ6vaf6C+2xn6PyePdBctihRVsNjxmHs0ZIWLcyKtTrPhLH
p28YMBZPGj1y2PZZ+DM9rfSKwwu29ifhV8rCV0Bdlk5OuqwscGcINEIpu9qu/EVFIhThzR8WFh+w
gcOHnHL21p1qtsNtpiZyeSaLTKx1SuHxHDL4xk4v3hopOafz62FpEN3rEU8H7VRo9gQbqsxBT0ov
gud6zNkuXD5XQ/PSuPmDMn+kCybo9x48CvacE8Pet4sBkOqShWqUJfYOGyVMgusaY76m1k50I4Lk
hHDKB5JgyzMJKuUxjhH5Cyiy7K6MF+1ArDvxS1L2Ne99miPndQbT8TDJvVX17jkCIsVOHLPLPgzs
jzF1FgMWFL2rMGVMewBbe7Fo/UQS7uCfYdOZU73N4KF23uKvdMyDCW2PQAjMcJDZ3gS3KeZBL/81
Sxvge6+yXUYeGikrm89Ve+hZhf5sQX2KHfL5E6azOlTE2cSCNlQwQ10+ZSAviHd63pztlbxr5ZAM
Hz5CQ2NDyym/JsxQn292Gb6i7Q5TKSSxL+jGjFdm9LDptS9zwAa+EYADQWsGoUhxX8qv4nER77Iz
BXVJmuFxrSEHefFhBk9/5cXyPIS9GaqXVTCA8EMbFLDzbY5iKmtIwkEvqPRXsL7cPCzu5r5UneeY
TckHZAmC5OqMnFHQNrkjwOTAlgJGLb78d6q94fMAbKHRokqJNLd+VTgAgPF2wW87Zn6NagoApV5D
MUa3XT67OGQ4Qj/0u5jnL+9tiulvys2ynTAfDDYEeD4FV8wdCEjISQpxUN9n2WcCTI3CJ/YGYbTZ
BTeuRUwf4HxJqk1LnA+T+mOoCV/lwOKCub5/kWYdHHxLYQINQBik1RZsKClXFrOJ7bCsTriBK7x4
SrNGpjxWNXVsxk6pnqxvYW6KMlcELmEtKjDFpdiyts/Wubu/9uU2f0kB3CjFpdmpjAUY7LMTxDeK
gTqNNmmguPJP1PZDLPGAkvnpq8GdGIIYAKko4ZzS9iwgfCFo24KQPNelmgWAKLpJ3MwgU9GbMiZf
IN30CvP0+vZP/m2t2mhapzhsmofBzia8BAH4LhX3AobjX+z+mSX1Rsq5DxG+HDs/4CHuZzLL92JM
iCuLHMjGNKqLZQKquBTzuuA2Vh102mN8DiQjb/13jAKMZVbbP85RvQXCky+j7nMItuBuWt680a3q
WTkSd6S0GuYkfdnMtKVznBpVwvVPmN2uYcfputhn6iSDaNdqxTwAX25mWgUv6J0D0KzhREF40U3M
67tBs12rFidY02LFOepCO3G/lcNOPZBMgMMrG9yYtlaRzKEsw5G5o+Nx8AQRVeDXV0dLOVwhNOKL
2347x1nV9O1o5VFZiGLEUNBQZetrkgCbI2sSFVnRSY9hLxZNoO/XMu9gUSU33E8i9yRXNJu2O3tJ
45FHyLoFL06qvvaNvvvZDkYLJYpE6IwT9LxpQQCUKjvJNKvGTRbJB4TIA8672MhLMa3F9KP+FD23
5rMjwiwD5AiIpvhAuHDydU5hgaKMz49ABsO6cUxxNyzCT6Unz9Ne87wTyu5LGU4qmwW8ghOYTCXa
T4e3RT7FVnD3pacoF4UCDrVUqKkO8eBGBk0ocGd7jS8jKzth2LFhnAOxQAedLRHuL0vw9wtOddK/
pPaHjylnBSzza/3bgHsSo0J0K2UlyDKZjqeV27Q8pwMyc9HyCiUEFA6xKXqnq5UPphCtwjZosafe
ddZwyN5lGYojGWVWMKjLGNHw/cIHJJwskAl2m09ggxl0ze+kftByQI/MQk8q0bAc88H71+xLwfUB
ZuBWThCd+aWYtwosvT7OtveSTN2Ao0x3SYa+VYGVOuU1iQMxxisCGL2eDQ9Ywg9/SQCFNZtB1Dfn
nCzIK9zGrtN9gE/2ZKU038WMhvpjW+QOiFnZ7eENwcNRvfLRrpLp52jvgecXS9lEdzYvl+tzgHBv
l7ieDnLZZC1XGO3lwgzVmHoSuQgmImHxpnKdvyn98YdImgjaL1BabXu4qZz5foLl3ye8585hIbMs
Kv/bL2UNHBnTiITloi6r98V7FTFfNGJnj9q+zK2SpGmTmDGH46f73eVt95eDXgDG18qAFaCtw2oY
DcBmPAC9MzYfAuzh9s/rdwNZuFheRnh8RrGLxvb0ZbcKg5rzEm/ZC4th74hsx7nncGFRlxKbaAPG
v2wRtNrrvZawPn7rXUXROLsFDMxXhpa3uMzEtcVxU8IpxpJEHw+HBKaGJ+cZncVjVhY1xjkFOSig
yAaPzRUpzRaxSQmQ88RlNi8rq5bHpfYj62SThNHEH3gHWzf1O2n4Zcu1w+a5dpVYy6HJoNaVDrRD
JuQMktukpDnlRTke+DQgY0fTXh3lUMxHv8OQRIVed4FOz23g3A0sCiSFJCR96GugvV0eWRdVd+vQ
uHDpoeqYPKiwJPSXuXOuaRGPCPFdFizncUUDbWb/Vy9GPquhwVEYoCeRGljKjBIj3+T2vdv15352
48cA2Cb5Vtvy28+R84j9UEheqNPW1Mp7ewmONqdjBBflOn5B3y9SiC+c2ubIMGrQ7XeGYVnfYv+s
T9N19NFJI40ZIOqoozUnDsJU7HaeQ28tzlkGvGrezxnV5+1yvAJmIf1KVGgRpRfdGswMsPQUZQPX
7slPcCxAsHB5T2329NabDdGJ5CIMcniqp4mN6b8OMBHmFMoISVVSSGGbKOpMzICkVGM4x3l5jmaG
eNJ/djI4O2Caqk7aQ1tmcfNpDg/16lEvjZTgUF6khg+oWHaAEnuDbt+rtAZWXoOx1A5QNZBWP3bW
JRnlFOBU6U69r0K/5+S1ng/6GwJ0/iR89zy1uiM+dRr59FAfeqLvEILGOF/gl52NtVR8yaaeGel7
KJACVKAWs8q2PhAvYQIVYoQPJdYeg7hF0tm/6BLA0g0NvqVz7Tp+BPs8nMf7SkjWHvwsB/4q+0Io
S2IuISLH6iVRpY/FkLxEjkxAppMM4/Mq2fBzyoPs1lnepFSsq4oEK9NRF33T6aQptYfdsoXEi1fZ
sqkeQlfFJdohRpwUrr81iFMPbxUYiUX51t1F0DmOJCc2KqrAfW1Cz3rY6n+t/fdCikwrpfg4NAbQ
bUIAU1V8uRU/fbHJ1HCph65Lz9HVGu9RWuJ+/BM/8AWhZkRPSYsPZWW84NHoyrwxS/8QyNOMRih7
2/hESgR0oRJYWg6ibLt5GsW6uxOyNg2NRcKdAhRX9Z7Clqvc0YI/1IcHmZ9BFDQ0m4AfXkQCFJWz
YCNIkQ3wQBh88gTobGL3t/alf9ArHrVokTbEN7hMqTtxKV3/gxMaj6VhPATikSOaGsUurOJ2cCaN
CIzIk1STVq91xDdE17TCoGgPIl/1UDCMGnrvYKVuOz7qe0vyc5o5m2ezJiypQRgW4E1Pk+bAoDNX
elP7LDtshD9ar8MQIsKMtbm9isD0Rxi11XwpxLBuAoSXxiv+NoI0j+5bLQY2N2p9vtg2jWrVNpx8
ZfWVP7zubxkEe7LtJqPs3XgxNbQ4LsgYvCO8SQLf9baYBhoe6eyJ6xbiHc5RIj+GJStE2rEc9/yN
rvgltKIU18b3Q4SB4Yw7DiB4Yb4t2mvwbraXRAl8Cu7ayGiHdb2Htvu4Idrr1BChmyhVrb2TEwc8
jTxkMb/M/QdmmkP5vv2orVHciOz9q7Q2rdVH30U1WvafYby6tQc8KiWeNYwftXgij4MgF1nIvWHx
K77QoCaoBkQtHQALmzKR029WeL3DzjOPuMX2089PtWUQNcYK7JgstjdWg4PL/V4D3ZxjavV4cbNb
yIwj6Hyc/pwvgIsOlYzUCR96Um7GHGFo45FtzAyJBDrLSK6EpsyFqGpc3aAf0BAsKkU2VaOWwR+L
gZOOWIOyTywKWrbRkSfTDApkrFAJpypcjNvrJNsn06imtv6ly8W7YnF30IWZ1lxtuhjQd0zan7lr
QQk6q5WXKDgDPZjvOUzCGMUMTlOUtAmStRQ8V69IfQ1sTwexWSGx2Wldrk0IUOFpOZsG2vaHaTlS
p8dE4MogpqD4Z37amtNEGV1pqdU60qBi7hj5JUjbe8BN0cRP4sN3pOcd52VT3dfk0gDXk1ssJJ1w
t1eS5N25CywUKsy8F9JAhSCTq5kn9ckyNouGc6DnTmuo+IL7wR8WtBpc5JMX4Ui+5oR18VZ9m3NY
FAVMfkjIuAy5eXLz+RjtCjvl8KyELmqpUwvEbwUILTSFklIhtl+wPnlhWKUJcSf/bnV04qUBDCdR
b98qkvFO3fiksR/sKbtT3ZuUOrr7iyuzhTCADDPtfliiJRWhDNdS+s4VMFzq1zHbcApXYNUV9JZP
HEnkX04L7d7rfbh6Pz6KxNz0NehSDsXYkviEoDoM9K1ivmBtF9DPkNOZZTMgnmA7zpJnacoxlDgw
BZsHecidWWHsJKdBAru1BY2J+v3iqiCogSOWURkXXuNL5t3fZf1Sq9Uw+ric/NxxgtUoioUjPV7F
MZTAnUD2oMK6PzPTwuEmLuZ1zevI9AjWEUFtwltpBR5XLnDuCnkuK1kGN1YRSObJVikZ/QbWDS3m
tdGmLv5PFEn4ddnNoE3cMKX2py8m5CuPzE24pGbuVsP7/vI+wJYrAMskdCcrWlq93a/2WwDlO9vY
CbXRUyKDZ/SHxYBTbZ5kC5rqBQa7THUmmzkVBGhyfM/fNnYdmWWyF7k9UN2f4FVb5xIxKjUJR+Hm
q6+q/5gCjklf2bzl38HP15LdBFyG5HYezOBXEaULVYBo7M/u219atNBGLAjGa+RZ/31F3LKq3vid
k9c3yCrXIzUUVBmOl9aqoF4in+ENVI7diB8WHYYzLOk9Pu4408XXpHy39GnPvKGwiyMPwmWPpPYh
zqXIWLLZ6C4RoEXrpjY7nwR44bP6D/tHfKI41ynO9WiJBX6L5bcX89k12O9PrjFe71U+ZB5+Ri1a
VRrXmxrZ82XepcHNDi7VYq9MkVcaRc8jabJCUhqRYQUg3nhBN4NWGgIzE6KMv/p8P/tvjSnQSaPL
lsuPKXYJ03Ki/+znePEWc3bJt/+yekNzs1CLEdquj11ELyyemc3IA62V8zW/k/Q1/BjH5fUkSSrg
JQmn72V2UkGTBOid/px1v9DpWsWjs4CBLeR19ZRVkV0fE4gRr8UJm8eGY81GMDmWr3Ls2d9JwqV2
qk9Rh32K8dC8FzqigzTJogr4WPs1j1Pbq1XCJ71XTJNVdWt0IghwQBwmFasthwBAnlGrgbPz2IjZ
63VMRq6sRi7eaTLjaxFpRIzqiX19csDh2jAMldQFPMJqqhJadWLNekVeZu9OsHL12KxD5vCtCW7+
7xxGjvI/qeRWzBpWsnPrkAT2p6+8RlyQlPYHjfR1nigTv2EKz9NQHYupz19I3DAI5NDk9oc6BHPM
m3vEu4oMA0khjLxGRBhVQFc7RkFzWkVxZRilQ7YJkIpbB6WR3XCCRdVKV85QNqhOqgMOLyDRSVRU
h1ctPOqeoBSjUMWNBGNo4aeC9g0ic91DG8BA0yvmXKivSc1KP9Qjnk+JvzxULjvTA92MakJYxQ2p
Iyq+R88cIp/Qu0456CVstlyR+85V9btLGLeZjiZzamdbCihVjmS6heceeYNBUSnN6D8uix4YaOCh
2jtYPAr/prFV9tb9YoN9CpjUs/ePszlp5I0+nSgRBNHFBfY9bV7CDZUTP3WL1skQqMr7PzFKOzjO
K2vKhKFz9QLkbcXobcSkXvag9k2SoZTXan4D0Wz/2kliiqDB/e23fAadjakiL/UB2kgJRcTcZEVY
sezsYvKF/Ma2ntT7XwkJqkSC3EJzsOFUafGM0Rei0E4eqjzLMgDby8purJn0KmbcqmaNLkDUso8A
Y77QkIaDLSWHj0HbEERf5HXPml8rmjhw/DciYPtSEFj7vrXERoNme9Vw9kMLC3IUrRjbyD9a8VNn
HzrlMy4TrXN+KNuBxahZIFsv2ibkihTACscPkcdl3NGAd0G9GgL5Q1iHxeRncND8Ji6n7sUSb3+Q
GFmOkRpE40dO61HTZ9W3AjLrIxhC7J9Sckl74mtrDh2zm2mJzKdQDRONmU8RIHmm9S+gWZ/3Frzn
FJ5CMcZOt7pyP7c6iovbx84Vkeb2LifFai9BsQhGwfBSa5QjCsvHAR53bENF55H7WHVlxek8RwBS
LzmIIfNhNRl46pSpMV8SGIPsH3+mW+a0tUvv0c3qVwh6GnEQJH0pgH+LUgqDufsyirKbqYOgiVCr
Xs6A9bVVcbcYhO4QuuTYA3iYZoMX+ycakK+MZ5jA1Oz2W0IT9OUCJUkoA9IgTex+XXm89Ne4yzmA
Xpurr9Ma/2iTnX6VZec/rC2BtzJQb/d5o9jnyJ/s3fo+Rtl+Ui5HFoujz2I8MZh3nj2oStl7h2J/
O/IqKIi77LaisuActa4rFqUdtfyqqtP8q816ymk47eOBBycbj+9rrLAd+78ARnNpEy0rWQp9MPoL
lkNXH49BaADJ+aE82CiSOBYRRAxMUrVn4xeBDfH3sANTl+WoBb8Cew4H4xYS39FpTMr3gtbjfD9G
8nLhVqblU882iSbaiuC1S48mHvjmlc7agofbOnEVNjK76db6neTp9r8hj1j2QEfiI7+EnsFta1Zz
EIUgAUVACI1+Md+cTVXPAXf/FbSucpTBlraGNtB4Zvog5sW2R5Zi+JEZynz+CKn4Ma3affM0RLkj
aAuM1uyzL5CoY6mtl1qc3JRim0nR1dfkgMpVxYdKCIL+Yg++E0zbaLFJBvBPKyoZBtr2hEOAL3nJ
Qgs5mOJygR82tBiAAKC4CbD6pKjzf9YvnTulaUervekH1g9623JqMIIM3OTKx1dolrpm6ocopeRQ
ou4GPfA7wkfXonHnJKidwk24TDpupJFBdJa7PXWPtcuim+vKNvahRmPfYZ4dV4mTEDoe1LdI34Yp
xbZKzingrn1/v3AsqDQxA0F4Dh9ewKStIcionOOZg1C9ug4VzyNM3iCjXM/vxD0bLzQFTTWJx8fk
r2AVudZHWJpM+I0jXtqMcKnUtLm/BL4WqUY8CwMOkd4UI3a/qqCEeTWwlic1m3JmZKDU4k/WHPSx
zCetvjSch/jP62uJD2j3onzHHpGQB8CSfNXH/8dOEegUMgBX7BuOu5BpV5ploZLqFkIK1RfDPzfj
bWxbwnwzM24bWW16lUKEFHTm9haYWiTYut96KWf8L+u16E2LKZMQeD7zAqZ3iX/h5uTrAEUdedyS
UhFqrp4zv87S1vhBma4QRghbloaGUmLkq21kG6RdGXUk/MwPdL1ZKdKB3lTCI4ShsO3VtAOoxAm1
+azxdEUP818HXj+KIponqvC1mJmRPqaUaxWaKzy6F1wttV+aN25lYtlnMCJwV+44GHBLd8wzPXFS
eeB+OJRBX7PH7b8eYirgCdoCGLnqRb/EoCeHmqLGtRk6JMpl4qZHSacrlKsrkp3qzuXvAxFDUPde
bySg1Jjg8e6ec8S+lYN47/ySUZ/13sTnKepL87R/OzsDXauL0RnlVDK15yttVDOU21eiBSRUyCYR
/YNYXbGUe3vXp2bC7+i6xdp3GDDA73iXY3WdPmZUR89P2ABUZPa0U7odrBuuiNlcD5jlIEy+yV4K
+bEBT1QaZdth5SRzi2napH7VXg7+t59X5Yhfn+u4MKmw2xA6zIBq+18uRrRSys7t9l+ZwminJpwQ
Wg0TdK7PdtAVYsgvF1lP5MEdizjuzde44ifIljiG1vtzC0te1JnvazI+90h2DjKR6NEC2TUpVFpP
vMFz6qfkpAilWh+W8oyb8vvqkCh1FwTZdCmpg7N4t3RxyYZi05RZ6ED/PrYDdOKzVwB3ce96X53b
L8g5nm2ook/RhFSyCwVX6r8n2RTyYgWXtSl9JEXwEzd2farcnoJZ0mJrHn9RtjxSLvKlWS7OakPp
bN4LSRW6TkDwCqKII5DoiWdPh3Y+9bBWehTfq3mZBU+cX2ITYVPalL/Ou174cKi2VwgmzHin7J0x
P4pa5hk7J0hrsF6uzrwdQr4JTmNrneRBU817RDeUNC9SjHiLZRH+4Lwjl4bBoC1EqU/KLv1ILTp/
uRQq4wpz5C3ToDg/dePMeM0ef5t22wdHdOgekBLl9QVgP3dm+ginPbouZ/UfWICQTRVjG2aoLZNK
P1lVE1dJZPLPHXzaInFXhqyPqjfXVUyr5AjxKR0Wdc37g0bf6dGncs5IdujugW1zWxEvs19wd3sj
AmEqETf6FubW24YJJZifHSw794l4kkbjEzFWhzxJDtvSPghLViZvQf3MwMEofCHh8Z7YWqdS7lFm
r8DMulK1HXYKcWFHq5e6Cp0je8fC8JMlE75Et6y8XrTo9UVHnIbv+rIIe9R0BZgc3IC0wvvG1R4D
OvfPSy/f6IUihhvWybT8sMpZHTnvEfbJZ7Pvopg+I0z6DjFxHxxdX7vCWQ/kk9inY8BrQEvo0Y5k
dZbRIJ/yB/eRcNKp/sx9jPFnjnmsvdOGuJYxevrnVYZSeHQwPgIjOlozh9Sp9CZ7SzOSn+i3pKZf
9OCp8JyyzUM9X/wCNqa0FQmIaiv+ALvlnWJ2U/nS1/H6ZY2PbYArr21QCx9v359siDrVZjEd10qQ
t6GX7xw84E6QGtc79+sq+lAwnwxwNZsrCOlZn4Mvr7QIvcCtMguiPnNAqXg8DXUUFo9udNz0N9Vq
G2p5sxHGYDfp0HQNxONcqwd2pezcGvkRv1TJXnrDXcNvO2khjiHHmbhRF6LyhwO7Ekm/UyYtjUdy
fIJ08s0ntI2BfPoDdYlfH2IjR0ucBJtHIRlhpPObhfu/e6fu6N9Vme9Alp9lsw9tNBKX1M4EETLL
ZpB5sQWhELvotNhP4XZ67l1TFTl9XNdIpjzezxf247rDlWQ12B7WkzEubqJJmfmYLl14Pt+OqJ+T
nsv++TpQQweNJUcqkZ6P0pKlYodSIVQ/VGlIpljPWDAAiE4IuP8OaYwoF7G89xivSIdYWfbKjyFy
njpWA7oFQ3LUBW3bxPBeNR9bsT30h9Ya4/JR6PdCyoROamcSrWRiGYc/qjQTvySPpGn++EadRY6n
XTzqPpSgwQlUkhrcRetPWf5NDqnqGxItT6Ktz64ppihFSTB5iFUJeH9dZugqzdzT5a3/URH95gIN
foUQHS32fW5p4kUKw2juBEC2146qbX3JkXHbHsV8t+JJHcNfTh3gGfdRr0vshjYHqwxb4oatxGo4
rci5fFnJvlZFFWO5quevFlQMstBa2gjOlmIdNoofFTMCqzzacyPJY/vUxGZob9tCznti8WQyOQtW
FWIdAc/TT+trWJ/K3DgOU4kWyVbqjmHL6vifmT3UnYABPH/zaSONRR/Dw6vqDZszmbcmMwoIVYPX
wsnsDzD9nWKh0FL+FOE1G5zRU/ukQAPsvbioDeVAKc/Mzqdi+oUBgIcWGcSoo1ohE4bRxh+IuwEj
ia7XS+Uh8gCP5By++WUBomsJcYPRTs/VxeyHM86R2OlRAUBuNPgTIdVpw7h4f5FWRapA70p75Dh+
TG0uqOk+wpgACM9KIbtT3BBJNqRdOg/QhMr+juKzN2GuROj+nZlD4LslW6sztosZHdJcfHI2XQOr
rpAe/26OngADznsKQ/qzezOewOVRiZtmbuagjs8mioIBBEkH0C2FBwRl1v0d5qomqEHljmQKOD26
HjBcg6+HrJ/hfddE9iAina3D9U5n7zbX16yflCMEjOt4I6czjvnwplSTeFFNcYgWzBG6IUaOysrM
S9er+MwyGpXjrF7MS9/My/OhRxI6XiDWxTbO8fmnUVdhqyEEtUD6nKcxtE54wElj9nNVP+SesgMV
+Jrwwq1zBeTkhcTsDkNlpA6gfbuXjaR+NeIzHO9aT3ykInVKkaEJHwh5E0rZDTONyWc9VA69jrvK
SuLQ4rZdRsuLe3l0xRwjeYuaDEbLPZiepqZvaL5aaNyLcgF0xrhr6RElBwOf9eDdzGi3R9G7xCyy
oR1LlqeK0D/rtTE/8KDa+DNmLNPtX37c0TTUXKqclZIlH7iW81Gb9tXPQGrc2JTzhXuiGeoWdmrt
gJ+mhpUgQ9mUbVg4kl8N+Degf8pdWEWJQQxymOnnvKyIYykWp4vAq3RgKH5fmEt4mHNqUlMA/Tqp
Er6UtcSuQZKpBVVJ2+t9OazzD4bg+WGKBTgCn35jW5c+grLaqOLXQwchouQtvDRhTOpv0/lwvRZF
EtlMg1i4NfrrOSGkuj3PGQR5BOXeSkfhKc+sO6CV0nnGS+PxR2zn0OrC2Zq09/JsyK4t8Xa4Pooe
UlGFFnIL+2h9UnqLAkF4nhKX1Dly/kcMXJH/jglCVvLN9OMYZQrXn71JuDjuzZF2TZ28yLrIfjOk
nr3VKNFxNAdbquYL+ZQa4p8TeTRp1SCyKxS8hSfjO4OCvn2ssNmRsXbYDaDDa5QBsDFkqT8+SCk5
4/DmkeGffMVROiEOIOQ7w312OJvJKvALFtPTzlQ8yySuvZXW7Uqu9KY2LGgBwFfv8yiI/KzTq25k
3W6YAEtbBWXqVUtkRAnve2LbaPDZptW6qXEueQVX82Ztn/njIA7edX2jJVv2BO3q/AuCpqkpASam
VmIWKL3NBeAZ6ZXoocyvihBFRZxstf6xe2EDGKBE5QwhrYBX3lVJMWeYgtc5PuZjzl6gmGPMoB1n
JXok6D4C/6AwZ977zECi8c1ayHU92Gph1QfCIUcrxCS9uz22RGd/sse4lcJK0zlO3tds5a5q33qw
G6unmJSpyOiY0bGyO/HtmdeCZouEUVE+/1x3Rs6eeOwTjUUSQUJSgLPoiMZRQ47u/9L18QPsoM5S
RaTY3nO4bNUG1Zo3tZl7UWjfBaeH7ziZ5OOLNIT065KpAeEiCVxyCV0DKtcdCoVRX6bz5AoJATAG
u9VFt6eDP8e/En+tETumPDSyGVLNeSk+8Ys1io100E6+C8jie5cc4nmQvbrvHEQeG1tMerDFp1wu
BbnOzgvHJ4OkDJf1vD26XnWPtndrsK1KvDzUy6QQQpo22LsR5mVa3tHtBtMy6Omh/lIXCostlYrK
pcB/bEsuDzsSj7NT5UsAHDdyBS3QLnbKDeyI1/kQM5xyWTJj0V3ZMsfxA9SabAGXBUzf08RyyQAN
h+lYLqjR7A+dAsXPN+VBBWJdUEmVmYjq5CwOHKP/2sbEm3beimQGmZDPV4nZw1kZAqtE2b/NgJ7G
Pae9h+l26Bh3kDN4veXHH/A2+JpCd/bx5ydPIcmFBsGcnaApS8S3YYhXFoaZIGSGUvNjTNbYFyP5
HUA1dRetVlLwVbVean5thp3LE3bNFW0SCsHuTnPeA+BomTayZeylVZahpsfMVWXzXuSOqdn6Afb0
4NgGFHD9m7DiIQfLZ72ztj08bUGl+CXR4c1MSOONpg2y+MLm8Nw4tgZWisUu/VZDLngBnEP3017D
yEIkcXMl8mVHWLqGuQGVQbTTUdJBFzAj4HNRA5LWoJgIY9TkoSfhGPv7r/ql5hicTubHKcmOkk8A
Ukatp9VCv2dhTXCTv2U9SJNKexbmt9WUicE14Tkm6qeIJ0ahl7/1HFkGDm4DZPAJLk4mL6Z3F4my
CidyzaFgpGgWibHuotNSgR63Km0jjWxFFzxB2oNiF1blEZN8L1TSSDkJ2jNU3A1/yHVcu5lJkz6E
nxCp4cI2bwBFwcdSLnqwyTVYa3MvFrwHPTYgWsySjWiunbSbhqL3uTsRKR/Id+XdPEv+y5XAhK8U
dG30USpHkjSWThDtiX+C9bLInI+Z4lbKoRwLgcJNeEHdrttu3cNDYYGPEE+l8dU657uTG0mUXshp
kJdi7k4SaD+agKmjnQmw6R3MDi3Oh2ZSFrW8AiMerKaNsUbHgZCkVXjoadTW6vE8BNNI33qSEJ34
ggDiDrMVJMGQJIKNVcLAjJm9Yh5/m0ckRjiqsIfRF1PtAO7VaRBTux8NHoYYy9CtZdbVf60NsHaZ
OSvd6HtvW0F+HKyykceZyzvHXzgOhYeUVZA4sOEnR7hdYxGplFLIbVH68STAa9XhiAIrjvTnog0s
xXno907NxxvBPloVkGEy3cDybSa1zJDVXAJka3Sfpv6MWwCIjwtt0puSQkwmIFg33LkcifmU8ugq
2sxPV39+E481Z5O3dSAbpXZ2fjhA1457W3eOxMsF3GDwF6kBU6qzRio/XslrxTpT5UDlpUtZp/jV
aLCAgc//nfzuUQRHJ+yNBL656TgIwH4+xSHsoW396tiMsufTYhUfS5/IJQ9Q8+dE93Iu39KXq9RG
HSknyTtda3XdjbC6BaEu110IXrjGzUinp4/sS4PaUEvIdiwWqefw/1TzgXL3sSjbmoDoV0VN3ln7
H2G5KtYOMbc3U1idZG47RQmFyOdlEFRVKVQNp7J2k5/WYqaMFw9h6CKtUl2Z+rUA7Lzwgc6qCvJq
PgDE9OGHAzRj5nw5kUKNZJkgnFbs7sbC7Mnlx7TKI5m+Xe7UcWLzQMbGNssQiDnLAw7GUwWVULK0
/PShudrzUH0VrGWU/tXEKMscBZ0Wrd6LN4qCSpBnlHW/QJf6F+a0MGUZVqOoY83QoobAyWdpcRqm
gKM1F1zj8Yn68enAVjtzv5bdbicVz4qWkUUGXbmBHGEHq5xZI7OEUdZ4bV85OTNg+WaNNlxME+Ve
wFB0qbXSA/xC3xObUH4xta+4Lax4rDChtNW7UNCYKeI2KXdo6RJo8AgijKkxdK9ak5Gf/Z5PJOl2
mbHUlQqDJPGh21MJv0WkJI/jNMOYWKPbwtXJc+KwmEJr9V8B/OicedtcaCi7ggaYdr9okMJ00CuN
Ii5TNNZd68U5BPPYxm1HVmMkLDR9mrPiYXz5cgfMNXAUJxbBIXcuS6HCZUzaSM7EPml+JUbszflg
3YQH6wFlrhDkNv+kV9s4BLoRVNnXN8ImNNJZA9gh3qnobT/95WfytEyzjFjXkA4MUGW0I0u6pdJK
GOdY8RQtsWo1I/TT6hsO5Ht9cu00YJUzcLhZ1q8iMqR031zhq5WA860ErQD7p4X1J0o0GwcUQ7ez
TT1boHlpe8aACQYIfl2XMBKrQQHVhaPTMqNxdU8CGWFznw25Xp29ctL4e4XjxwM3lpBwS4SPkQUv
Kb+dhD3pWqISaYDjlDPR149Uj+9hf7VQPRGsabIVNrU6Wsyk9ffQVeLrdSQjRJbwMwuTb1abPBwk
u6OVuXqALdSvEqff+dBIqMl3mLq2hq5JOHDVJacIh7wKkzhcimlc6LWWuU1w4M1Nw8D8Jpoj4vcx
KNvkNY1GcPphUVUw9CZm0Zil8V95BJq1yiWz7tcK6WfU9OX7lpZ5LjjIHtoAro0DKT4Y17RNdD8/
7WS6MznwLjq9X1qxmxOLsOoDzx1XcO8hSrH+cNwt+SypoV4aXXzwFBWkcd9g9HmNyrPV7HElI7gq
ltha0xYXfWhaPu2pUO1nIvLUdQt4hUVUiuYFWRZrgLQqDp3LOcI9/hXXKC2EM8+PGtXGtEBsgSuQ
Zzb3Rogf4cnqye5dEoOr5omypjgyFNBr6EVVtP3BOnLLAD06UrZprCXBSvSusfRWyV6Q4SiXJY8s
+doQiQ3afVKgAdCGWuB1m/FKdcB/xF9KCGsHa/TS7twOxvZU02YNupCN/d9RzIdKJYoeI0ysW6hD
p7jQN7OEwKXq7Dl8ScD2MuYRRULw4FUGXneSVv3/oJV9/TPaCFSY0WxSPfzlo4hvWj59ZkvX2tsM
AV/siEQc5gtO9DTF43Hyl2I8D2EfasEYPoCO9u9hyFWCH4G/XzsSC6ZIW5fv7s3g9EdFrB9pm6RI
j0hpO87SxqtZA2Rj8F/Uyww9Txjs6PgUUOeg7CCIxufl1UlveFtVd/44lY3qtu8SHs6/trBVbNgx
+YZdNQsaECIAPtDtimQnwJBlZrEwSX/3gIsebct+W+x4QBytuY2Pf/xdK09dEyJb+x3ccxfKpD6J
GOTYbofnhbMPF/pWXwK7jfJqCPQJYK1+T9ktvgFKq346DLljEaDfN4wADYNr5hx+ccyBQDTcYuPw
WEAXoOCQcV+Ngm+ULeeA+zKguPblC9b77mf7pZLD/dBDShUsFCTyzIHfaNb4MKU/eU1Dtw9vBOY+
ONUs9cEIxTzVHir307bb0cJd7Jc1E329vANNjLS+UWLQ8pkN/48/WMPbTOGKdQvtw02ekoWXwYSn
PmH/B5J6hWl/F+q+9YCvsGOLlAHCjkcOL0uqygJnZqVbvjK8WyHMmlMmc559BfrRrZ6RnM4y8keB
Ra47npeQZyWshTu6Il3SX+P7BZ9WsP9nfnJlQry4WpgHiCqKs0NCptWPFdDWRs5dwaZMrND/c/2p
KSBBJ9dHw3q/4uwk/z97oP1me41+tjWlI+fOn2wC+B/jtdAK6I9drCRwic9fFe4ThXO9UNfkWYNd
/hD8Etew7Jnfaretr9fBalTwb1dCFQOEpCMVigmHd4eAyfTNasPnGSux/6YE44nELF3LiXNZAIR6
AooRqylqOleVb2udPqoxe8gv0yg68I6IQb3y/NvkRmvcuIlF1J9DWjd/wukq3ebm4EmdnGdygpOG
GdO4BIil76miyXEvcUsL6BxAsxB8uafQ7V9AT9oxC0rxjo0maHpYFaMAft697uVXljYOaeM1qLnq
n8sKyMe/ejRmFn917bt1xC4wUk6fQt0jg6pxw+fIba2piCei3CkHLowGCbeU08sOPim/KcYOmgDN
IWSp6pztSHL9oyQf+vnIPrM46j2GUGJ2/HZl2KG5APmqT5rKDz2WcI2qR8hH+ZxD728YcyDhBCtO
L2Fm37PWdBqWnmZAV6UAzFQ9BSafPmfrLyjZJrNgEA0JkGRFEi7ozTwDxqt2zL/7tKE7lEKla7gE
GYP8rAIcs7xbFDCw0e3tNQaIKqC+oV2VMWWna0Vh0e0+MG581L4cuS6erWYysMt/CpAlCjm9GSpY
UpyZkhNP7/fWihZUXR0i4riQhFPxwbF2wPDlovJJK6yQ0WLnMxibTvjdN91dPOwoT7FBgizt239B
CraEr/Tx654t+ycIT8ZrK9BSdHO3bG1k8PaKQcatNDTbbRw0M70rV0qdkbU8I8cAhZtBOydDHPq9
4KX+BU5nEHJRXhm742SnBLRRGly3OW9tyVA9utdDfrp9Lv4onN+aHnxAt0g8Ery7McPCpD6gumeH
mfBIcpmXSD9P54VFlXGC+LpiaJfpnXLhGjUDJmoAeyE80KxmORtNO+tjSa1pL8z6/w40aHshwC9P
lg7L/vXjAWxrvIuQUJfkf7f+mBGsjR3UdD2B4uSP00xLrvxDW+zi0YhldHEtbCBtwybi2O8k9NVw
EJXtbzmR9MBiSN5iFv7nVuz0OqOeXvs/uumKENkPm2L8FumQfo0g3F9JLYfbIdMhOO2UQgATe2hR
k+/4RhCp8hIBvaIyYRN28fbhKqkILdEcVVXBTq6HPUcsyZPyXS75NnO02mGT+Q5XB1omV/wQt4+h
N0MNM4rFnC2o0zE6NAzereW2Dkh00oDa6RUz8uTGnUApiYsVXN289/f1IN2ITKdl/+luVIrh11Hx
03ehlPBnFAO7bAQR95umdiAgj3gWXPw3GWaKe0f/9G+BCT1AWSbMXL25rKraMx2gn2WFR9PudUbp
q4QPlQjaD+5MDSIvnhgbz8Y8TBc6UdPZV2dRZB9pH6BD65Fk+nTyNgLJVgLXt5b96Fo0xhDf6ZQN
33baeajDPk5S602oUJY/VRvpzL1s7gCsiWD0MYWUHwlWeqdeY0OI8n/GguGl9SnpQwnzzwWkDBPd
0tX9aCq+2pFokRduA50qgffTw1Qx0SS8vnDcLa+ZALPqf11JyNvIHBRQLv4FoTJX2Mcvk31wAYrj
kbH146eniN0lm7scbV4ln5qacv2VSbLa5zqaoGOj+WiK0QQ87a+mr2b7ekqpjsGYNPwS6Kc1YnK1
rgXD8Ekv75mErqHWbNmhrlqZJoFsi9mv1z9Nbzn/UlYVqDY6o+9YokrQ2t7ufw5fwv6dcn8ER6aJ
Ym0pfpEFJhY1/BiO2ftpZ3Q7pZGz305YUE5k9LyOxc+v63hl4oZAgqWA3LkgIsu+z0bywVjXg3Xs
KcJXiYN7aS7x8C4RQhyw4qgttE97fR2pFZ0gjk2zS/PRacbPskd5muyyl1Luf4+EX0luDNJDkDAV
skZmjq3lGfUhRSzVjjZwwjsGCAB1QH9C6myc/xD8DDhsNMeFa8XehQChEMKkuO4XGrSrf4zEGgWz
irACmK3v6WOy2//rUVmFuMuHWYe95N6/GITAzgFnsg745csMRMIyfW5qsSO8DDfJPdEtA4exr4EO
yPdoIxO4igcKJjSGNAwJ7Nq1ysQhY+afuzv0lGtXyxmzxnn7gqWSuvn/sD8D09t02xXLEGZT/iWV
85ca+kvAkvSX93ZqYWHNgQS58yfGevlpDcX2BMHRc3MKbNCSXDvhsR9oc+h35QwGrZG4qYtFD2l8
dXuRvEkxqmjfJhrk6IxkFMhtcf590J5c1gCC1jD8mbCerdrafx/44Zr0BfrtrfHCvtFE1DBJMtKo
6a+l4sCk+Qui8VM3Ymue0KZUqrqgiMaO8xboIF4GZRYMrMLMm69YGEPvlsOCtoHSsODgTkUXRWLo
gGlPapl8LVo0zRytIkPmW5rjTPVxFYGY7HYmxEQTxF6Dh5yIftqjI6TdxcuvTaTnIBTYr2hrNgK+
4I4MxUFLIE06BNViD4MXxzYuFI4uZsMBNLNAhmia5qinmLMfUwoQwQL6whvf4H6wDOK22DLEB//p
CRkAfOvxP1fSiNnVW5dPku4SvaI7jpObmyS27XVWp9ODSoKaizYujros9xYNZr0gj7NnNNCb7Reh
LjJuBYRoI9w3GK8gAvzEsS/wACOSQdkfuEHJd7SQEjsenH0h//hC2qceMGi1a5vvNcEmliRwgqfn
ddh2SwZw18DRubWTXV3Zg47sCN/MMA410sTn0OhhkyDP3KuceSWJZgh4Lwf7AJOcBxlhIIQDzBNB
gHt+2PlZSBX4BPr86rksHMUkMlrfqgwB8niYIj8umca+sOKah1HKqhDf4Yx9RZuyMEscTxe74pme
MFsIrhblEkMYteWUGIK5hLvLnmNCXEHiHbbhszQ8uEWhOVRMkgaYmzOyrw+mG64Qqy5Tm5KFB50/
AG5SVxVW/iC333U/oKUoz2EC5RFwtY7gOhJsdeHuTCI6bIr64BReMfKNwypjhX7uyN1JWAnvePus
hX97szGecQSd3CfgGH1gUIknX6reaGMLcx0EA283dChBh+ZKGzAE+hOU1pdNyU7RAw6yMqkdtjGk
Wq1hbqH7JSGZls77PJwz99uEIJzH/nc+woaPbiCHO5XfpW9+yhBUXn7tEL2dXYxBKWWSIXPciOaL
kmnmRvcfvAfxRBv/RmM48p8RkR9F29W1H30Ncq1RztiVEdLqTVixgO0m/UmM4wu1Phe1wv60ATul
68ma5md/nCjOEm+RaNXlHO4G5omslKbLkDarz15/mbPxmZgkqD3rHM3iSovQmgc4hhbISSGeTFKJ
g+uCc7D+yZwKZnyEKX62mcZKFaWefT3Iv8aBItM722+eqD7v2kgLcB+eWRQwjR+KoNKhEBBnCwg0
49TBQWZ/CuFWY+04ORyvbgcPuJEguWki9wWy3ewtNYw513j2O9t14TPh1qQhG/mbJluI+yXMKXnK
v12n5B651LevrahHhTCK+6PHQ9nGGYuV7DbkTyomNNWm0OVkI9ZRXBw5DEjBcnJiV8bCOhZMA61p
zoSYCpx0WitJpknJLnzWB25IbDhHKmbXN9AqFRJdwY+3LZx9F9OIVJvp5ek87REC72CTDK/BECcY
Q3ZgihdAUPOZjs6pGLDPDXQrSmpzBU4Tu0k0Mfyfl76rXnwUcmQu4I2cdRNdXLNAcNuhX37244fW
FletyCroTsN6bQrLmehnDhvEecOxo1pzbRbn96W3waO4SAdTWQ9X3/HQgq4WaUVaVnn5QY1xWz75
yku6rcA5d4nIXehRp68Hnjs7lV7rdUorRP4tJryTN/BHh8PvsH8vrtOuGBcZP+p5plt10yfYukij
4tP0Tomszx93d5sIX2GkRlJotG9NrVWo6gbsoONdBv8bKssbO09tO5mblkNot5SWGVvFUVIVVT7G
Slm36ARqD6orEbyHMmflFyMChSXuI7/7b3YkJUtpiiH73bZOZVwaJpAjggmWbtCpYSRiwJjwjR7b
olyBhqdxyAOmE18x3TGhzBHe+Or/JFVH+9atE8qryTs4p4a4cnwDpK27RMnu8r/zHCPiWhU4MDWq
HRElcQuKoSSOHrCBK5CjO3ze5xhAcfL7Y9ZgSTgAqMU+Xw0z0OP8kxYdb8Ccd8Nr46wtkwZnjR/H
/ThPPNl381GRH7+meYUQ/+DnXw6QnNMvZkmfgM3ci9cioTmKsDAYPnxwWia99MeuU25oxMxrYk+9
fe1dJ/fNputV6cQXWis+KSssuK9OGvbZMqtlXkhuBYUKfrX/Q9gbs3bR6/JvqyiEToPPB4u0xGAi
15vU8MixP1Zv8vhimaAndVsoiEfcj54va+Wz1KrZ+gBuofk9dzEblPiZbtx+ed8+yflEetAi17rv
5TNZA4+KqKWZCcLFcLGTFdDtdkfQ8VMPbbbG3LseMQZ7RrR/uraDLZdfMF8SoWyr1572LTFeCbDf
wASXsZPg+4innRploCgmBA0GcfatxejbasSf/NJHuLPt580d/OyQgF+hg4zdo6kvtYmZ/mkDDEIs
LaclUH3+k+nMPlOSFsJSWuClXUaOPnIa2UuTl/2hUuPuOt4+X79lTkftOGhZZ0dmST2KjqL6oUk5
7+U72anFiW+yUBqvgb5TID+ayFCLy2Z/pNx3PoR9oWb7B5uDeZBvYyQSBGvfMSk9uWgdtiwc3SqJ
8qOt2zZ0Xdpt/IpS2MK/1gHCbUlWrNVhXvBbdkl8M37aAQuUazu3EZ0S1xpb2Hfy8m9qyWVLM2XM
vKmEO5d+AUTNHpvMmsDSeLo6BzXKoq8IBUnpgIBhq/FhTAbmv+b55T+JZiMy9vSee364r/JbEVBh
wLRM+zQ8eZStKmREA9P9+vxfCOY6Y8UZlGIYIs6GVZa1Kf0K/H0i3bTNPUfV1HHmRpuOM80dST0+
tjbKabJ7G1+55MPf9L/+GnzOpK9s3DDuC9pm6YGuRA8l1KfImVJk1Z+EWGr2SCd2sVerOulOnPqD
8gUbYnggbV+c8+b5ZUN3YuBTGhNQVkxVzB30mmxgtlQjiRee7j/i8KxeSWNVGAp6LRPNNjmEcemL
YROGyO9/+mmZ3BExhxv2BX16XNL3RG/KQkhUM5kWsnlGMdmgnt56VcKpl6zzb8Cg+fLMG/6uwd8C
/jQZ78tBJLKNnKxVVRHxD6jeQQbjPVsHytbGATKH0y9nbE14KYeuXJvC3OF3KcpCmBheeRWhQyQk
2F6NiEykjWv4qK1mTJAYovhAplt1ASLvy46E+oKVz6OL62orq84glRn8+cg1W+9hBrReXZyRXiGZ
DuxKOaz5HeuQwbt2ahxa+68VTjIvUBcAWEm30VRe94sXCHMJv3xgwjEWKAMLkW95roz8MGZPELnu
gKWATzaYZDl1bZyAY/QYKSwwNmEbpWEKLEx8VnxCc7XuRf6igoLVHNzSvqo6XN7H/3Xkqt6EhwxO
K1l6iiTYUwOXWiSdq6k3cNnxkowoR35oaxjSsZY1GW0DS7/45vaCGNZUYCOGbWbqbXDYGOQmIWO3
HtjRd4r0jBXWL8MAAfjPPR42+Sfva/QPFu+X1n7VGBSGZdYAtraCpqHfEc29tzIvaJoKCBO1ULAF
GS9wtsl75ctx3hRHV8BvB61mosXYXxfDamYtKNtJAXfRmK17+itcTEpiPpr4v0ip/IUOGf6YBkwf
M8RYGLfuVMIgai94/8xNlVeTNDxtmx9eKq54QHuey2OOEFshWLaQeZ6z0tULYpSouAze66uz8ioM
5rG0rVaDQMtnumtjjPqrAdi19zIYNbKGDPqjSVwgKoBwacUB9seJkrrVEx1tBYwEYarp5UjZdu+O
X3cx5Ldn2mNKmH5ncRoQie+muvx1tcYyPijuErZTUsxAaSwQ3eQ5TTJsGtslU03vIifxSa5LuC4z
H8jeo59p4A15UjXwDVXAiMAvjGFbVQ2IkjTeRX3od4eyLSb15WeItT11P2yVNOfdJwXffhWeu836
7A2GqugfDuftVN94TsO/h/k9YNWHXXPs/BqijhNRue8PIanfvc1U1JW3vMLa6hbzgyRfn8TwXaO1
YRatfSrJpJLFvJPK8OzgWz39eicZYLZGEIcW4zriRHAHF7tdTWr6nx8/KTeNm0any5dPfxg3+ItO
vh8wEsSAv251q9Lx3aw5e42j1n/efFSg/OMhqjHD3ElWhRso0hgvPEwei4MPtZUboQOM6SgB1w6S
nwjQFsKLGZa1KQXlG+GqwfUV4Qzzr6FTgKYE+DuvBfz4QXx1g+5SyJ40vDgVcXYt6rljsWg8JaQm
fqdqkH/UMm5ZM4Kvk6Hs2VKLStoayM6dVVMAOBbj42FWd30ifTRyi/FjrEgVON2IiCMOkwhB19au
6LVjZIpZYaujxbKiY5tq1jX9ULo4SRDEkZZJTwE4VMl/g8pi2wPOpojJXzciqZIj9E1mpTGNHvhx
7bf1FMFTs3tTphD7lXUAFoeSSXN9g/2Lp3WnoioPz1wSdhYPZ+urywj7p0YjyLLmZCrc1BHr0ko5
W6qhMdK2STyoDTaCdExTX0JGE0gCOIn9jhDEstLX1wX+GLpDOdMUE17Esenu9fI55i6SDiJzYZHU
2+SVTPiu7Xfbq2Nsf/ROVEzf/uDon9OL7bpOypJi2MGpMYSlbofIqoVay160QV8AXM7Z6n+kxPe3
+zfYBINykLa3AWVzE2OH238BleDWfdf0+hN7xHsP4Kfm2s0mJ2AbhaS//3KCE1nZYJtTrsw0HVX1
yyJNKM/9VJrlvnUvyM15JwTLdv8AJAri9JCBrNP8+HX1tbQUiPBKmR+DZLTcmTMisDjHeQcJvZs0
OyDA2oLH08EBny4FW5aRooMPb4/vlFzwdXtsUifXkiDPHRAXqIhKuPj4b1ww4Orh+cccOZ/guJPT
VKt0GhMfRjjSdMv0EWJZQ54OLre3FZxKUy7FdU0HcIbhfPgDH+1crI9KL/+Cjik6Df5Dz2k6p8SA
J1wn7iPsXnSLLhTvBAxwltulN1dcpercBiVSiHz9RMPsoyBLpBSUPmo6zWJlTP6KhZTk6TjfzppG
WIUtZmz24+5BuvATJ14aQA4y2RHXLsLW4TEt1u9pY975Ec1F9cfNobSbZGjgT24+Pl4bB93hbaoX
EdaSmCGeBLEapN5meY8dOE7YbcgFJBLk9a89DfiRTtYzOG+iZE14LkXNIkcyKa3YV5UB5dLr44Sa
Wp/6jGPbmhX8cK7ckoWFRMefYaZt8OZFurHmJe9AZr2auUXNpDXcP5c+hmZrlhvWQgIVltqcQtUQ
YkSPO93Oe/BbAnDcn9nz+MJ+duk4AsieJl4q8ZA3gt5ewgy4UgdCOTYqlJ/RrUgDBywrd1Nm70CF
21MnoHqvWX7M6zGA6swEjJ6zsagdA+JcnXyQzY0mguBvj0rcUsvXRgnyExzghtg89kXkeuFTItTT
h7tQ8Ri6KUR0x8fnpGncRRSgWGAueonf0y5zD2ganqBil4vj/cG1R3+b7lbvwrpoH5tCfgVFMG9j
k1Jz6OFnMc/4Pa2B5Fh7HJj2ay/02KKVPc6r7BDJRFIJblBD/qEpVQVmJaF5Ohsj/mug0DJ2TdJE
OZecuoa7jLcIdwGIQQ0NvMnZPJdWHdYRn64FvqE96oZ1GaOlnT5/XPLPERERuz1jr0sBdKhB2knD
VHzszg87gSjUfaKnd/1kleFgK/XIEcO2OH5q7oNjVdN3cxOT++1X6WiIgiSQaIrwPQiiBLp13d/d
ZxDqEK+abcGaq+jBWaowrWgZKVkXWvle/OST/sHCavX5zW0uvtw2I2IbABDoimB3dvzDbVaJ1U+V
Pylc6wRQCvlq2Fd6XWUsR4k033xyE77a/eT427+8onc0FRFJeivU0Q/J7TYDbIQSxYPbN+FKRQmQ
ENUrcn0G7udfLwx3jVpqG9E/g/ue9BDmwKDtW7LntToHzW1mgpRhp1xELIEN9weL9b3Sgy9jo6sp
34pHN2Rp2zp8aLwo1oqy2rODsF7Pqyn70+qSwfNJYEL10wAyJHgtZ6t0ZWwFP18ZzG/VrB1EURlq
3dJcUsgxLYuMVpocfkkfY9+Mg1OGCGzss1bQrWQaSQHS5D7ImOnqnhgn36uYz8/Pjk/n4n0Nogg6
+NitJWUif4zw1KEv7POBcO65UTgVxnVAQKlAghZrfu8gTvNnLyWp5HzUvc/IA6AFQ0F+ZC4py/4I
mF8ZJYXe4gjutbB4jDs6+l5F+173RwHP9xbPd6iumJ6xPgnx757R61sTPS05IcbLWv0jlHqtT9pQ
wXJfO1EIWHN06/N7dcWA9fJfgeHiWXeavatcf4K3NWOk8yTcsO9A/D/1JKGIOeYGNteClrX2rxax
ZePgx+JyU/zN7ipSTvIyvG1FwLY21BHsHw5OyqZQEMUnSNZUgMkjEIcP9l5O/Ge1aWeaQqQtwQJl
PCk2pwAQE7DLP/R0OfVV5RKoScuTpV61Vm5KFyMXbOXohLZYFNlCz8j7W+g3DzIRCGWbcfh9pWHK
JCBkVFWphxMV2lWGTbWiCJbHcM0GI+/p4gcIHZQqabWwl8s8vmqiwtpMP4bZB8PM0qe7I4wrpu7x
F96YGbCnrTCGd5xo3mt/EMsNfs/SpLTXBGZcFkKitsZw1t/Ovyhd0mdOJzyXxJMi5kBQl1RDKXe3
o/08hMVweceRk1akA7kLNN1MlSSorOKOpUf9OjqE34ij5OZd05uaaTj0ZH42dQLHKK8z/eIg6neJ
/kwNs2UB9o8sjFYW+TyI6WuvDlOIs8whMDmMnoyDDitr41xV/+z/VyxBWhEeeQFc+ldukudO3PsV
4yHcRzWrKvjAf3n20FkD6on3XNimVuVbD7jEz5w/oeD35T1mYbAwtsQxCpGgofX4sg1l7akadxRH
wkKniohGmvUZpX3TX/y3jPU/QqKULb5JDMDZmsQwlcNo7C+HVDI4gb9/NgGN+NORBKX/YMFpiIe7
pQ/0VemRNvQjCYMVyVU4FGufbJJ4dGdpjPACc7FbayM5QyYwvQgNzNWWQdSiqn06e0HSuyU/ur12
xAGtDYC3KyVGiAQByg2ExgftzAbTrSTxBQnYQIyDs+PVofrSqn5A8Ev+MCRuqSTaGFDrqSWL1AsH
uKxSjAGCFYhK/S9EuiWYSAVu4qLFb8+S5lAWr/G90duX91WEUlR0pJ8MeZaFpve9SEE0PqrbRHO8
HIU1K63vorY2i9+3PJk9CGkEjljpz0DKkcDhbFcjPPw3fn4vrM5BR7fHIeo+gxe2dChT3su4yD3D
boB/eAut5FoW1DZSOR96CTAst1rpBrU63VCUCBIxZeyA7+/Xeo+//8cCS7W4gfn6IYkjrpklUgZn
ScABFrOeXvUtR5uUSxHBbLsTfuKuBfRrmZUKdbh5GnnVjWsyK1syT9b2r8d77iGaBFyEzmDyBZn1
yeA5vlKY0zRDq9Xb1kT7EQK/g7mVSCc4y/uZJdRQ7H1ixI9kxeA2YdtfJ+6cuAwEukIgsIUEBKnZ
ao0KS6ukbfRXhMB6DC+OPygk5yptI/MIg4KOLktitlfUnanzdhl5aPww1jfrd465z2RJtMcUxAyv
T5i1hJQJP1XmD5sg0FYwMo72m4joE4GFkGhYu0d/AtQ5DWIQ0hNYD2qS2WXsw+d5kH3ypBgcW/8V
toeiXbHaAFNNmoE9wpog4x/QgfRvKukb+xVM+I9NHE4te68F5rcOwpf5SIK5y/zMdahu13qgOdSW
KNWNeFImf+Q5MEcMIqHbYGU/BlZiIp/OLsNAftbnbS+cqvIef3jNikuFVJ6NQOAN21143go35VDh
xmd3iO4GusuBRkyutz3vK8eKyZrAhFXzJs40dTUUzsVZ/Jhz2XxO465hxdWrfb3mzvDOFnrFhadN
j0BtmzNZ9EUSB6aj+qzUv4ir1fp6gLk3Os9+2t6+sNVeyUC//rQFf5n1J4OpKjCArVNOCNMkfnwL
xASNgecuBUdaQGhCvEt+CdG8tq9iBquXcnRtLI7Flq9B9zXUaBt+HKLo7hmMUTVNaJ/Yg+axMTzm
QgcNlNJKVd2srJI9JoXlzbGkkwI0FPbfBSARLE8y7URzVsm+OLoXUL5habXiAj4JyrSpm278Vq+X
Li/DC4R20s8NiXsRNgARDv/PeFtrG15kK74PyNoKjdEOpSLZ5lTgkqoQMRDLhozdf8vUNfi4tfUw
y6xZxxo/hsKOrluUsz4e7ka2f1AkmHmhlLKx+USRgYtslC0G4sfCO47VIkWTJtzrw2FHva0i7wN8
8fjodeB/woUsj7R6X7CCRJmFnO8GC5+fPTQMKKcbhYTU7Cwu8PdUbuiBa4kWpUGD8SjE8U9yc36G
PHDcr0OS92XxhQhZglBF5fxMJ0gLWvWBytkTEmfUhYcv/WNIjf0ADVDhW7oAf2p8gVMkGr3EktCn
470W/NBe0jz6oxDC7DX//YTUjh5El2gqxS/GoLZnoKSFQCqlMtLt2uimpdCpFgrdRr7ka7wsvZVP
rDoKt+Ns3t0e7ZaS3OqeKTa2zeiERvYN6q7UeKgVuIIO+je0C4YlbzP4wuq3qRPGqHIuC6jmjUnx
yY08OMbFMcj92DAzcHxIN9tHzZkJGQ8oL3AXt3JRlOJ6AasgDOq8v+THmBnguK88t2nokIeWdpLO
DaBi101Y9148o0SNxbvZ0sBoL8cebPWAFMrSbanwMOrGEktXGfER/Kls2lkVOcWqsHtfjULQSL7E
L6U7dIVFOpFFx3OSjSmAp9OkAspMkfbfzQhzLijSKGFiqvDHK3k1k+iyJvn/uvxNxlJYk6S2Mekd
brOtbBYHAM7e2kIsg/Exjiw3FHtkBasmus7d6WYkH+Aji5AzhjsYdw+Mfq0fZTyNgW6S0jjexCPG
B4deHNIb8+pXtfI9k2zSslxfm6bTeUufBAGpwLWA+Ngq47xKyTxcn+BLkRJxDv5pp66s9k+uF6D9
o0ZXOuW2PMAXLrK4YyFjqjnYVYnSJKwYCYFi32xOELD+E8JRATS6bL7dawHWDeEsqK2lbSdF2+uF
y70RZFe1Pdps75sKfQs0tkzncN/B5rvgB0uSwHziKv6v8ERn9NAICrLlLqmq0UEbHQoFVp0srvou
YliCeXwnTrpE9HVajvuzWEBZEFL74N/qz/3inflk28hAJsQ7H4Q+lpjqdVObkRektQGczop+8pOr
InaxHYVlrr5GHu0GBoJK0rd+PyS8fJo33MBDh5vfinzZgaJzwhP5rRp3VRE5E/T6HwjcTIjg54ZR
tO/T0ZRGIPvWkTcOiPMdTSY/aqZWJUcM5eQ6NJj42D+LFvLHcDsRHzDdz0m74EYBx3A9lKGeK9n2
0NBLtzGoQjP4C/IFjk0vbuBNZGYV/Dr8RG8IdJKkAD0cW5Z0PvhDJSkTohMMmV39I1Gd+NRVNPqu
CLcYhhoswC2gvsMZxzTdYTG0TVfb4nqhth4V0BIleHw0AH9yG4smtfAtB+GZieqYAFY4ylKTPjgH
BVWD4dgd/dHFiGCwCv/aD/YMkPTUb81abyzj5V2UtxNpVtNXj+cgR4JqlkfJRE5s7PMd//IVRhJS
WZ63PKAZNriHrwnX5ZoZ3D1DnuCYbzdBsA/Xk+ALs9ctCr6F1tIJcDsLhF0jXe/R6Ig7zAZmDXP2
r569BVZk/ZtxQFKRwxD522kJQIO8ixitkJuLllnht6KrWt6cLoCxoR5zZyWkYYBwNl2BrL0UyV1x
sTsXVN7rpGMZaB9xYH8S9Ey9DCj6+t4zjt4DFMLGyFOvs0gDNE89ccKUYpRfRL5f2uV4a+/WdC2V
+yqUS2kEGIfEeGB0dWjfCmWO2FfveHgTprcqr9yQXxsUOwuItM+g9Km0VTAlHc5teTW+P5Kc6n6k
D/x707Xs44JNzQ9VnwePpKwVl0/oyzIUoVnBEliKKqGrNs4XcD19SGmURBRTknZviQ8SarH7WQqf
Y3Fvg7DFiGhQb8sHCy5Ro/V8OFfCZWHeMI4S0fx/W1gfD6eEaTMUJ620iix3YCZW+P4BBb4ItvPc
acpRzpfPhwEWW/8fGMxFK1iI1jFZZo51Ky7SXSsNj4zLZYrHxgbS67c1fSMJqTMr1hD1ePULTUhu
jHfCqbn/xvQTb/BFD/ymdJ8Emt6Tw3VDjOfXOBunaRYwz4bqjy/iudAK+Y0Dapybk644hfa4JxyK
fcFfhCrJGQ/wuDIlBo9w6DTJLLu2e2l9qUP39IVoDAJeOh918fBaxJDBYwa5kp3z9qzW4T5rppdj
IXZA5oGADQwyBAdx2nP9QKJXGm/hd4MZsHgcQG+SKCU8r32nwNdeQMotMMpqWH25VckXOP07KeOe
UCH8qV9NtsWKDfhL29rt2TqKw1vaxtPG+5zBECdZZ+vyfFSM6L4+6Di/4UxZwQiNU+jPquk4bmAd
jTIfwmhotHF92JIecvlP8uXpdAqyfM1RihjjtNDNcNZrrrYYbeoskUD8v+SSvYSpus7L2o52aq60
q4Uuyk80jL+a4BgW0wSO7JrywUzTz8p6GcbWo9OGdZYgBq7nUv9ZTG3dxi4vvLJUvcBHnsTIApqm
ezrwT+mrycONq+6p1yDO178umnf85af/3nP1WFFJo2B3FT2fGzsapiNecZDWJA4mYpPQeB9aPaBc
1nzHMS/jXpRMjVuHOtJgnB9BFdK4ke9Co+lJUXBhq1CHEJQq5hZ00gmDGOjIE6gnfYizfirchvHT
sTIRO7JUQBeIuNBmrZFTdjVoIQOz/Zlg4q9selLKG6rasYOlFlGFHzu9Nh9KN1ye8+gvB3TGJCCK
4fHJRLvQExdnQqUJB48KAcAaJ1CE8CdBbQEodu7JmnK6F5To7IQ6tKKdKCgiCzXNmxzYPRftzq0Q
q21shTxZjm0M1gMQ7DgZbSUWAntZqrB/GFHbxjrHUyNaBteAul/esfDtu7p53ZTs4KT/bG7VLYb+
O7KMf21k0TXzdokAWZfx55r1J5X4T3mRsAn5KOXwUB6jqqz/zXzAJqih8CH26ZhCrxJdxvBz0tJU
MNjDDePq49yuaqfRNN/JQWn3VTx3z+1rHXSC9Y3ttEs6ly0Heko+FyNtEf3BgHR9hK0cgYlmK0gZ
irC6HP3/xDiNR7oNh3PGDpeltuGleVhVTe3aLdFi396VXFBJ5GhTGrys1HkrHWfQ7ZklTfK/Pgy/
bqDvL6MPtRUnG20jLFTWSfJtxogvnWESJFQzRyjecYIAwEUsdwjkLO9bWcUG2EQSHiehORnjqBVp
8PH/zPH9iOv2MoN6C4XlmYFmNONhD4XxkQKflig48KsQYMEkTjgjN2KBMf0QMxHEnbD8B1fkYTkB
8zXkNUV/nPAJq6s/a/vXIQt5av7ky0mko5LZj2NAcn+2ZhN0wDazCrdTFl0VTxQ9S7RZZv2nUHQ6
3aqcDYn55XJEAPWZO6tyNW9CMlCY3w7sWmIJRrAXxW8KmE6//GcREPt1cPUNAln1lJUIRSlupuQu
PEsc6jK+ELXYiLPvr7TRs4vnfwyAxXV3NHJrQrk//8UAR9KSwF07htDSExmD+zHezlpo0MH1blEx
0Dsa0vq8z0t3D/X56OIpk3vnehGMUKX07mCOQKDeIKC5GV4d0gDxKLHdHSX12vLZF8abNJxXti9y
C9p78cWkLU0RFAYEGsGbIaZkB/xUueEx8uFcoooYsm9xn6dxmmtudXFYw725UW9RQB2gxmH4p1BG
RvAcn5NfNb2sUMfCkUZ4r7OVEstt97QlPdjNPDKAnz5I6ANSiy4JfCEqF/RykZ3Fzp56GI+acncY
zidAcrdPgL7o2ufcKbnsWHcu2VLph76c4HxGSVDVU1bVNoxZsYYIHtkDt5KgsgKLe7dAaP9vwS7M
tpEUiKaqFddeTi1tM+3T6RTwfKmBy6tMMeqGSh+L3Bb29N04XGxXISWbP3Yc9+0e7sT9BYhGzXeu
EJ9r5GISYI3S+Aj9oTjqPdal3avRLzuOM7DUbeJZ29seXlRMZfXHwWR4AXJWX1Ro9e9Tw0lMNQq1
Ql2jF9b/BDNB3N4GLcLs3D8+0jRtZiB/0EAJDL5nJRoccrJXuaiYfs+6yAH78KZCiMfzuTh/ShWb
l8oZWcTVCVWtAMvnzY5SEKF+Go3HIvFtvirmlFUVCuK2l4I2RLdSL9ot+9giVa7p64OlLEkXJ7Br
g3nQbI9KiIOr2d6GsdvBd2G8vkliYztVGifzuwxlAY1jmIkmGCKoOJMWDjPSyTGuj8S50cAuoYMH
vb9xgcBcupHaoxISY/1947zrury0iM/PUVzyYgAxhuqx8RN2E/q3Czxqau46R696CK8m6+mzVZvo
CwPUK2EAVTxDPcIuBBx0x/OZFx49lwEoBWpH6jLRBxkhJ6oCuNvRJ/NhEn48qZoUTiJ7+2EEFi5Q
0DqZiTIbHQvSRgGdXFwQ3cIUbl0MC4BQWXygHclfSKjLNdzN3ZySjIIke5fd5HJgssM5rs3pBRNO
t4eaMUk5b6hIp9VXFjMVByPomF06PUABtolIuLpm+nA91LTF3gNW796YHR2g7/GlgJmd5rhBrTRK
hPtVchm0gFvY62nxAiaBujnxYTeshLZ3PmyVTa2ReOMvUPGNcOx00US4kFOvTme3KRMKGScW89ut
w2xoY8QoksJkuwaFL/evKcnNr/5Y6LqGOTZfjMRzvw+ATTQEHR+vZMrawzBDtg4jUGN/zmQfzlzg
F/riH9NxFOAuNCb6RckylzswaWkrt9yXraB9g/pi/q+ERMR0FwN81FIfUb26PkKRBIQyOvBGTTHE
ipf0dhumBREvdEEvnd3l1nEP06aKXD3MS1waX39uItvuHwtmEC9KUFAEItyW3b0u9Js1RifPeTx4
wQwliCpx91OReGDrYP1/Y47hUkYhK1uBhN+6oinfOVpAhPXGuI06b5ObG7fz7jToovzwseIUMukU
vwfof5kSTfd/B0bw00X1mfMePrLx8WSwJVZOouZDrnnlInqS3Ra/2EDT/I4CdELH2xcUPmOLMzlN
dnmziYAFDOb/NGR4zuFmsfVM8mYNcxu0fnhBnDEfPOekkmc0KTGVLor2RS1/mvCgCmoRSHNT7WaI
lNJ7uuY9OSO8q2Vu27ysYXkJkzbI9MWm4DhLR/BqOVYuO642lrYVq5pF7ADOCI64LJs9ONUiL8UJ
0Kfyk6Q0EebUaHOKpfDg29bKFLtP2s3RUvafWpiy27/xx+IqaVCz6LZ/YoWn98qDsSEImkVMQPVm
9xxU0YPMjNglu8SsZV+TIuxAHc9505RYoFbinRGWzAiKIah+z3UaUAIWEE9TWTWAVTdWLyx2HpBK
umwx3PJmPdRsSdYf39X08HgToy+JznPYCjnITdVHVFsptiJUO/DTmY9CqPwxp9plz1x+JoncVhyg
EmJ5rDE6QeYGo6Hex+WwYRVcFJ8dfOZqnoSDpmGF4/5+OZix5tEM/QAQYsU7cWFmiN5gAPcLX/7Q
1vDADipQgzxQ+3wf/aGPl8NHZBZ4YSEwLXgB8FFUkt6HGhMTVPi6jx5c7fnjUsISsJtxyVfPNMr5
g+ftfAwgF7t64+PZR1uwj9Cl05VGvmhqxO+rUlrzq09uVvdWvdvcqVUyZa6SejY6wb8LOo+Z1h8V
OZZaG3WDisbn25lD1rCh5ApDMzjPsT0nNzE6H0MdmMHqju20c3cb7z42Zt8z0KdXe0+Iob4JgnZh
RpZ8EbFoBt0YoZVanpqeSpBeaSHTt1aQxKjFzz2ZqiAOfrbZ0/h6numSvHkj1z5a9PB3PNvjtqTV
HrQ0eGUE4TGv+3VWL0dEdyzDK79x3s5cNeTqWN+vbus9k3KspFQAdZXf28TRn0Ni90BbZ1lVKXN+
NxmmMvYMBZXFVNeZbsrlIa8DrEMlEQvgpinE5F3Hsxy+fAKJjYhvU0/U7H9KFRYKa4fpODzdFzOM
sOTpAOJojQmurvwcZTZOM2pfHNrACbp3SBJbDPCjtukugRH6fk8XKYdZaA7BW/2IrffAGxU/JD7V
dC+W1tWLi3/J1aqIBqaN/AshgB2+sKj0pXQdtKbfATXDKyTSwnvR/TTJfxfETqZd2X5cnVLS7Eg8
T8fZuHXgelAMs7/2n72aUcNJD74w9SfOM7otGO5XQ09zb01W/e/HjM6B2zgtTK/KY/WP1wBBJbH+
PhktyAmnqn8CwMjle/iFpQYzZmohC2Bppt4QsdIujoeIc7yep7btyo77bC96B6FSx+PiRmpuOuuY
7T8Gm8BANp33gXV8nDvlBpaBDkU0Y47pkYiYMhm2xiJXDrigb3eFs+sl3KeIJNSbAM2CUx8PeQ0L
Uvsezrx+9MOKYxg9FkrARY5ASZxReEYq/1NlpiJGb0ghxP1+cBzpAy8XcxpQizJlBUch3EoV1JGE
ZIVYwimVDsyNOhrazKBbi5c4Jnt45n+8/FV7AuwG08RtGjWCc49q54KIP+hWWPfhUOWqrYuEdCIm
cvumOP6LDAQ5pT9mnma8HGb1RMNsfaIpjMIiohy/d2KL1TfoaKfxbuSKVfBRWBwum1bC694Wgvcj
tuVgZpCbSwcy5oc1qVLRfJtGezG94+mffXjBRWAYhgjzkTeYl+fy1UopPRBbOTCc+XE9CO7mjBCW
5kvdNmEfoShelxKqXY3pFLHtrffZ3ASjWc0U4KrNlEKpFzoOOSnmjrhQ/lUhfJ/pxju0uFMek7iR
nV3IiJ/E3Q7zwuRxNIBXfaRGJm6O1pO7EGTkzhI918Biaw1Ydz8RpO+EWx0QskZU1PN0Sq2euPtB
cScSvS8Y4IMui5w+ISN0LHzHi5P/Ja76xxaXpQ2djptk672Opj1S7o67fkfGQ2FHBIWacWDxc95r
RDR1DseA2xNBW2n6dDV846tr5CkUTsZ+8AfzUQ/ZJwqwQ/vwHoa+spNc9Yfjqu3ldIGVRboF53Cy
TCxuEBVGtUFHyPT8fX4E9wSCVJIadD0r50o53BZ4SkoPJZYir/AFn2jxNOhP6Txw5IShYlWvbDN+
cqsW0I4Dd8xAraeAesUtma1BkFHgsaTi2uva7/IZAf50oeS4hsKLI6e7oY29rw4CbMQsMeOFQ4Xc
5qz+8X2xD3+dUMheG9o/c2Zg3LpVVtO1OESc/5m6UcyVUtznJ5QAFaf14eNNI9c65B8NoOMeo44j
usaQMGRjq4RybPbXFhX/jN7rLwoOcYYFO4SzoNBCZ8fdMvWkwFj+rMZi/oaZhIA/CTAkLkyj2DOF
6Q2yR+FWU89YIYhl9Gkahkp2lUf2Phe5ZictpmAAGngptH7NbvPn8VJ28F8ad3kkui9KQjs5ltNR
6J1mpi+qHoWOjrdWAPcropEsMLHWEK8P7b9HrLEEg/oc2HytnrwAR+OTnRQ6TcBXPUCSmfaZMq5o
Rkmj4crWYf9mXlobu3CcWtbDEC1VUjRWW3jfdI0n9rd1i1IakUiPenNiKqIGIxUwYTW3J7fYpvsA
xWjEgM0QJAasbxxXBVrvDXqWtrIwPDZEk2KUnu3AjIL2Qz5enFQt7Z9piU3wRA/YM+sS/zCtWrqq
I+aN1YJj9HABEDQjnfK3OO4lrlZka9rjtKRHjKxZfpdeLmQyBXB7VPMGynxb0oIy6CTHZr1G24+q
hwAkOvX3Jp2FZqi33fzO0Q7f6+9EX1U9wUcoS0mRdqAEk6uZVSEBogIGHYiqa2JKyl2Zn5Vk6le2
Z7P5p5PelNTPPvOmCPfgaWp2lDhr0rgvXWUDu/M5GeIWSsCJcJJGs/M4BOtFc57tGYyenWi4tazd
P9xfgMi2nK6XPp85G/nfXm2hAj+t7Fr1yvlFZxgSbhA/gjwOPFJx3SOfcwK2fUFvfLS9TqvXzh12
8xaO2cU9h75bk/jKbhPMA83ps6QeSprKepHIcBlQFS8DiyfuEKJUarKJkAG1CxnSanvpSRO4j1o9
pxWDWRdcPjqdk6rFJPweKmM/p/Tv0u9t04sN/yZBmIxy/IEmhqCIZQZ6WfAVgKtB7eSgdr6afgT4
rnl/jerg0RZh4/Qjkc2zv0fVD2HJOBKJQvwZP0M7jSZSIb4mIrHqvEWpOLk+jMypASA9DzvXnSyy
B+q5QawPwWJUygFBLfMd2PsEevCfK4lxI2hlfEbMYbRxizPj5xWmQHnOTbD3fRG7oOLQFgPN6exu
14Ixuy9BMpc4SUZ4qkRqWxDjvJBsECLvP/WoHxAdlCngr6dCFXqdu0Zfh3jlx1fjjQkF10q0RerH
cSly0AFPARQjq16OMCNlF4Uf0UbYqv8n6Xf1s7elAGvT317K4Jl8fTjQja1PtuJKT1hS0shGH9SR
/jCTLV4Vz7plc+UvjNLxQHGJzo2djZXHw0rttbqgkterueiNDLbaDMREczsaaLwdFLWph8lulZUz
F1CmTKHkHL75+/4lBOvZrg39sf6XseABjcfiashIlcWhEDTthqB8rUcu2eJkrGPbGvkLaI27R3Fq
0tjbaoW63ogqHdiXwArYViXyr4SqUpyh3BdSq1TgCd9jimT0ggsJYSiBKM72vjcHjXMhO8bOUfXE
q9NH/CA+QqSKTH4YOYa7RBDg46sYdx+1gELCl1dYbpMBURWOTfVhLTQ0tlXuk13WxdfIYja4tn9+
K67bySfrsp2IYPxKZ7QPJaopgbJJU6lJRO0JlANGYLGc8JAioJoHe3BG0CNbvLGrPBUf6lw4fWkZ
kZKmgggtW9X8P4IUNtDhNzHoZ2/lvMutOLJBwc0ezsa0g3s16LkTsqVsNKmCYV1cPxAt7rrVhMUn
4pkCHT2vAHCSuqk7hvEgUMqpWDOOZZIJAr4z8XSevCnud9aGyHaz1LwUdlR6oUKr4xPsH56RqcKT
ZWZYngb44MFIZuEVJy+gjie/B3tB2CMVlysmWh+O8Ity2zWu1VZe+d1R3d59Ox/l+X4gcx0A23VF
q/RabxVh37wSOeqiYQmJLuoVZZe2t4RDIOWr9x2suxXZip/tHlnUTnqDyAfSfEgN7ilqXrMBPPVu
Y4PLiInCOH2zz4qbDMb/9P9XTxN1cpO7lU5Zs7j6/Z2nSC+UXmxi8cCe63qS8+DCuF0PfFOEg77Z
iHaNQp6B9pj/dJv5iIJTrCPEv4V92O9uAVdrQg+/O+1NYet/5XdyJZ0ovSDkdhL2F1x0wL7IHkQn
2uLiTkqkKDuO9KwtRzOOLgBMSaCEThJMNUY9r35X23YyMTUchtjJG5fh0GPMxwQz/iJiz4GaLmCW
ZsHkPUXiYYc2buvQRXmW9Sxq8tZmKICY0bpKu/Vy+vA5Sr64ex79435+fB8K7RBxLC+lwV23JI/e
pU9C+aG39oZeRkCZmmH8RoIn+jYW7M8BmbKV2iVmro9kxMg5DeyCmt0jiDfOnyBTMeR/02hPc6hb
QATmCYv4SqhkH3vcLAVJjiPvjKYKBVgPyEa6NXCM/4QI04migf1lyhz8uXIE3k3CKUURlEBZeGzU
ZpBYEiFCZHaS/4AlXLfi56cyTvvb6L1RhM/LggEp/UZwhmDW42KvwXlYOpO5O51Gf0/Y1kO5Dnvt
+ocqpqcOfnTRdemC5JJdHsNsn9zTPmjj6NRXsGUerkdyZwr8rftNcXRvRU/wUhUlf10NxaLUGL7X
KYvxDOrI9a3PunbUacWVl7W531GrSmiMFV9T/0jRIi1aaVeVPaEGyQzZ9kI18t86Lf1kWvGh6u2e
P/OIK+B1fgi5sCB4zuhnDZ9WH8C4h3gtrpogBxKDpKWm8lIGigg39D+9EkJuA5p8sI4iwnGvJV9N
Vw/YF7NEo9HZkG/Odst33+iEax8Vbr+jtphyMPuq1HHskYDoRwhXJZFpPPCCm+FUSQt3T/GrQ1jA
To0H6CQNu00Riouy90Sb4qV1dHIJhwJWbGzO4RRWtyHtog/eauaFlU0F+blCUVhoKxqwSHa5WYF5
4mt75HRHy9+4FbXzRP/TU7jwPZtAuJJos9H7UC7GC7rLivHuPPKC1lpUgK5/eAnngTHxhhY/lJym
oFRCy4AXPhsAfnYwf0H+vpHsQJyCl+SOdrJp2xlix9PQuT4B3lWOrsPLVJcUV1WyicgDQaAoRJaZ
pZGNMJu1PJny7gCXxRlxdMvqPy2y+OxLZotxGIK1znc0lG5JWngYahNOnCCqn0veVWpeEQOrtJfQ
T68ZHmHpC0fGAb1KyKgyCmq0ou5x0abF2HP33pxrzog8FfgDrNyPDCcVYC5xbwH9hl62zCyeWTFs
c4hvlUnklejXAD4zzgsemtvMPcoYhRlt6ldpvYXdEVlsi4SZheb4h6j313WlY5Gnhcve1M9fNQMK
gWj+Y1JiThMaYGL0mrwAGzIWgYr+OC6/5Lk1LTJ2vW88f07bznHxGpch7ueQTqYXQFpn1ve25AAY
8DEDrvP066LczbFbHsj80MKjCX+tbfxe90iZcV6RkPhcXWc4TSH6w+HtJCNi4WwjIugaK2m2rWv2
c7jELgHog//+K99V0sl9soshtSCYor8iWxoahiseGi54QkDxYbM72ClTfWg63mMr/yymyQb13Rts
06JcXeFutHGHtI6u8LWDtSxfkjBcIrUNUsC1RMuGrDgp03u5sfMV+4jz4Y/JnKjFKeoCackeSsoR
9GrjIQw34xZsnmunTBXcTKITUnpZLv2HgvcBJtYgyEjjBUfwTg93ndDYUJvpOdfWV43SEcP9uTru
CxxqCrMWUwBjko3wdwj1RX7fhzHChtOrPjRgHdMA7L4cr6xGzzs6ml3betc9X4z/VmQbVcd5AZdQ
S3u4OGBgB/5F0sJx3GlOJGzF9XtNm9M0617GAzoXe6yMGUXKbXq10q0euAZvdEtfXFqKAr0eefxB
fGGAAeCPv674xojZ4r5Jv4LQ1eaIHXRVqyb53X0ZS0orGkKFKbaq4soHROXdrX7mylF2pswMgxgs
+zt9/rrKmiAy+skzBpzB8XyPfoOQ5MsRvZEzsHUzDjkPXF1AZnqv2QbvJPCzgxB8G2QaL6nIURMh
ZDanSSwA+IB/poMi9ovSnBcJOV1l+DykW+mkES2zIJHVAjY5RNzGlKIYst0Qo1RBXYSS7IYrxG9k
YvOw4XwSLG1/vAFvS6BnJ8nDZDAmhfJI34EZ7H/7mtL9LQWTRvxxcb9MgdT7rb09eoTS+suNarjL
dplkkLwaA/MoGRoPLRos/wGnv9vDpRXA01GWHHt+A5maRfps11dhgi/E+97zG0nPv7IIvT/FW3M3
GqEg1u8cc83lWe3n5obXr6atK5EYjaMBUbvS6pUV4dtNgZasf/RUWJchO5QcjmpYfqYar7hKD2nH
JEAL+wM++uuGuPHLv2T7kK4QKswYyqVGhDnceE0fAji1nMCN+c/5XNO9sR8ZuW5fE/wEPbL/66i6
rOXxBiJLFWQp2fdlTGoR0M3aVzKSSW2lFCXOlwjxyR/zzAZz3u94375druuMJ+eGJIdS9/DgD9OO
IcuCLOa9hbQwMQi1I54o1XwBX5q6W1Ubdy5pYYXKTIyd+Mi3nspEyoJo7b//Jmo7H54RQC8URc/O
O8lPWrTbYJqCouBQ3SYbKz+OrSiSuHC1S9AMkTvwd/3L/CXNkGxwNnaf33f9VcKG2GAhFT/onjqP
DZ+QD7Y5bU5lcE6Es6hjPNrxl0HrMVeCBRGPULDP8D3+a//ER4EGdaG86xcs4Zn/2bL4oCYrFzxT
OJw1ReAoawiSpMhrfeVPXHMPfi+60M9m+mVHm5+rKSFat4dqns/uLBwC/qQJ+PNecV9+122vHvhY
axivYz0xiCPQBUCDhGGzy41p7oD201dPLuVLYOLXaGdcTqdPSDE+xpEVpQT5/bXdk0FOq7nZVqDr
5Lu8z6qz6rj1ADQAsqNUpss65tdJErmMcRIpQbW0RGfmVds6zeceSDxxVTo+/NQNc5j8EgpqxWan
P1rpn42j02yQSLWuSPmv9TRvTZWjfqlgX6mC0vDQj61+YvLICf1M0JlXTvgCuHKI2r07cW+Lsy2x
XHECRXBMEdZHgIlxuNpYqZyXrMwGwfiJGvW3nPLWS4C4xIZ7lmM3f9TcJ9di3UAJlkknqbluDoHM
bNoI2NgH4TqaNfZ5XwV88rWE3m24GVZ08RTWJ27xZl2IQLwM4t5jXsdakUuLmNF0NxPMYY3wZSsb
Kn5GHS6pl12Z8FYVd0RzzXiRXCy6/UjalawRAqkIftGgKlfNC9EjxLoOZkwlro1SXLLns5MLQO2f
8eOk8eTvzTjJLJpMnnD8sypIYVknArC5ycIeUMf7lDsNQUh1Uv9Br2E6+HrQZmy3sYD0jxUdwN1l
CNwSqbNjeUSH1lypTHfIWgsWZnbjVDI0iNS6NHujtJrYdBVbA9xjF04HQDgPWKYJXYOfYuypeRRZ
7/7UlItRlDq5NuEgXcRuL92Btnjc/S8JlCqrYFAXbXtUMiuob6vik8nUydIJFnDUkBZLfvyFZ2P7
Tg22WN8alGTwcJ3uB7fDvGf4YgxGKGREbFyDfTpdTTjqzmlv4QRFNIoJ7mi6ImLPj5HVDmu6Sb2H
4QOXG2bPCi7t4tr+DE2zMVWwjRWRAmSK0Q9Ruzi+zuq5cDYFgOahLtT/yYxATbBfqN3l0w+eJXVU
qe2Am/PIeSjB5Evf+AIbFLVmBr00PcYnMPyDxICXxl6rpdjI2HMj1VsybB5cW/V+ByCzCt4arp+V
LnInV65tN9OftNbzOLsASN1nbgFdT/iqKmseXMFsDA/jW0AMmDRQtzZvR6Sqc5Vp/oqcR1OWpaxL
BRJfF5La3gS+424ghgsor/ZZ7hFRdbOYXhuxrFaaxReEouLh7YaH2hYMAX64LyNq2RKPD22vLIJ2
X0o6z/Umu0ef1qDXBMrXbFAr3riNToIvjqlqxe93A8tgk/dcuGSRgA3nyzqOym7X4HCBBtLgeZph
4zdcJ8XgqZlmbcuxG56k3qlpV6DsupCvMnIh8WU8y0aHlsc84/CTA1Olez/I9jq2bjF0Wp7VS+uI
2Mn/kGsw3X+QxeZcmCU77XtPZ0J6AOb1BxoYaRtbPty19YYG9hhw3lm0Qpp4auOkwasz9LqhtF5J
RrIM7VAUUNaWkjovgv+PWsQGMpq4ANUCCD8hyYGHPQcG3aJC3Z02M8QX0WvCMWYf1m6ye4cuMLZK
SG8gz9PFuB06crDAuKqTnT6duQntVrLlnjKhJSTglT6OptDf8L8ZYAfTNBMp/W5oISHyI83a2kvO
gx4Q32NjBAUscjtVgD7htkHU5uJeCZVpTnnBT3BYGzW/UncZzwN4B0vqoTfOJyDrKa9wsn2T4/RA
X50R0IuGXL4nIPz58JldZIrfkgFqR5SznWh6berJIAfMyDEHy+mbgR4VGByvweRIf6ImvHxGnFTq
gZ7lZPTru3hHJm9DXNNdRtYnAkuMGKj8sp3nFqTlhk1qAJ23i4MbHRdOLSErlpseY6AJ7kplin+S
ppwZwORgWPzTKEKHsaPpq7Bv0YkzkaGR93BYYyaXO50MmfFlr6r2rMgK0HXD052MkGiSMoWjavkA
hYyaZJa8NImMrRzsuFIBevk25KWP6Q/UB9cUG/r4Gzxp+WGQjMy17Denz30nPhH4O/YNmjH7kM5U
K7egF1f7v5MSMxq3K/qHWFKO28AC8jY1tSBCieqU5zQY6PlNby7/ivyRaWWDS29UWKWyB5fjzqVR
9mqkmuk8i21QzB1K1/QIaSYcs72Rv2h8o6loobDT4rDbNj4b9K/shNsaStfBh3hPCtZmBERmx/lC
64DG0OiC/bUTdWvvWerJNnRzxSDaLzBZF0Y+4q4HI2WffOwswfo/xHzIGwAYJbxBxcDtgF3bS63c
mg0byQvnf5wClDQQq6uKafAhECxpbQ9TpuETz9SQ34+u/4QIFTWK5sKvtSgSJ1Dw57MK9Fbrnc7/
WpprV7mG/4gRkOrgFyeR/1aDHBeESZoEf4FQYK1MOQzrrNtI81maB1ml4Z4EJxxdUSNMQkdk8HFa
X9WX6Q9K75WF6ESiy33MwPPZyVVq55B34saR2DuSFK4hRp8/W6L4GJVgq63zCdRhDb2FliHcX8cK
z+bXYPmUfxF2IBJtM64Ln6rXJpFfOMp2K4esm275jSt2q5HlvUb4ZK7s3yOkNmpl+u3EXEYOdwEk
P5RsTeUTC2dldAgy4A+iod8SDdHcqX52X1d3Ku00W9g4AvewSibu4Wnec9+SmLiEvwwaIAH8YVEa
5RqGHOTkONnP+wfasBnrmCTOWuYLh2twoVsrKbXFhgX9Wq6mSJywqMQ/qj35Nc/P5E67xnpdttWj
0O+6eYmV6zE0EO5kTDnoBDG0fCK7C0vVYXugbCxG9nngybNcZ65f4oB7mMe4wMUuhbH9z0G1TZ9j
e5Oa3LFNT8HDRK52vvSpgW3t1S890eL8wLu+dJNg/UWAdZ6NKKR7vmHQhCYniohRAzPipaq4kNzC
tpUv7nfmWya5W4pHSpoTOaUSmpAkXbczi9kI70/6vEThwZo1mt6NVEfO1nDeUKtEkZ2ovRNBihm5
s0ponT6EiDGGFLM0jcXOxE1x2g8vwyjUEUiEBErIKYjL6MNQ6o5I6aGcgog1zkxscUn0LjE/EnxS
8zjHDR0dx8U/XL8zoA1Mq3NY4mYpZAPIxIg2mJ9A4+GxAnOUjU+1qOe9TZEwxOudehY2ie/v+iUv
xhDe40M6WaBC1ASdJOEtByeQ5bpKhOSwR16dZy6exlfqNJzXrkZrfY4D/8nQYMnck+B/xyQBdbIO
0wMi07CgzC4ixPJGOw81/DyfgIS3ea/FVmi3QHxFR632QjQcPiy5vnDjz6yXUrwJFhVTxktVkl04
1p9oL9INjZF07qJRQb5cn9iXcVxNDPGXgx1LONJdaemN3r+NsW/Os2DPiyQGhglh1lh3oUxFCefq
c5+faHqZo8k37BrMKXtG+Kg7TFe5HG1gD9rCXjDEYCBLgjvK/o/EomF5LeQS0GGShgBjP85no60Y
NDkGAdN7IxlR4BjIk7k77QXyCTyaTuaPcP1pAMnGGbkBqKd3xIN2avUQkdsBnu/ptBTm/pnd500o
/8/7qrksFb1Z2/ck0A7rNKrZIkaM04aH5ub9P/nk8vJcpndgG/nBYjwY5+Mlxgw/P7HfWWJVE0sq
XJntyQb7VfT1qyRuT/G5SqIUPUpx1vQxxEcQbsYgw/5c9mPeQt1LSac2hSewoiaoxxvdA7aUDYNB
lgRLfI3WAPmZhyMmooLdDRBeY4w4IvO5aJMtbROZf7Ox16Ayu4Hjob6zOORnB/HH3wSYdhXW9RT1
Grl5Ix4eJMDTRkXrHW+AF76eciHcP+GCAsnHrEI2H6NBMBe3STt8lcJasBXNH7pDD5VapHvy2AE5
50fPl5xAtVdybzNMncgjmLO/vzdjb2vY0lLSK8w/39DxLvCYewI6RO/Mly+SZjkhbF0GIcdHGhJX
VjtLI0ii86ydW+ZF6fafZh7zp0RoVPO5TUhmgXbcbsScAqYSk5OxOu0gb560b4BEZ5cjFldM/cJO
P1SP44v3tWjt20cKaDgZYmziQlN3wn8AjAnHxUkvbUwAOpy5kNoX3FcBt9NDmcx9DvlRA4qaBqh8
lAYcEsSCrFpOXifhPrBqMh6KBDIjjpOKkX7pmJickFgqGu3Bbj9F4lRMMrruJCWL/ACjkuODnYB/
b7aXaRkI47oSfsGZUYAatn2NnAT/apQK+lXk8fjSnMSuIDEOGFrxYptLR2doiqrz8KL2cnB5Xt4S
uMnMtl0bxLZlxaMaRATj62SF1ZvLUBEXKubY49dZwtrBmkNiUxw5Hv9xOiGNI99Eer8aBjTPTSJ3
VENFpTuOAXe1qTOsDvySgReu1BCy1XvqGM06OyrOtv3hVvdKjJoTkgMB783gVVac2o0lTaWylv7M
MSmwXefenDLZxfpKOQ1zoY6FK85/J/TScqnl778EGRod4UcNKZAeZ7d7HMr5rf1qJJMp653aEMAM
if1hO8cACIffXn7xW5GPp2uPTHo46dWpFZQeplXD/1NdwtwfBOvap/TUT4n1y8xp+mLE7/IWtczl
ZnzMPo7nygkhZUBiqycHqIicXYA2Bi5OGG15afV57gWjS3CUoWTYzc1dCDwrl9v6khMPnEaPzADt
1isW2RjN5HTZKZGcojo7bp/e89/ayd3ciWQT3nS4oK8fHXKhyomSgOsducSfaw6lJVmEu9A8uGtq
S25zvjAMNIbW7E1ld4pSnpQOjktasDfuoSz4XPhu/4i31uzqNdvkdcaI79yHCcC0mBbCNQkSHFXt
JNQyhxMNYFA4MjNGkO1HaXv6LNOIl13MQJAXEjcaMqwAIaz60KxIrQT/qkH/nswV8+l4TBm/dVWm
gtmwAe+1ggefz5Ay2mgtubHou2bL2gzov9QoMRHsyIZ+slDNi3hNJP78B4WmHbAvuVkmUEAlk8XW
Dribe2WN2yCH61cOrsHlWePXZ9AlkMtUtgxDnCMvIddNi5MRF8BrBqKOvgH5d99+/CUCOoegScSR
y+cTe1iDws1AjHgAUqF+yqO2mVRtCv+bkJf/mUya/ptTdqPCsercR01/seAu0sBuw4EAkKRGtEwi
J76ETgDpgsbqlt5U1kaWy1uaeA4SeDdwDKU1k5dje1C8qvzstJj/5C09LhCiN9XM9W2WA48hT8bZ
VvCeZ6XvvYJ/vZv0Ly0EEVoOw+7kz+NEboci/AH4PuEHcm9tN74Uy/7691km72x45qvEu4dtS7VS
qzU4mdUBBN1BH1GwYNnNqP3ea5f48ydrbXBDdeSNfdDN/j7Ax5oujuI0nk8ZSnVF/GC4OCFOdb4L
1MswU8z16sxZU9iGoGb6+xZURiOicWI+DrSt1aRdH55Qs/eB6ATqo7FFu7EeNNTzb/Pg5hIRkvm/
vGXmfdJKO0A7eLAZQYFo1HHH+IhgjOHjExAeRy5sxRMcQPeVOYBlBZIDNRRoay1dgZ0kA71b/7oH
cIQUyDmivpTA2UeyBtOWfpw4cv1vMTRMuwiZbDmmxYFhMa3juHy6WwzEHZFyReQ3X6vfab/V+rGZ
IyxXcXsJYGyKnYJGk0YSVS/CCE3XQZu4tdudxBbEubwhxAaOJytAs3NXBMiQYIZpEzPVoK2T7YAZ
Zx5nK/gsnkYXO85GK4Dg/V5q07eC76gPy+mMvyIjhFG/JgAfsJ01kBPanOLyd6sGWP7j3emFBHTT
EduK1U7jGiQf/WJ5PcuDdMMyir4Tj/Mo8Bw+L/1e2kL/cqGBbuII4Cco0Zi1Plg+v/nUrXgqogrP
Y0l7tW3ymiHceVZ2H2eidYe3Kvu8ySJRxEEWgwG0IrCtqPEHAPmWXsqat5pvuh9IGdlMiZnx6mJB
eSi0FbRd4HMIWiPopiGrIDTxy0hevspolFNLJ6wulf0VmYFKwtavudfJFqBjr3dLlfYrfL/OcYqN
LN18p8pJkzP0w392j5k+nEpmpY1/lF2P/S7+8hYH2HcTX/aq5i/946mCzuYX545bS/SjiU2c4bcj
hWM3O3dyOlWPG1U7e5GGfe1eOTM1cnxEO32eI2lpvL9FmrlpOrTyFZC5OsscT/c4oDE7DYcwwNOz
S/atnK5ZC85GFrt+/CxeuctwiTgdijgPtKgf/egtnPJeSVzCe+d8KLugIfvWmp4yUhabc4JCneNa
b+S1mGeG+RhvyjkL35CGcebIH21Cqj6hhn0PKx61xLEQwkZrWlpSO5DhQ01E69SToPDQ/ZVE1Vfk
DmPcd7j6Z9AsIlxSoXAeto+G1QkXfTCKosgDDZa+8hi1Zxh/DR+FC1YxMny0kGfbFSKOuoccjOKd
J0dz6ZQTTBIT5Kj9bBgqTlXJdnPOuxmUEuRhHa20ID9+HiiwfQ/xKIdMj5VD/tlYTacY8YrvHeI9
mTijjzZ6Y3i8ZlLWMjHh7Le7t1amzUbsAg4JeiLAgh2KukXvcvkThoFe0aSHxTVStoMaMDMGxXll
Uvc1uWnMoMnOyacLko5VWBHoRplcVR8ciC/gB8YOprq3yVq8PrW3WbxzvOs/Z78sMs5RbcHe6QhP
iAfwJx8m7PoeT7jl6Py6q2v0Qb/t8iJNiEX+hrb24PYFTcYmbVd1Dnf8pLLuV8dtGos9hV5BnMVy
gXCsf/wwq4aYshqN2w66wZw88nGX0DN+SmKdLZ9AXr8HcsZy7doUE8Aj4wDBnmzpqRQk/EknFTEg
+Ctz+3LpuhX/B98UyZa+CzeHojX3B+uz/h5gohAgJJmGfXKbnecdEtckzmvj7UfSFfeAwGoIpgaq
o+kQyz10fBdtTJDwZvhkCy/foSRCbjEjKGtR9dX1kZh+ZK02pcF2NZxCwlmIQiXvJsa21WmBoiMP
mm1kJ3s3gTaQTJgm1RH3kmnEVp/JSmAX1HHLtFKFtVxWOC51kZ+RyTvgypjafapKh0kdvjzme3oh
MxKYU59QzDXqV75ETcF/Gd3V1t7wcKLUUYFfm+Lwlw0X2QXm+wy7O9xuorwI4F9IFgDi/Ys2+y6G
UqrkrT8j16OWd/UfOjgQSVV5+d9n4yXWuKTK+dZjvDDRF/cPLFfRx7WDAWH0G1ne6aWn5VJmzR5H
2lAh6p/uuwi52BzLFrg8OUoy3j/ENW1V5UOBVSnp+/n8rQcaTLNh4JpDzJDVqXZcbc/j9hb0L5Px
9JrB9VmdsXiPL1jDXJMusojIMaxSoX8UPBo9FskJEicWfwM7nQeTnNt1uAhbW4e2T41WUwJXPodv
+lvCTg8nl/vSo+3mGKpygwqeq3TEPlV7M5Yn1vgY36Zr16x4qepmWw3q4zM9myq1b5hK+OdDY+mX
XF6ZCjSyzSh/O/yMRAZm4NKCq4Esd1vQroc4jMamxVeiAnYBlee4DM+5Rs93amFyLxe85xbmB7BI
U+mnOsK8F7+j3woME43qljHDmkVmvBITu54askmvnU+Y2BeJVGZnqyWqFmgHy/MIgkTnxPRcq2Ca
K28KTYyK6R31ruOWhFz8SvX7ihupU2yDC/rEeFeN0EwQGhiyLEAJejtGPcbrdC4x5AOBXt/jenJT
y91BWSgQ4MlCylmsd+hBu4sOvIO8AejQ9ZaHj6AnOWcndlWFNlOFmPavOL15AzlvonPtpCPh6vTb
h8w9nxQCAnnbNNUbItwqA2Q6co1bwgYOezVyo9NJzMznnGinYKzZA43R+59d2cSHbi5dgkpVQ9t8
PaCNCYGwuTLMbrPRg8Tvq1zUhOsVPFiDNOY9Ygnx6Tfe5UziEdNy2PsL9PcTq+i7clVjIc49JMIb
oKaYxWXKYG62WnRYNZ/4AQfsIgb/xs3eZO2oEKyY26+ophoToTwU3A7AAOqi2R7l8+rhz/5BJNEl
rybwSrKuFvt0xCpyHLDTVoUkfhew/fktg6axKq2hl0y+HL+ILv5jfk25EDYDhH6aSl6Ncgt2OX8V
kHH49xfTf5jRwKA27HH8ZkxRj0yfR3aRHqEpktnJTxkYHyWZ2aCqGab8M+kIsxqkju9Vi3VKGb0g
88lV08hztyWG4q77csHouimsdAWfGGR1sls/RkqMnrSHMT3R/F/OWNcMq47xonhMEHgOZ+YxmAI/
0HZBrEX4IqKNnsXkYf1nWeetowGX0pVvlNJ+00Ic9UOR24SY4H1HvsMabm5jKeE1Q+bhnXt5Gm8h
sn5kb4pacTEPcR4JikyIjwpA/AUAOpe2ytRJfi2nyIyeliezuZmljYmsaQj/ehh2gd8B+AHTOkjk
zJzfP9c4XlUbH0CUbsI3ecTlTqCYwKs0QxS3QR8k9TA5CwsnG5lEEGX8rxQjfhWmkZvsjfp9x49q
Qte7dNxQePEUU+FSjasI3zi3r+7L2CIW9+QbuviWMZqy7tZaegcy1SJhPg/QlGbRfIBvpfMqehr8
H1QoYjOmYDATGvMl5eXUGD+zTjzRzirAxL9AaiANp4GrAuKpdYTtuzhF2/t5Xg5FuIu+OGSxNoS4
JKQyiK+LwX6ofriN3lR5hOfpNeOg8p03/E5EvJb7d4qnOIKqJ9WZOf7F5KVI+ATQDTYWl2HOlAg3
/xDDjcr1DDJQ0EpPwI5x82OqdCGlST22BbkOmI9vF698uu7b2wdSYDOZENVRxe5R4iAY8iUvD7Kd
mvgfDudoaB2T5tF7xDW1cTEDWPBH2Wozn/GhyrhMg9uPsXmXmM86pUwS5eCSfUicFNxudy6eT3rg
uT5pOAVHkI1NFZQ+RBFkPDi/fhdPBjhme4Fs7rMpcBgieNP942IdqSPIzZR1TiJ512k5dijCJzkC
+xdUkETLkDxkVoDaXr9+ZlAQEcpSlzv/Z7bKgd93lgrscNpa5NnyAA5vCNKf0Iwbod1ekovtyGAk
eiSagV0vdcdgvccfgNNToONZRmPY2onHdQg3pAnGs2Mq5qruXpnr6aFf7Xo9gk0KbBljgaHWi5fU
AydI5904Vv84X2uu3ffkKcvbojBZj/Yx3RxynI3N4eCRNf1pl/ddxmQePHdvEyGO1YRhxKMEZXy2
KDRzsrta5kulD/ZOo+TM+EDyjlZLk8dvycZnCMR7LxNYf5SrH4FEH/YU8XyY6Cu+Z44Lb8cxwpCL
EOf3ER3typW0ni8dTfo/fnVZRxDuM+IVlzuPqqVkq1LvzQc6zWKUsDOuxNE4+AtDjHbGJV6J0ftV
Cn5NTD0uJkYK9QPcMrrp0G/zOnAutUlnLabcxzO+LD0Szvb7SBgE/YRbVeF2KKNAcK6/zi2+mzXK
9fqT3vsGe/YR8+eU7fDQHeAwT03MukbOoOKYlzwXfo3B32ebEDixhFNiHnBmkB1yXR9GBr1DmmGc
zsCVY7fLqp7ml3wPlbYSrt7FtSws0h5hxpDlD35naKa9zSQW7nYC+ti89nEJiMb59YdReDSPjzoD
br/k+h4sSdsg8qlbxBP3IsvEgQEM013iSlhvrTvQQPBOg26HCpSS+3oXZCOaG86bslJNPSrxRzvZ
a5SLY/lPKKYzROayULm/EyZCbfbQj1I1GXlmCmrGvHYF8K1ictcDgOyq5CRhBc/6HLOtpLKLSkZ3
rsQMGedkXtRqmG5H0Nzft8LzWzMJ0gjF7Z3X8KCLpudJwWI2NUvJWlRBd/dUr1mH1rZqQASA7JxX
gxdyn01vQJ3hDgOn7KrteKslyFlmWbOFE3IxKwjgYVqjd/83CMFdyNSJjxBZ0hJVaKQyG7h2zHfF
tVkdLBeHJHqEIMWTxIb3mmxjWSpmteB9ffA7IygdGm3SJHvlOQ64Lmxd39BOxGsK/VfpZbFv8rE1
N9w9a9NE2MYGki+5M/baJ6wJRu/Xi9FlsBl9LoPlrvb+CsQcjyJ+iCTXzhb7wbZREGOZn05lJ9CZ
3Y/a91a1MGmEMmzNFam2elSazP6CIGtib0QsUGWVpdaWCgMgsOgNWnN/rWgRvMXCmOyJImCZ6W1s
veC3z8JVaYT8J1vQV5KK8VSLR/VgnkQekPRoV6NWPF2wS5lEDW2YJyUcslAwl7Jkl7jGZUf9AYkz
y4sCvFgJhCKDbk7H39xr8Mc8oLbJ77j+qQgzFslsxsm991Awbm+s/9aq4j1jYH78EGXBaMXXgKFE
Udv2IRHUmqXnE8Ju6zBTg6w0pddwy/PNANOBTxwkKZ+yy+crChU/DfN71lBdcUQiN3eYO4L7FxSL
D8OpoB4Yx9+e6zRDG+RyVsz+qNzoexDnm0wNzfNiZNqdoAMJi+NRqdbKU81Kma7wNXIlbb5xbBAl
bKvCEnC4aWBMjXIAFeteuf2veIwaylXgv/eCRQsLhIgwK7fLXReuezvfTaUTCKjBGuTSTQ05FD7y
4ITeJIxfOdnssup+DElqjW+f1oQdPqVE67WzlUutapB0ZvCHFQs0hY/sHCd08V3LKXe5xFv3aXXM
lzln6I8VMQ8QJ2IC4LFngf7BYw1fevthKBKNrFr+7785fT/UuNTwKvSExxU25J4a9FZvvgT73Jcz
RZcZ5hYa1d101ReJtVht2n+cVoS9sQkHrOglhVwOpZ5NwcfUvhfe3UVBysd7yz+29+JyMuHIX0O/
r1uNgbgK1L0Th7/a46q8R+16EvhHA7VKNJKHIk5Yzjmzu4VszvCOxM4+hu4ieRyMl3cRMUpuB+p7
wVXwBchAPtruK+bwk3vGSSNiVT8aEATEOM6hgYQ0D/52jwGAHUvcta5UsFDm81yZzp+T/O9ewkMr
JE12HLAC5IzJTv4rCkmHBKN3d2NUhs5w2H/pJ8OXvdy4RqiM33AQtZbdTWAJ/jD80HaPbU4fXjnJ
FbSL4poavoNztRq7DJXtbNAuySZPR3nJzKp0vpAvFpBgiZOO0vEtFtbNGluVsiy/XHvUvC7QtrTL
KlCfva/4F21jhBGdSobbuX9Iro6VnbsEj5s4dwlqLPrikE8HgCN5roPLN9sf/CuU17cYFAv2RfuW
SJ9dqkBesdqKcCbV71H2TGIePHpAIHvmQTv1Zh9E6LZd61RwOH9W4sYdmRXO+ME2i0afA+GPdlNU
8TWTMXgHsaFhRwwN2BdufVhVXh2toy9S7hjU0H73j/Scox3sFhFuVMtAZ6F4iFC2CPUIpL++JGvB
uzLYnRnKXDL9lcOAbkfAWKGuwMobzYPtOcCTfg1X8NSP9dGk49I/xCykOCLQNBzenPmaDZWx5DEH
QmUQpdZ554EdZ7DWa+KnKeWYnTJwZQZOdipJa5hQh/Lz7zKuNVThZ5BbUmUPhg6fdpn6T2Ge97E8
WQcbKbb8fLnKZ0/2iP8F0hz+TrInrVFeLlSWzN3DwD4KOHzRWzXqEY0pYXC3ufUHDRsLNmtICO61
X2EU/SchvqY9c/f29iWxLLTzO1hatYcE58atC3USajnOcJ8x0P5rdP8/SSB2HQOHpylA2fw7B+7i
txZpok3Y29Dv5nP5bfmSYV3pi1Pt8z/CB4a6bCL027aKBH+aT0z7Z0QvIXTkb/CpcsTmwXKS60De
8n8+oqNB/cKDDPwx18hWIz5lXvqxk33isflQCtmBoBHA62ftAGlZ5mYI2U6wUj3a4LeO4Ja8oDld
0l3sC+/MgYsfHv1aCfCTELegu67Q+kxS8TXZ2QsVZO0a2AJnRf6gbT3toGj5waSfOz6X0FKPowdx
naMoq95PSLYbFM5jqpZSmyGUC5kPrLfkpn8ytj87U8u0kOZwIdlTJkm2eVzvlH029wq+VPK/sZwJ
PHEJxWxkmPTqwkymeV7uIcq+MeYaUK0+aqNu/Pn6ISYilErhmpg+08WcK996xhnXQZKxuSEMDYrl
GAbjJWdF1faC0/a/TlqbNFZxUtV8Nlv1VgcxT1MqJQzq39inrdbp/hyYCasiHlgKq7rdO5fyi9B9
ugx/CmIOOXwUPeeT83ouLdUjph62g/WIFWqj7xr+rQJ8uXxcjkv9NKOMEMiuHpgG9zxgBHpt4/J6
P2rBYryI5kh4yeIoqjRFAarqAJ+1dWnR+NSfzy5GRSV4G54TtoGOBqnReIYpIAcXu3DGTwi+WYUW
d3AQFIU+9mHn+La3Qa5MJj8BFTYS8Uiu0FoCQ+tA3CTYXeKum0rpeIAm1cTXqqcp9WR8K1m6QLHO
1ltTV/E+NsK2DjVHdpKntLUtpVjlCd+4Zg2HzZUspVs7/iksK6MhTw8qbaOrZeWtheYoBZ4ozj4Y
ZizmoZcEYFpjGA9CsaOf9RtvRwV+ovf2xHSrFkkiTp6xELoUCiDLLpl/F4BnOrdmfsksBE/jb0VN
7NrCB4jZX2PlH3Q5BjFgEjMgNZYSNjjVak50QhzikFDX2UYpWpYKkonmv282ArJUspoMWy1s/Y1m
CkNtO6aeAteHA85wsptfuwLTcn50GTcsoZabDUcI9PzPAtBKeaNT9Phsy4nkZwCjhbHXNWP80+Vz
BcKVHgxvzMz3MCnKSgFTgBgSMqxvq1wZb36X9erwEvTHi7O3bnFUZ31EW2NwoW87gPtFkMNST30Q
OsigBmpCz1jcPScAHwhFcFMoXykZmdXC5HWEUtpeBcQ+JLyy+0s99l6IdiTC28Gt8NRLub/jxXzW
swT+7oK3vMRzFuV2j1DpIAjQYPBnkygko8pqmss8CCafVwUITd2TYWBoGYnSVGz+Ty/+D35LKV6h
g/W252pWZH3FHT4jBnHE01eLdLmUh8d0D2o0I1O9NjYXEccCmejHPJ5HR0xVByitTPlRIo+RqJFu
G0W/98u03znFSKVAx7d1VkUSGKlo/rHmyHsSS+wuybaj2RgODN/VsGSbLryILgb5rwXDRjyGsOiC
EkUpaMKHVIyMOwhGkTcvRM5THb7RmO9b6dcnjmZhDhkZv2y6zX/xF/KDML0kxCbhFYOceIswr0nc
2xQoaK4TP2RdVaphehuhFSm7Vg7uo4/v4O0Ywi2h+iSp3zyUzOMlL8MTD7r1bAQqifSp/DLttczu
TrNbwh6hRK4Ty6sZJWH+AahkqM1HEfUhYCvUge1wK0GhE5d45iuVg4+qAbUPl8W0gf1RJIIon0oU
C0cD03PD7BhMAH/s4a5J1UWs92M5FMkUX+yt+peRW6yOouRAaO0Sqsu8j9VyZ63C1yTnJr45wyT1
vxKXTlRFTAgShrmNkgoFqBXdEbYx1DM6doPqq7bLLIxxZ+ZGC8E3yIRhBt1NlW5N+RXwkVB0Zaru
uS3rXhEgxMKhIhPCBM0MsEYC+pibDSg6HdSyKth0Iha8QIoHAxCQxQJhiuFERtvlCQ6X/Ja+W/zL
cUcfrUn2Y0ZkNB/G5f9APSiTVMF2A0KNmOR71Z6O6xTBw+JfhGAoNzrpCXtMgXZBidbYuwoFZJkV
XEtQ4MSeNPUMsoU5qwgs/NhL9PPy8/znO3144Zo8sZ4UYJoXn06Ro2IQ0zbFetHkf5dsDQCrZkZK
XPt7FL2V7OFmgUyjjQdP2w9dOLXp+vTPOYzd/8bCjct0l9YkQ5XISC9bFwQ36F9dY9mO/5oAcdH9
DBRtYo80/MXz5XzoELx1YpPGrkTOWKQibH8LWGxbrW85z/nQmkrCmh3mhxTpm4DshUKXTz7kstfR
0SHnisaOKJI+NOsJvQurXtjU6GFOIWrdhcn2z5kJd0yuvH5Lv0dSgzojvvrG/IXfg0171/cpntMh
5cvlEK0+v45yxt0/qj0Wd+Oyb0MWv6wM01RrOSyaYZUaJ+85MQZg3GEfWu2aB/+GuzE6SeaWTgmw
PQSil4XSa5V4590K6UC6sA4F19WdZaWWpisn85g50xw14ZznbnZDidIc0oyyGLNTJKO3DVWxXfTQ
ddRG0bm0oDMZz03srxwEX9cPVjq6Le7GLOpt1fAgJBgIxr0WuMtO7YZZNMa7NRBjzbDoRZzaCduv
N81tW2vgK8xQNd5uu2Qdwr/Gyteddt0JFLv8Jd7PLuwfMa/E5LCERf9ZjiZ6l6dagVebL+chtNd5
Kj1CGj1sqitfFaS8oG8HV4AEjTbgbILXhP8+537l+282w/9bjIu3nZWaUWG5aaRB9OZnN2TKuo1p
7wJXLThS8E4I/h4A3XWcHlO35zADCALqUgCbvdVOi+50TjuDzMXQbpDI2r1NMWT+4mJle294p4E0
Cq/yZqvbJASabGpPxHvbBUHN4RAPE9OmGNloCT/81dasQRuN6EJFTeMBOp+oZaQuAYSDfSOFCzaA
m8f0IjVWljzOd7pjmpdEmi4/CMJUT0niz3sY9gMmOdQe1fsTvxIAfBI9Xk/TykRk9i5NHF2Tm/Vu
/x1gNZROBC8imGE6Flzj8+m+TI4e4q0WmlF4w+vPpycnou9tBqLrPgm+lOAz+zHBuAWw8NDWyKFz
k+wUUj8Fs4+p7Xk9ZOYtCnY8UWu6vG3liKlMtmo44VK56DpeFLq7P7VHEnofb/AiV1iLmksTgRG+
wezsx9wcI8tgAOJGjLOhcOjLPSrHjChCjp93LVyu1KOhubLWy0XbjSRI6Zmmp+cUyWo2FMNPTGQt
5Y0sgwmQVE/R4L+HFLl97OYMOOxlpxRoiAYgF9vL89ZUWc3NrwgBE6NpVgX6NGBw/S6S+FThqA7i
0kK/OGXrsI3koQ2QUpC7O99ipT62QFhxbE+3XluVK8m8VHUBqnsc6Y/pg/YJmn9LInLxNIfNh7Ib
PXjyfgQYa7txvhwNZ8L0rBu/2JBXtwNyjNCJhqVjSAMKuXTdPaPreMl9x0av6ZTE9PWn16UAm7Uc
3PZ8ph9GeIv2caoP0vzG//FU6jjZFYaxH5F+wmM/5uhYjpplQXHbyGADY0m49o6+XDHcvHa34OA0
wwI65SaEOSvKYqBfKCiHBvpYUr1j9+cuEjbuvt19uhmctg/w4Jducvez+yE6dkBzzAffYASIgG5t
oxXD/Dlj/5iWRAZYxIszxb+Kk1ZOzB7L7czduu78IZ63H2g4/OmRHRzYsm9JLLhx0y8J2no3+Gez
XNUH0uJx2cZTFdf7biBe+Xhr3/DbfIFxsxo7eJNe6chjTqGk6D8RYjpaPMOHG9d1+RyCGAF0TiRl
xepGL+kPnL0ic9vbjyVN/aaPBynM566oH9vaqEFMnGFVoS+mrz80RrKquG5TcLprBkmU3CWfF6sl
3gNvJkk2wtcw7qMQgAiieLvhFKgcHwcs3EgcZvw4A6NXOnADCMIyCUlfh+G5nYYa5HTRtBPxGJMw
LSG8lbk0CCtM7CZXCiKeUQ/abT6CNhchq8k0rjddiiOG2nhXX7y+1ydhtwa7/4cJZ1ZJQytVdEZx
EvMRqMZ5tvbbP8iDzDFvlE2sxibOH/bU2JV3yZlk+PSoXFuvYlcehFaPR93NhvSyQnpQo4TMZnog
U1sdd2U2z6R8eDsrOXei9OivZlhUryUWg65c0liwX+Qg7b4Fj9GdacupP7YhdtBP5RAST5/3yFdK
iqqpyjC4X4gHhNgoMNMKQgxWapmVBRSUidSygGNeKfia8F1BvZmjZDCMjUbf52/1lZnN0xQIk6p/
2sL615OV/TCypnbgl/EDww6BhhKF+YwcbZXIroxYJCV11C/eMmY9zMG8rlla5Vx7yEA/63Nai9l5
ZIaCkOkNLIBV7UO+n0TXaPm4CGq3b3ccKjWyBboQKodWs2y4bco0padM7FMmqfxDHLxPyF9IsQwr
wl8CmVatEY3dOFtEBrO4mgfo+i0lalogH+2LpgX/zdVrjOYYm6HqwRdEZndv//mLkuKJ/Yx+WmJv
ay2M368LeMHNMI+TiJQ86K16Q8geEiE1+PcYPRWz0JEeXbKzeBRWdv1rUTCcYskBZe5xCFBBQj0J
yNydyjfa3uBjKvxnhOmOmwXAhS2mW1QZux+Wuw67Qa29doNbxcka9rawaOv8SSPFt24tqbXPL/Tg
rj9IPiJM+U6pyHOrUe0c2Iuqtfs89efqMLMNSRoRqQTT9W02gp99kKfS/Lb12wQp84SEcq9kD9B5
Z+KIxo+E0Z9h5BxJyZExheq+6Y1AKPYzWICiwlBkZvuRQNljSn1yhYTw9eZNK5vbpKAi2e5xXetO
7oHipWTamR9VzbE79N4Dnv2ex9BmBrsMeKaSp0aY5IO6nwgoKAtXHjBgtqaBCiA0bvbHFhXOIgZH
XMtX5lVBlHfXkiAjhV0kbJOvYh4TQQX19LBVMdyxorenF1y5+qKxW1/x/Ta2Iu8rSxb+CArU83o7
+ieIewXIVE4TUroL63d+tFut395QLIUwrlzXpgWSo7kAp5A5D9AJ/K1JOoOhqTYsoj5Zsh4dPMo8
qpL4eCn5/qjWIyTi+ulrjRynXKb9UPjDlFT7ANSgQYaENwsLA/vF+lJ0RsCMpVzCxpvZRaNnuw0N
Ob53s9nE660Bz/FhXggU4DU905iHTAoqHNMsNeDA0YkjjeaqOBdnggadqZIQmXIEQPTcS9XK6sGY
yK9MIVxBYDq38q7WLdQXsZzQRKnfOcLpuGZDamAcQT6mLo/xMGhaKBx7a8e/UhS/ffzrJGYZduUv
vfIGZzW3COX0JLZlXVo0yzMlNCA3h0QqRT0UzvQSQpjRqaBQNmXYP8zfrox2GxW0j7LgeGhyLN7M
IsTAB2t2nXUkwHalFOvEp44N9chKL6lUQ8ewaw448fPcCQAcieRSR4F6i74MOSRzrEoEw2/Lp4Vw
ZXMLJ/THu+YaoouUvEY9Ls5HdQwpmfKblTar7OkceA2bmn887ecIp4Zns8tADn8b1c7+WprtfyjY
5NicUJaKFV0rNr8eHlaKyIcuOZw8d9VMbjogTLujBT3HYmrGqiERygxHIWOp5Exqym2/8aMIfNx9
jU1fDUXUMLfqlRBFsyKCNm66VdziRXupM2DULO4U3wl8/NWhBqtTmAuSYZ9eGYGe5I64UUb0f3AE
PrK6rBHgVrDgmHb5fdq1zYQcj4WHqyIQFHMtkSfIEpx7qs3sj7y8wYgACd1Msr/rJVI0hsjKqiGd
yFnTLae9gBq+nBe0ZuXcovUuZltaew5LLmo8js7vQzuKL1ZEZzOHMKkWBiDKcs6eNIwoltG8cmrx
NgH8VryQArboSGnrtAkZQmz1lICcwfVshXkwQtVieUsM48nvVriHmjyYAJXR+4w84RbA7wmwMyDO
cAO3T3qOkdz5Wekqr+BcrHqpAJetdbplqxHJ1LhvE0wcJ6Rbkp5hTYJxASnayFw5oSfhyGNVoRFe
wMiKQlxMFrbpiVo9R30d8ti3lTQjCNEhmhq1Kx4aL2ykkpK6KzhtSaBwXHivkjsfoYvU4Ki9Y6sU
wiYDlqC2WbFEyNkxkXfLCAQ64VKM5+smnH0354mNqWkAVqR6ILpCKaJJ29ZvV9HmcVfHtYohC3qE
nW3+1MsBJzswFqVsMinlnz8LxqZZdP0fiCaWvI4FHt4ESJ6xcTG4FutSX6YUvpWbybJpQkqISdQj
pqGnbFEAzo4n5Ng6wU3NQl4L5m6VDv6fk7j7s20BLeVkde9WaEdHbdBaXB+zvHLXY2h8cI4x0b2s
XSprFjzFxUU80mPXGmI9qkhmEO3xrRsnLRLymDcHEI8jRDFBXyOtGT2ZuAqj2VF9t0DSpTMkovHR
cG0IU1a0rgDwjeOG3dCZT9rzyfs7oi7v0omBWg5zUVtRjWpjk+62JKagPRtSJxLCn8puR4j0FyqH
2XIky1qXqKlK/PINlU/em5+n2baC1ee4qU65f1cGW5g8ow8Vc8JHJBguBcQTnUT3L3hN0qwzaXpm
qEaxckCLMsT7JKABRl2ZoSFHSibJ6WQmOtm/a8jYxXESKQ7Btr/IMsSF9M7T4WmeA9tF0niYZ/XO
vyUZwEI4c+o9FvPdksnLZ2Skwkf6Zn53IFEGqrmtCKdUuNnm4MK0Km8VITn/ZWXq792LoS3W7ASk
/FBlZb/npAejvQAH6G61CCPmZsLMpA9tcuO7I2YxxXH1fzNEGtb3nXMeiYFvAWFV+MP+SYFh7TG1
lfX1KHpyRGOCIpJwYAOWgc6g5BLw5KMVlrM3kWVh/uo/ghds/00+4M+vcMd6cLy/7joTgEC4Wzhe
qJyr3AAJgtkZ9xkec6xuF/ypLZDeD8B1jZ31wvlqatz+xZhFbGU7kaoRZfoUa8dwXzBNg4IKmyUZ
a0UNyZyPEAoL9NBANZC8IjhViSpeg8ljwmdHAznkkbbP8/l+AF8N9nQb225Tc53oZ3L5gywbCfze
1D9BrI1Hl7ty2ZbclCEljjaER4WXTyiykjBOZJwFSZ4ZkyHPhSFQgkQpKMtp1sULjiYGb3lrhaoo
etYLVs7VB644gfgO7O4yPThWfa0ylre4mleFFkddtIcALgr62nc/Tjzs5RcUkT1JUsdRNIp/uBIA
MUJoglrNEIeN086YxjyFoLxYRQiQKRNJNvqzTZY6o7tc5gPQhGDRodwM8W71s1NS22MuO5IxZTHb
tDxIlA7ipYZyYEsSi3g3VPTWOQ2MfFX/dfxdYZXD9X6X6lBUhhARf0uFjt0H2OWjO8/K0knOtWgl
SDPAQwyxiOL8SUX/TMlYR0fFglzlNW37tthwvvxCqn1PF659W7xg8nmhaN18pLlPFt4mxbX4zeHZ
9jKiHocwS9/5+t1O8nHI7ul5QGkJcn4dzEzm9gVxhtS052OUE1Xr2nswov2ehieyXsJ+8fDdEYTT
AR06j3BX475tf56uCrLYTil6rOQL4ML5TIf9XA6WKzZ1oH934tjF4f0YcpzJ/qD0jP9O/ZXlZMJY
rzfzC+rFwEypWjIVWwI54B1Ab6aNRGhIxxLE0xpmXP5J9EL7FkW8bezDBmtddCf8wjgsI59ukuhi
2zrwSxvYGLuSV0AMKYHx3k10XpGZTm8NRHvJ+LzY+H/+r2hPzIVL7L6Ag7XaUsdmo/jFCHArlDeL
nlm7Z/466kMtFzofhDOJr7/N+FRa0Zxb4drlwIl7RYxWkibjHXCULL1MpjFeIh3AX6sANwN/2bDA
Y3vEe5bikw/8R1ZFZ5xB06jAkJtB54tPjZab1qkjZp5qsGigIY01h20Pd4ZXkGw4KFMC0O1kIOzJ
9FXIfGulzpHodM2uV2c9g78/rTYoOFzfXYeIgsuHVBU4n+/uaNLDv43cE4WZUpIb0YUj8gfIP35i
3IYRbeqage+bs3eSURe04+tV67rgd2TEgui7ndLbMNqXLLI+dxt4JYdtGRok2KQyo/TTXhMguXxW
TUw+ZX8hMADIjn7uyQUuSo8WbeOAsr4dqf/n/k7qswvWiEqYifpZ5G9ivUOkkWpUu2qx2SH7Gexx
f0GvxzWZ16K1H5D7MVDmh5DKgzTQsG9uO0djA0lMADR3GpeEZPteTKAHGAI/W15IbWTVQxNEcdWy
1yxz8nY2fB1DWnGybjXg/Cki/JIqRa7XK7Q0a/2+/EQ569NiSwLasueaogNrA2Tsyo+r+5/UbJ8Y
dSbVpWEDp6K5LNMVzjci0dvYNitoNsvc9vK6A5IdEKNDDE6OkF32PU/1GAIJYHICmecoEYclI6vY
ReEzZs1x87YlXJJni/euBmphS3n7SKsVkaiYYZJU+3yDwL7/sxIdYgP66CCKpXLK1ZUaPKx9mIIN
DWSIoHYBPwz+FtOZQmTBDy2DZNAp2kURhN6XHDGoyPApAISwDu/0U3uQtbofC3Yt4Y46+T/vhBMW
4Hqqx6dLbZMp+lu3g0bxpOotWJsDJcY29hWQg7Eub7b6BBssiuqX070EN9m85JWrVwQOXk0yMxkw
2WdPM2kmcChqF1EK6fpbW+jvJUcHqX49OXE4mAsnkKOJl3bqsXLlOdOrpSy0KA7r3qh27fQhwIjV
yYl8BuZ+00PnMXKqAG4M4JkX4Vze7AZVrReCkcLhZ8ajgzNTE+fl+sshqhjgZkjg/UHDeLe5ERKT
VFCSTiJy/9oMFhF8h52W6xC3hwtiL+TvLY+G4gum+Lkl1QJW5IPOGZF34/u7dIMldjUBCkWAPjFe
aWIPCj5ZoN/pJ4yqZ78xCqXk2tJApMOJuR/N2I94Z+jtAU1gk5NVnq5YTciL996uF0FSshC+qn2V
cmXPnjW4IbV2JrsuteQW/MwWhbKNq7yFKufpKBVrtdh483MkTF+szY5W0G/Hs4xhUIlzUVI4/fMx
I3hCvGjFrg2GWrvhB2F7NMaaG1QgrBSCCWe7j9vEngMkA402VDfgbrtjAO2+YiH8J6/HJiD2xsSW
GfysKyn+B6q8BWsKLuTbtpIBNluEVMbyo/AZH4hygRfjv0u61CQhEa3qyGrG6yru5cnsTmufN6+u
qjnJSvovooetqGrQ62RGFmJkqlgiBW0mg6SXKo+j2zDCeCI1/f62FXZc3VVOlghoUQ9XtOd/HL9b
Qty/XfpmUSICzhtS49H1sKr4LVR+ac/+gKlMDOHOymM1tnM55AqoM182vs2bSUV01ApKELLrfE3A
MbANCJtxzVqipLmG7tvZLuvubhM1ZyQsbtLbUtVfR3TNDJQ2CIA7LQdxEiRIVdGShNsSzg6SMG7g
BgQMWwin8VEOQCblOG4Matd72emJS9J4t0iQaa8ccqlvlmc3ULM2EAULpiSe7xjbcUT6IGbD70Ny
FBGqLD9AWWNXBRMIjNMGHK9OyJKDsuzGR4/DJYHOo5Cm6MDB5KESF7wakOV83pe6mI4WjPbvHqxZ
M1Bhx/bNoiNlE9uLVLTh7pVdQRp6EilDUrEzbIBfHNxTH2Enof7s6S6Ca9ba1JL/blUIZCrcvrFY
tPXf9eZUhTLnCxz2EshhAw9LGWStpAe+hApAHVGUFq9uiX0pcRs9r5uVg/UbsHxPYCNjERV9HXFu
8BTjEDAtxNxc6465uPpLaHhMxU0zCy2lk2VzIKiNQGrFenvcFclw6EErmOShZip9qDXq3c1dC17p
ncIiNlZdoHysGSo4X3nr2GBm7EsYMN7ywz7yXvEl+R8F/xARWEVOpT9KW3K6aTHua3APx14Qm/mv
tichcxivyFYhgIfZ5+uSXhoHGEREk/XY0bj3JfOT30TUAahS+QXpiRmHD1ZgzB6DgBI7/OTk9QnI
kaeB/xNkdKH9weCwD2hJGqY0FZRXcf9jZNtBDQsDjRM1VoTMCyhvBIK/8ijA+GM+rDZ2c6vHMUCi
hh3ppE5I1ofG4CnrtZKydEhLpXkWGlRJ2J+F/z0XQZV1BBbeOmtFjn3yf6ns/wXYISUTONjGAurt
AJjqiT4FAMVq3ipAs3KqiRJxdGF4kNLDD2ubQDGDdTki54dKifp2/Kem3s6UW0QFH6JXWxCaoDaF
f9telFH7NG+1tirxDJYatkkukf8C2BZRMQywo8ZkCtihhVbdqFK7idN9qi/mU8i7AGoqZiduPWve
h3tokqW3A8MmiFWmBRUd3LYM2ce/0wTrH6QMsR97B14I/rdJ9ekl2pz/e1ApF5U0CTq8aMxeMxRA
g/Y7avawlu0qJkbK2TsxB4aP4hTtvIJGG+9KostR57M4TzCdmoiJt04pWIq+Ay5Y9isjLKF9UDO/
eIUUa/mMGJS0TB/Ls7/TJkOH0on1I4HezzwTbZrEK+AlsAy8UzeyhAWIWz767uXOosbexYqAskJs
g9kVgrZRye7l+k1UmzmdFT+4P7Y4Caw5oQEEyiVFTlP+C8NTviaS7yoGme6pB0lm4UQkWYcJAXLB
bVUGfVvGggbNcrMtJR0s5hqu1PkFVF63J3V0RvonRMFt67PF/1DO37NRSCzblNKVH1GqIQz4BlV3
x/jhqKcck+yCr8EV2bjzQAT+zp3KMQsCqjYgWoVZaqnXS6NBKJ7hI4BrdsrVWLkfJwQVRZ5b0jhu
VxFnWnlJkyZc927h9TcvUspM6Zi/Co5QlrXlSFYRin6gePcDsI9ZnUUxHraIiB5LkwFJosgxHF7T
PZ7Bqs1jARN/B2TtlwOgv0C2iqca9sp7DHNyjIQYZQanlLkSruIWaDToe9JDKEVytwPCBdkEAIVj
GGpUGwcOpfapgjqrDtmLmxp+1zoxxCGuULl8uoUBciQm/1evIPt8Me3iyiolyzWZJ6duB+dUbMEe
a0XdUvcHwkOvu1gT/vAGp0DV+CYQOJMw/nEAiEgV+mfBKpnpMX4fer6F1Zg5lO5ZJ2dcPAhEimfN
1UzQo29GgEUArZR+1aBNDFq9+shBN9gEk6Ck/nbckU/kVSEIThTT0bGvjtbRcJRmaQSgpFjg2Kws
KigI5IyglvChF+uSefFc+Ls0trB/MRC0ZBBmZNatEkaBPTFrGkcPYhTmlD6OJ+M+gJonfMmwdhgJ
uo5C0UtyjoYU86u5R50HDHDe0Q0XUpVZxDmJDHIP4uwca/skZF74usMq/Aq7gqhsfmAng/yn0xKQ
hOt8gC1bAzOGmv19uSFMWoC4KevG1DP704Vw6qMXknzOzBPbVN4ZTpdRsTy/ydI2EmHwXJrqCmGn
ovbVbxSrR1Nb4Bd7GvZ3j5rIcjgG4bNPkqNoIS3dRTFv7owl5e5GxrAeWgk7xvB9wfp+ysDWc2ql
QVZ9QFQxWmgOCQTPK9OVoAmGw8dfCafp7IkIxjECYg3x8fkGxFvVeHmTVzPnYfQzZ8y0xXpQeV9D
O9dmsJPU7bFWdciHdSeprTGRwWqDx/YzbIRjbeuiCAFkzw9FUlQ+KHPm8vLMiClPzBum6vV6+rdW
dk1YAGFXYMnccPU6T6pCMlitbfHFib+BM9n/oyKjpfAcMYwvxQP3rs3W9UIVLCcb2b8LasdsVcAU
gwPkj1jP0TROBnswZnINJkjDL8fzIrgSeqZ2AlUBteLwsYA59EZQ1uhGZLTXSPIvQzS8YRaMbgKe
kwoiyYFtHsU6fqTnLj6Q3wUsMJLd/gLtR2lBbM/Rd84LvcOa8LuhBx2fXSiQCRuP8D03tGRyGV60
A6bb40FlqijteOXPDkoPf4XQcP6R41608R5tn0pNxT5t7MxhxU4an9H8jKVS1by5F7pD3Qd3Mh0I
Tzl/34l/qq4xmxdTXQ/CSZVM/QmZsvF0S//LTFb0t+vmB2Tq9QCM+HLA78nEpXx7kug7wcEo2WaP
FoArEk8Ve1Q54FqUYiXGQM09tUXQV8OUYrKw91PbkhzvgtkBNoWqLjvLi8d+yB7FjROLFQpeGMBN
B0HncJyaSonYcwmJyaW++MXCkP0SODonw0SDhM2ZnmQZdudc0+YRds96PffM7oLrGDwr04NdJI8l
OwBLrfmKDHxqmxs+x3PYoOtMHSXlCjx/do8btqCT8gmCOUhpP16uaGQk2ghfeZ6CLBdkQHNCPTsZ
y09kiGAq+N8wt4BQLGGTA9YPd5XqYPOonYlsir8JVbvteWvA5FRCRRJT9gZ/RzKc0YvW13xQHaeR
6td5uSlfMoY1jdHmG6nSepoz06AcUXH4+qRFP9qcVCA/R3tK6qvKPSxo7TeP+N3oWg7y7OZJc+e3
rWgEKtCGQYVgu0KWBywDIBzGBfe2O7g0hkF0GhQ2bxWoqSIsMJgnAxMPa3hfW9cAmXYu9fWQ3vuQ
82vJ+5Mr1+N0IKZoUqA4H60sQngxzM42M3rF+DPD9crCtFkGy3z1g0SZJFOLJgxvQD/5Zxsvt8Pk
6m3OnZgz7QTObnaexLjPObXxItSoOgp/vfyc81hCn7qlNAJWEC1DLjnlX+OLxxIodoPvOwcfASdh
nVtqandtiQNlb2kz1kC8KDgT4/cBFFMIciiy7EXcO60jMhBC1FLQ3X2wwtzWBO+uFKvD3s4xWRRB
xDrTWaJ/115OGrqHx1Jkff3v6cqCGlt3wEl+dy2KY3HDdY6Ut+qvEhvqSVmHmZnIIvsoD0H+wqoa
aXUkAWYbDuiRO5Fxkq8DUVjV8F8gO0MeiyFo7B8rz++7vm/LyQL/jynEB+Ac7qWrpF5tbnTHcukV
6vXFv2lHjXlbF51Cgf0E/R8XBl+JRHUGKsLzMfM8Tsoo8R+N9xE5kDpivM55P4J6F7ivwQrSVG+u
b5cnyObnROy0FWLEbXlPw73ljnyg5cDDBbhFqnW0R6icT9ndyJYM0ZKjLs4P6jILSEE4n/PAFjDo
U1S4Sgpf1BIGwY9aiTV5bCHOQ9JZ1PLNYkxEtkQ75z3+a8me96NU+uBs3bNI9UIZ+ihB3B1K9E4k
+c7RgDHfzVZXry6IDlgNiB5i3ICnPOLAzddLxhLtvPBmcCrs9nZouO5kpGGr5yNXW1Hn7LbOgIZc
QZbYnzVlzPwGHdA+76v1Yha22TsldcefK3IR4wkJ7g9ycHuYHSaEqbhAun81Dd5xn6qbXOd8kpAE
dcAeEOnQPwFyUdw07SQjUIA4+GJRJFoqyofzd2lneetB4OQBagylWmLKNcucjxwNyOCehSUuaUga
B7coPLlBs0ZKyj7s+ivdxHHJP8TZDwBjvEeXczgq/jNCU5Bnn835A02NbPGUk/TxSHXE4GNjsunh
T230ASVUZjpuSAid5ZFYMHMVIVkcFSBNU+2OdEi2wKPBqESFXRhg6yQ9TeJdeNz/OSImo/tsFH9K
FZMFUEKNKiR4xbBO7pI4EI+lIVn144VgPHHCf/0KfwYl19148crpwTZbDBS/OB42bDhHCvBF0mTs
G7V5mEl8fwvDpU2prIeVn8eb0lgBH/6lobFFZ9x+jkEEOWLBJJYKrRWG/IeQVsVJ2+sX5iw1VNiZ
naGgQmfn/ELg4p3tN+kzaPyLGebxDpkaPQvOBL5EOWnmltFMdIFeyMobEp2o7ZEj6lXGEUB9tcQJ
BlBwrm3+s1OdtRnvft3NPaX5W5ZVH5kFYZkXo3YdcsUybkgu8FoooUEpmsMpXPybcJJYOVQGpZF7
6qaVwKbIKhkKkrfpJ/F+d36I+kbnCqfqjNbn5BOETibnKgjejuwr6r0D+zzH7szC1a3QpRmH4EQw
ejSAsH8RPJCxx4EvUY4oPjGetUBp3zmDDIG3cI7NIlKiWLFDdUqjxQI2brIIGIkJSNVbCBAS8rg0
mVLh+CNP4gYkruX2sMgTsZeymZcWIgqnE9z1EKpcsUDaqopCxAeq23tsLV02IVWcR6HJrLh47hfE
hP0oB/mGgwXnko2CPpGV6jK+hmkxNDZ77WAo/3Wel3CcecnbcCAWObk15HBktTHp2CncXQjeao8B
Dn4x2yMZxa1fI/Qp5s0V1LPKvY+oiZ+f5CiWTSQB/eJS/5vsFW7WAN5L+VbV9Fl2xmzNm6WFxeNj
bgQeNQKvbc+fvWDSHlVuruXhOP5xd33wyxgLEwwBpvPLgitFug3ikjvzjZa3kWn+gzwdKxz/O4Ox
dEe+8hgBTgINBxF0tkutUgg6NmdoBgqMexjwFltmka4UQqi7KeMhokAOj4cR70FuDuNuuMha6Dq0
7MCg7VgJb5aBLFR5v7HXRltlW9to4Cw5+cVTogKSNL2eFcIOF2P3+xes9Fbp1ulWv9if8uOPY4Sd
G2r0nLFuD/hG+dRAHv37R6qan+4s1fFqafrDmJN5XdmwmCSWbM5CnENDGOZSkwrsXttzUBZ4LyqM
K9w/AR9/6VHLa1UNiDjDHQG6afqL/0WbyJAH72wr69y1Clp99OURPymISsNfeEqYmREifoxXy716
it2KqEgYXmrCcy2mKez9Sd4Zcroti2SU/1BpXkK7GlBC3jxdSzkEX+RJSE6oxAEjUW0+3JS3AZcW
sL6Y5h1OtS2SPGbcOa/8tFfxL2ARcv8BVOxkewTwVxKXlCRrmI3hWu82ifoMA7+I2ZZRdBkNWVj4
XFTxfkbYyaJ3MI9KYLT3Tajjpnm8WgvXGmcXGZLPMeayfZZ6hfuCv+EFzonMFe+JZ3zuqugWKDji
xZFuh447PJyhudYc0kwUatlYuvoB7FwopMKwUetWMCcu7cyqMPtJp3EtahPcNISMQcQSPDFBi5D1
PJm77cgdLzqanPIlVTn6kqwd0bBsrR2i27e8owt/FVFDUlyDIfW0fVLbYfjiox17lIsAmbsh7gn3
kntsgq9tlmDsgJMql4CQn8MoaDTD1zYOgXsGgUMDLng8dT0Ce/tHcNu1yK/P1PT3zPLf5a9H2MlT
TJfudNjcy78K3E6HqV9eylufSG7X+1lZWg8W+gag7xBPbkqA2QhgVN5ccUaB9KxaTZk+8yv4HXij
QRPR+pYGrbVWJnuuNAW+Rn/dXH8Zq2VskLBzIv4j/zNjxRw5JFihlvxTbP6+GWp5kCVYgsyhr/6B
9vqlYuuyEnnZw/a1GQ9nc7G7e0d7sfeL0dsqN8CHvmRxeTtHNjoX0GDZF+gHaV4YzpMD+p/2pxk0
XGHW/prMlhWW4aGk36Yp8LCaj1MBQfU/fyIokwCEspHnUFCENIkRVET/+l1q18PQZ2qczGNdZApH
7BY9bwjP8SKuoxrVp4kaMZYO/CEFfQ2vHCHZ7yo0w5kTFUeHjmKLvO3DexiUxCuP1ta9QD+V1SzI
LTRGMIueHOAMz4QMyMqRJ7sa4Lz3wMGQrIqgYthxoO001bQ/J8NfPHe87BSvnqHrooaellZfEEuT
QsRsBBOyOoDht69DMLfQVIiHmnuOu2/AfAnsd3cJFqTuUylx+W+PRTyPujVttgi6RtksG40rp3bJ
gYhWdL9FashtwuPrnXNWOtWqPIe2tnUYOOrACxcqGIgT3h7o8fMlaVVSYqPeuoA0FJCBXZrRvPIg
tKo/wDV1m06Ew/1jhtWk1XqxiueKmInTJfwZC7ocxQp/3dVgEckfjoH5MvHztYMvE9f7TII3exek
F7NsfaBQGoKXonUVDqDP7w9S6Q8ZvF3oyFWuf0xB1esGqMwqa8MT/d3rLC606d58pgmDQ/inzDH8
gK/wWhyVtSQmntHzRvk9CCeQRbUdaXenmGcYOjPBC+3jQXEZ3PIuCHfzrJnAWqjd4bDQdVEkL9tY
PBjU2eQoQVw5iuq5mC0A8qANLXNJegfsDOBP4T2RuAeNb+1uqWKZI2hpK852XAPmW2bU6Uyt+0GR
cP5Cbpoty60vl4jjHXDCjN5dehyIqUPPA8GOMP/qL8vvFDX5PfTK0epJ6sFFq17U//ARAxHTZtb4
AF17QfwtDV17V05vHbq2+s3upctresjdvWLQo/eAc9VUwwjWnB8oYR9aoxAOXJZ2vjDVFI27cX92
IxUmD11FBuwq7aq8SVTC9ixiYGY7T4EANawliKkpwTGDBph5fM9I8MT/XM0yQh7/48FxPhO+tVbj
cFQUlI1KALEwckRxGKMamdKBMPUlXkJm66UPdqmGEtfktxTrlAQb16EXrDtZWQ9quiazULdpKX1N
yFLBd87//FVm5XW945/jYsejdtXY9ZwhTBaFzpoPMb1wdB/bB+5b8IISLsAAjuCowTnQe6CaOflD
q/o3v3daauPbEyEnC9VoNcR+7xAl0P5SfBBLb5ElT1K7roKRFhGBMoEnsUApRucPl1mwQnvUt6+9
4jTP+efdyqg6Z7mlEolIbaAmoxhirTiHugJgrQcPG4GAgxExYyys/biXD+3O6YlQpWDUr1AhlKjR
FrFAFNXv/VIO2mLRYrP+bkTDXF0OKSHm9+3GOSa0QYfxsS/Ni5cuSUDW50cL61RDL/W0KmW7U4yB
TOUPLdnPlirCEfRw6Bb76uwaosgWETsmBKNpRqRpM/trO3uNuyl/l2g9JL2kC0z0WOShjzAAfS0g
L+MCldNE0iXA58w3r6800Sxicq2t45EGEHFn5k2Vm5weahU1FH8OB5V6pbBMLh1i1D4kJYyatbav
vNC1bVfDwDzbvlQFbQI9T1GcRzmSG9KnbiiPzLT9OqSJ3p0nPlG6igeY4vasTnLyViaIC6iN5xC2
Y0IA2MMZtQdd+naSSoiNqhZ0+CCXwJQXlPPDCHEvjx3jBxXF0PfE9GpBgU1dV5ZEpae043rx0KHg
Z6m372PA1oGHLg1ltKUY2x6UJJGNWdbwrQUYG/CXtVf3fQIFZLoOoa25WzMUmWYkjQGtlmHE3SvB
PtUXci0J4YaDmuwLY2cbPefe8BXY+g32ig7G1oML9wTr+9ANdgW7kTskEtifX2r3vZuLuHVtXDe/
LqKV8wy8RAAdcPaA9SnywitbZ0+B5u1ypXTMBp3xNtzdmfQbEbNkXfhUx8AxCmWb2dy0gP9DH4SE
vQMuGMHO8mhX6rntCZpajxcY3Hx106ZfzgqoUKyLpqVI4s+RCoLWHhaGf1DHXnt/SLjYLaYRlodw
s33WeOZKfuQFDhXDlcht0aL7DYdLe6YDStlkyXeKIw1uvMbmJ2GkNlsUwmhJWz3OQ4FqZhLVudoE
PZlMLBNoXJLXlt0+K/d3OGqDljcdX7pmC7QXlCKXq/SwUibcXfmE6Fnwwk9iNIcByZVYWSnLpCsw
EQV476uh31ryHXApszJh5xnhgd6UXesBXTpZhxUJXzhJVGlIvOWg5FmIBcEmvD+zE0ZRVEY5PkiC
yu5OGop1szHHsmXgwZl+xSAfqfM823oK/I3E3V61WP2Rx4MCdi0UV++jc7BCQMsK3545OAbzHooe
UkP3Fxxnj0cGYdOSkBCgKigKwkyoTlRYfLT+xW17WMAb5ZbnkVBsjykY/Wvoj9xW+ZFE9diUqIw7
LajkMOAniKEIMpPvqfrAYH0iYce4N7bCQ4K6qnEJR4zTEvCqja3Zu9apHhMpqbFm6IQ+3KawWN9V
onfDcTziFMAzZoxk/91z9YL4YCkEXp7Y+eepTRITJN42V9ZZ11hJ7v3ARfFM06fAK1Sd1+/huhcy
6gWlULtX/MG1Tiv9Dpa1bim/lw2XYlfDmqVcHhBiiv7go1CZv6u9RDRQE/r7ZG+SAmswrCu/4NmY
RbouMtCYuwS3HI7Pz1qQIOZG/o5I0CPLoK7GDPA1f2nM5/pV65LtKymws2ejOEkbWwEE+ypezu0s
ppCuYMePbNjg448uB43QYAuGU5f4EbO9+hgVwWZSDPPPYwRIqbdxJxJ4q2KEdQX60xqxQXyRVNXX
em3MZTf0clOIJGROuac7/FJSSBGAbRWSD14ygq+6iBEFUPHl2TjgcGnbh0JnaZ5mRLmYZ1scgEL1
agdg/AYplz6j3DPiZk4oJQuUjvNze/RRlpEqh2tt0/PGjTubsSWgC42fTZL30KynoLQDeOkI6XjD
ZPw/Ob5s1nyEaxGR9LKvuKWkn9mvvAaB+xadjGFLsRbQow0D5IgQeEOHFEBmte+KKDaRLBszAhVU
hkOmozUaXPjVumuArlTxhSP6dsorKjdA5SMHsa8HXsPZsNLRneBL9a76TcdUL3GHTrbgyaXde1N8
G1Z/ldfBKbg7adl9U/SVMim1C6mBkpyqmVmaNrA3yKnV2y2YK4//6WmV3FeyjHfoadk5nexJsb85
mDjqmG+Sdf0Oekf6L97kGsNMoLLf1uV5gp+mzQOVoYzmvUWmkITe1BpN3JkswM81sGvp9IE2pGbm
IvF7JnGUr/9vV/AJOMhsErAoLDdhvUpUdA533TPc+xD7SjKUkwbuDhOyXR17nN2QI6FeX4S2uxEz
5zG+8dQenGdUPbLIIYb6ZbTShvIZFrbTzpsm9b+x9GmMRq1bJqMXzJIzEA3t1INa/Pa3EO5KJDnK
ggRDj71DpUaOTbHIeCnRkY70+WaCpB7Z1hIfLhQc+ZsN3NcEeH/KMpAUr95JR9Ol5OrFzqri9jQt
9XvSkJFzaa3t1fz3B0WlQ2nAhFi7EQiTCMo5Do8Bpunxod/xjoh5EtpC1Ug3PYDN0iG6U1Lmf3SW
fNtutkIgmSF4k0wXxsxFk93BDgG54TO++mEPQbiamgXFn7+Bdj9dX2ArwF71c4IetwKz8ab3qyMy
cCgvrkvzyTwSrxv+z38F10oC9xz32cRDtc6oq5y2NsAvramFzT+4Wq7/+VIF+dn3Ftp7E4mRUVvl
2ECNPjUFI7zVdoIUgC8mCtvUEa+t5KhRaktQ5WMDENb4iuoRsoW/05xsvst5bRWafUg8Ny6bHt9q
Qi13js7G/6kOTsqgWWG8vJrZWn0jyCPdp+hxtKWPsK4wsSoT2C8N6rpBU89nyseRuQG/4ZhRJK3w
gv7zK/dIGoFe2TvmaTDEkk9OJCwmiEzFBLhL/BaQwO2E7/Ki7Z8/EDkB2ZlF2kwsdXid7wfZbyFK
fQfcY5HOxxOcIR50RdzF8hluFBOmn/Y4rGii4Ie7LmY14DAPvQ40AhC7r3mWhEpbk/PxH7QyhYjm
uHg5JDPEFVBOCt7z19LSaUouUPp5/9W06nabK5zU+CKRnDOyHCO/WbDDOkrEgz4OT2h99Xyifhwg
8wPiOgUrE6dsPYGzjKF0P7ys9KzHQbu03BTWeWF/1XIE1n+lHkOpubf05cxG3jNoVMYDCa9SAjZd
LlyefTgiGe4KfYQjPmX9126orduNBmldbOpszdNe5RE8Mxb+w9Wfq6hsG/rxmBJiMN2TdPAQ6pKT
2HdGjN/R8ExwuBaDcLilSQRtte6a1UdTGlesa6RXZ7obG05zPx4gRDSxjCevYkCJVnv29UXnM8QT
1aXVVHwLJSAUQ2zVzjtV36aOyUzguWHBkK+1eGadtK2iNI+fvY76jWWrX62bc+wxaQwRFVq3OIqK
rF482aNqKzkJALMTHF9OmXNg521Ff35JWM+tWJA21cjQ4nq/trJJPhLZKlrBiFLO94yqKjf3xO+D
e8d8kFX6VyiMBA5MonJ3Rk9tV12yHxtk5oLlIfkrTavaVnjZBJJKm4WCTztgoDFC3lrfh7lnC16D
EekYXW8p4WViQBTPtxLN8cUjDWOyWbvnkUWRoITmIm7zNpN0rq6an15nRqFpJtbLXMI+YWXoFb3I
SkZEJj7RhXImrtDpoJRNip7uLAMMamAx12AQ+TmP75gMA7tUXJ63I6rJtHCdsVdSsqupFzOr3HAE
QHYSrXokRBRYPTMfsUE7RSgJ20uQJepGnjB9pFnoBDPVYF6gJW926o8eiEzYmtgPvpG2OPJMhXvl
pUQnfAAQaCGZYHx+SG3nXlN8twktoXj9o9hnI1yZ5CnqEpTv6H0zQd5M9QvHHHWlTDeWJIuwkLVo
v/K2vQaPrQZ3hjAwa5iPYJlfMnOMDKtx3uxIAQpdH/EpLQKv7q6oDdh4csHWEeMa/qagAlaMqQ6F
ORDOgZ6uYRHlKWSiLWO7TVyf7mhv0BmzLPHcjI30cMG36xHv014/Jj90sKwCBL7SNmnG9E8t6XNR
DQGrWRjFtT08hFTrfTHerdB5cb3DEKs0xmHya27hcmFkTNAAM+GMVDpY8jXvPD2dFgQYQn2KfCDp
ctOvEuaQL0ollw82t5l0JelnQ7+6maLpuQMxOIOk1B1HeWwKuNFuvrTKKiG/JVzjDQ0QGnYPfvhc
5BiKKMAZi3Zj4DA30a8x+9ghcaO/Dw0MGE10XLrm1efWC0/J6W2hG02V0Ga+gJJ97li3TU6mYKo5
7Pfgp+/dRiLD5hVlG3xvUzii4cv3ZVUr03biTNHPGwjLJXAQdqv8L1ISH0DOqIXXtfSTGkXKW1i3
UaPzL9GJT6SQx8ER1wQ8fTSb273ys1CM2JfvzDGKK5Akw529jzu9K0NHWFMEh4MMMfu9GciuDBfR
/teHt51jXTtA3XQ5yZnkMAQrVcOuMz96yr6Fizsqdau1rIxlpqrcEoebT5dEoLgWAdqEEPC2mhA9
O9UKMt5xhh1gSn/E2OGMnHpVjZ8pZfgCP9xQtM6f+8X9lF7z/pv9gZ/aJPC7XO4RDwTNuWXN2LJR
KuUIWeGPXAXsso3s83dM2gAA9UpS4x/4SmnNdNXRlo8m9GrhzXx+ySSKNAiswG2PemGDkK77HS+Q
7Y+N6ZiSsTbEX2kY5WXeUD9cLJOU7abtJDzB8364QJc3EfND1KZcfkGEvBher+pV5gefkLJs7HYM
CSuIDzt4p7WUb4uR47E2uSfHvWL2MbRS/vUBV9WybRh8hk3+1Vbp++QaDMia3dEiI8LTxYtFgmTt
MytIgtaUvFHvsPNmvyH8Cmy6PhMqWXJSdcnyA93K0/I1ilgS9GvIGu4NXG0Jg4RU2J30q2ioGjSs
ddhGNwlaG668GpnCA+n89cMPVtv/+bQ0TEnX72F/Uuc6nWCb2nsrEcmokdv/5fbCxXg72nh5Xaqp
f960tNwj06Q4sax0B0L0RiT2GpH6Fkumy0lBPt1CpPACZYE3ZgCPIiatr31//04apqPWzibK78Z1
v9yaBKf5FySeiInSwo2dqtJcrpkWJ02IyZJ7xYNbwqZkpWSkrx5lMti4XrMfAfWifTmFminjPUkn
y8tX/8bBOcZBhoda54tpQ3ys1Cpr/+pZalsIvFoDikVfnLy9c8tj8EOSiI19ZYG5rfgod6BPrCiK
k91XLlXYS4+o0cp2kIUY78UTLIRuE9Er2QbcMTTy367YxjqdF6A9rYS5mbDphPIVV3JmCOd6CyP8
v9Fm0SjKu6YD+kWX0CHSIp0HzSE3RTFGqGH7jZTJT1QLC8xhhK2jcLDY13efdgYBP9DiqCuiRKU2
7SYBRS9ueIUp9x5wpAcTs4ona29Q3KG3XuFRZBUOy/Q22N5To9zCcIGgUL42tzQk9YUw8JVGU0Y+
jCY04+T4QATNWUJyIOHX1yreyt/bv09UeCnLEG1e+G6XgB4l7FjQ/76vSY6eYgYbfxOv1fsHkkaA
9m8oKwsKdAlBOAwpNnVRRxEPQrRcrfEQfEbKoH29hr7805WzIkGJ44D/E6TR66OUG3UuT8CcsWqo
xgade3xEIoXlh4i8gcTBO8Ri5LDkskzFUQeYUjwxpIJ3hRDZCTN+P8NmamQfwTAvoUohm4HjXKEG
1q0AYQY1jZiL+TYxAmAQ7bIYs3UcQnah+SPW1KYqoKql5k4OaKkiLr3nJu/G9ck81DAQfiFkrHQG
s23dU/9d0QKshZBaOeTwPEOxl2XQZE+u39tdyfmUoWs0xYKgZoEQ02RsUZLdE1jc+fVgzacx04pv
u/3S9S8MJLrRdOTHNtIsj3b4l9YHNRhvr1s03qPhaku8sO1y+/QKZjex8D1TmJ1zDBic3GvMPgNG
nQTbgIe3qpv6A6zJeh9u1+uZPxq3znyVlBZ036ZlFsCEPDBrp3jAKB8fJgl/s6Ypxa/7zh4SSJhg
WSCvuNrHAPLOtjcGZ+VU1tfOIu5xRn9j410y9PaJ3blM3T0EuGBoSjKfUJpu6MSYOzwzUEDXuKch
+6VKOJwMDig0K5DIjpMnsx3mDOSIXIB2w9gTsy1qx0Su+zLhB4UPnb94iEAqfM9JXZZjTKDKdZtm
WIjPwid0Q7Qq3C7rexsgkbBPZWehIdtKxC28YGu6o2v8o74+QNuBZ3ZQXRV/NFHje/2ztcOJNwXk
WU/4v8VIMoVJLcs827sZHcJNOYb7v0n7UNTannBnaX1M5StnQJG2N3054cePz8x7oPm36yJODn+6
fA10PgAxEbaPAVFAq7sFUxTcVi+Il22p5/kn6hEQERiGn1gM3Kpkj6m5SAJ8/djpA0scfmv9q/EK
QwtZNh9MA74vwBg7Wlp3m4qNFF+E8ZuSF8SBJXTONv/plhr0ihaHFpg3+KFJ+PCSrq65YinjXVI+
5ZXpAdBcFIgdwHeOslPr2q+/DwN8br9YabswQa9aclMgjWB4YLWYjrFONio/RJE/hfwXpXYAbZUL
+YqfnVbT+tD0M/NSBZu2WB51Ge8wOZyMsKllLsFsTrRw9li+iHiWKq71m60hmBIooW473pbGCaGj
e4p7iDCKWrShY5V4SRqEBCN8inVyUnhepQAohA4PNwuD6+nIvAV1K717vbgDk16PdI6mNzP7tdzB
+1eCDhSyHwgJetA8P7eAIhdblpVPk2CotL66MfynhQf7Rk5WEPAVo/DhiZN/1WcKAVX1S5A3XPh9
8dZdR65dCH5RBTqUC3wSwLwqDDz7qAdgHzy3NczNLaURh3eagfl6ORb0FCvlriZSMILJapIsN7rY
w+7G/jJFsJsIHFRUqymoSu6s9sZu24h12ubW2DmqyCgPpzCD+NHTrAMmPdG7Iaa3ZFHHtCnEqM4W
TkMRZFT9Dqy6/TgBxZ5i16/6gxX+tvV2j83Wq125eSsmW0ss1Q/E76Cm4oGO9xPFzMuX1NVpb/3C
4tN6y7lO2QfDnykQtaVKbhibbJf7jjukW/8M5WhrCow+0yjYEpR2O6dwNCJIKrZc3qBffpf9SFUB
0AyelDo3WsXQE9Q6hLchX5UHzvgdNRorW3FDDEIbrpQTgpWZwg/zowGl7qn4L6WZOVkV58krvkxa
giOLH5JW3dmOeQQBohAJHrDq5Cg5cZGGrMCnXrUGQqV5Q1QVwA1qbPeN/yUIg1nb2x89v4Przntk
6Ami8nwIkUd1pUruiTM86Hj6JJJdDIQgJTooFhitaS4ObIn94q8fde9Dv0DKEfgWv+GRERy5zBBq
HddiBcYDIYc6q/o6nDJ6GOZk8rK66jQOoP9r49YxM1S/5lX/c6z1fHkTzD1Q2Og2Se65Ql6JoPtu
1Uf7aoTGTDE6qd6rB+qDsULeO/SclpWqnaDpISIPRE2jZRlQB6RKjh+t4UWYMU42AR+Ll34uVvVc
m0r37b4Iwh87lE07mXiqLvNq10Id2pH8LNSPCpTHWKFX94oCHxLSdp5eP468NyyocxyAoOEIXKpx
M8ygT1yYXtxkiWNUMDSFMNUxSb7yLfG84M7qmfsEMm8J76KSb08aQhye7ID/tnLmj7zb8SLFUFMk
Uioiv/Qq85dUk6bP/BTwCXkrK6VrJZ0xi+V+YMut8q0U7dqktSzpTKPp64AuwdsvAnr3Ozq//tji
jgSlm0Ot2NdvCyvN9/wIOrt3JQZaAA+pywJdsOcMLsn36Gg+wwy5gPB0QlZaD39K9A34lcOizxlI
adenSVTpxXtnCDNrl1j48QHVufGH8IxSZpKdbHDQwY/rTu4kab4mBDtd1VGFk3W4ezVPssz8Z1zx
kvy6nuq9AsP2NjyzBF7mUViwflstjTEbmMkoUkS/WVKekgV5wjrMVulp1ZwVZRpOjuDhW1w653qc
wU55LL4BCi9NnvuVqoyP6MVxQRhfOFtqBPI0lLnnfAVw4Ew3eqcfWZTQGJ3M+K9e6YE644hJPIMu
W8ykV819wSu2DMlGZDY3QI/IAAmHGFKOo1qGWQFY4ZQlqE2yC3e4ufwRBXOw0iPVfzna0LzKGKcB
lbGZPSl7Vh0q56CN4NU/OwrRat65HiUcrDdr6Xbrgws2DfHxhOHd+BrE5vQNOLIP1QLRJ+5r+0+M
KiX6pRBnNMGNKr5pwmo+9D88cPgUvKenEBQvqz/aPolRrEQ2hrvVs8yqM4nfFMyIwTYYIJS2LxoV
OM6Y6m4lJVqPC/L26RO56C+1DRk57ek/i7lP1CeLAwmSPUpT5lbJeMysA006QS35Ov3d5pgIpzBB
iT+2vY0mvPlxxYoYbC32M5UHQt0QKQUogljaoeMx86B0irwmGrKS8u6ys5mSpBQVt8QXrjC7SXvc
Al21F26Fg2Nqao7w6EPJHas9g9VyJdwhVS/eeXaIs/rg76cmON5KeWrzIK6j81AbxNh/H1RtroBS
eNoU5L0EB6gdltSS3k+4brN4IAt6RF5azIef26kK7XZpDBbzTzpVrzRcdO0cFh6OSoh7RAXp1KC9
QgZQIZBJy2adaVBEXLM8MLyU9sBGvj7AOC5A+n9dPPEpRHAwuZLcjzVc7I84jqDaaaLEkjmHc2cl
w6q5RTwCUxGmZ4Ivak0z2LyrrbAI/qj43TumjkdEmyXjmuue+mAv3+cFLPhotLbqG7KfhhM/tTNZ
e3kOnTPkntoFv2Tk/RPj/Txi8VMpny5WQFqD6XYfRDGVu6xgxLaN57u4Kw5AF9Ie8GkBfpbxCLgp
linl0VwQFz62zKKBI1KrzrS52Am2oNGm7EuFUih0IuR04tNOPPdINIM2dW4k1fAghqh1scG6zHtu
MAcCJOzR765Gw4fR4cf1F+IQLJIPrfUTEzmwTdqFZWXllWyu8Ms8iDn07p2g6MibEukXtufofg/W
cUglNrnJwfekGIiMGcvNJ2e9uSzOQaixS3fh/Y4Kwr1vmeO9QcUvq/6XTfSzJBaRdb9NBiGKql8r
F4kBS5pB7qJ6sTL3+0HBZppryCW+GCXyLlNxi3d1rCClrvob2lwS1Kj3sBKLJFE5tGcOaBKG/339
VJxwLnEzUOagbl8AvHsyhEkQQoBlVbr7pZBDucB+VCYhkb76I9XEzwPPHKfiick4LnUOqy0UkeYU
WykmAwJ1sr2GrBsxkIR8ZOSJULL5Qhw4jaVPEA0s6OMWNZrqfSuWR6CR9sJgaCu4CYsNmTzkPKQr
e+vTnAbW4Qjo1cv7LLXFDN+Y0ZNQDjge/k08KzJCGed6ycoJL2qyC2BmKFBnPq0Nt4Ty9neZ1VcR
lyOtCMhASq4Ya9DUWWv5H5SUah8ECtD6TlY+Ecwo6EEe0rZTdV7nWC2vN30ehmSf+W8J94WyFCnh
KKpiaUZWAmIPDjx2iNF2iV9X14WoewHJNNjmbT9florZt1CY7CQPL1wH/Q5SiiHQZ5lU1rRAQJqn
EFv7/8eqrlhfzj1xca/Z6N6TCcN6YzGrFcekwQZ0v38P1wUvnVfsXDUMrGeqc8TiSqslHGD1CpaR
YSM6vQCTCzpsX/iygACeRHk4DuUK9EYrmnA0SUj27gn88SCw0clNY7B9Xovj2l0A4XxOb3QWXF1X
TnKR+LRz90LZszSunU2ogCbGnOSgjNjQ0pNzusM5V8U+KEvXAK+QHxrIeubKlq5v3TBLNtj/42N2
ECBAcqG3wg8k3mT+MKThBntXIIrxQm1BZ+MRpMJyJZYjUlG23c6+VZV6HfxlKN0nfbA+RfHB2EWk
VB1TKoYble/cq4zyT/ckEUCd9NzN4/0JnypPjrLwYlEFjXt6vnclrqs9KB9YIGg3Sr7Cho3zAkff
kd9HbEdLnB1AeCxZGUIAXyJA5KNpD8C2QQsrmwomRq4rR5HvVzr5AuFJO9MFVJ9cDicqsb/bETM/
rEm+sJfOC93V5kiPX8Rc4HOZnmVG2W1bMPsWftJ9LbLH1mcmEVrB4qRiUuS26hWrI7IuzLJMXuzC
OLfmja+oy9j8/lN3og56b7ND7LdCrBJHv6Kteu6ElHXbiX/qCZJ1TRwSRzJ4wCkcsJAMVGzvBYQI
wfk9sLSMWo0rx9mpTU0AcJ0Oa81BrzVp2yaELAIWhFosgqyJHwdOnc8HEmd15xEYfnxjLhyKQkHH
2kKD/uzQo2pngR4Lcp5/KzKi/boWPTltaLqgZc+az5ENvuhD+IAZ8a038dSzpLpG1q+J2fWH+sGZ
BE/tl7Udxn2r36hfczRC3kB8jHb3rIvHY+CIkgEittLqUgQaG3U973qvshFJXdF28xvgOLdiOgVm
hrYMnLS+eDOrqzfKmHsNdbsrQOvpIjorK7OgIslLvQjWTYdM4OQvMipN2kdUwQsQPX+2/kju/ja7
Fxz3ISQusKHALk63nFA7C8OGpA4Dzv4j42N+iIK1MkUVgPpoTXhLpukrLeGpe1aL17rZkU9D+MI/
pIvdELjLhzKN02hjb3T5PG9PI4LEL5IQmMyqqjMmLeGf6HxI1AHPyDtxLVG29beHuasimfIkK0UQ
1Fj8OoftxfMmgqbkbdVOS8ruimqle0A+SUhjWZLegrHqp0m/1rpPp9SteQ0GFSfu5ewTMOfnBud4
MQvMY6msnf3kT6/sNEXa9nPm+3T10TX0k1ggvRbq10qnEKDhr4IZY4jNiZsO5ldnH870aoqS7e7V
7KJZVwCJmFI0IwKLT4hcxLM+0DzvMYHTeypaZfUgM+5l7vsEOPLChhQTA+h+DUQg1is3Ggu2QAqe
Eo0SHM5/2Bzoei1CoLxSpiD13kWsb5JQokvO1u23EC8HJmDUwfrs00XZ+gzF7+uFfvCic6Sd/s8N
7UGCE11mTVJp52/JALteGbKkbO/DVRfKh8ET5+78xBZ+THwlVDgnGHc75WPr6iD7u1+WMhoVNKcx
CVa0e5YjBr1UPvy7pj/AOKcEiZPA7WEPld60SSlGY2NjFL0j/sFoqxglljY4H6doW6QgO2BDbewZ
qJBgkqv6P2j7in1E4oAvNWRhO6kzHte5Qq3T0oBjzq2mhzldJuThU7bj+DoHjDPmXiQxd9ENZrpW
rutX3jzN06IWNwmq2K8d+rLJOE0VXPCDlJYhpEujv47mc6AnU9nfJBg+CDdrfS0Cx+TFE3yVvw7W
c12tt3o8IZ1D9NERz4gcVW1nKE3Cgsew1dmeEKI9RJrO5bTJNWNAZ50vzJ4Yi7ghLQXVfOKDNS0y
pU46NpaO6o223Rpz59JRkXD4jgLbYw1C2pq9B20Xj6/DTJzhJJvAgj2S5hnh6gK3LSchZK3NSQCr
Y+LLtAH0hQHC2Q3J6A9SrERtyk2ZDd6wz7Fe3cCkBTcntAqtBmBbw6CaKrHM1WrQ58V1H5k5TY8q
i9Ks7bCbzvW5tpvVChkXeMtxvnzWMSBDWzQHj0se45fKKmdT7VdpIEYhQkCrfSUJ18dnvivqFsVb
B6be5myJTsMRVd19I/Ima0Z2STJ4OnGVbOi2L4oZCtNw65bgMR186Oyuc5Ml8EZ+1+84NePUSASk
q3S5B5XtcI9u8qyCsnX6A9wkkcaR1ftCT6t5MGtCwCNrx3Rl6SMU8RueyRbxtdsTA1MNoPK+G5QI
j1qfikhsFGqkDgrRPjJ0F7uSOc4ld2QbzNKjrAbNl6HwYeytEmfDOjIK8WJHIbeHkvhgryzfLPSo
m4nN6nqv/dRHfusH/WNymGHTghN2E8pANQvATO/fJ7oH1MXX57f5/8LpUTBEikjQjJ3rbq8V7JKz
UPy2iEXgaYvhsSRVQIIj+AixOLjbgRshTwWX27pE7bsxDjy3/u+d/OWZiFxEfu9TCchK5+sYLdOt
tKeJ0nC8Cf8AglymopbnVOM1fgBjQbPCcGaGfX6sw/UPBiKyClxsDHcmc7BtZdheYPAhkbvyXwo3
h/iiuQALi/Ep+e0NvflvaBvW2ef73fhC4h5/NUaSa3wXWlVYTxIYZA4Jnjn7Yy4933+3XgebsErE
bZS4zOBOQTeu+AufdaSM6gbqpDhlEffS90BKlm/9vS9W+SHg+XZboWBkJwChPgJrJMKoouwb7skZ
eetk2QU0j6VLWxvUwTOETLoUxxxirWD6kmzr4Aoye/5LUI4PfRwVnBme7YdEe0fGme3wcWGydpxN
nexEKh08Ddyt5B3ooj2tNe8wOSrt8S7RodY1oNpZj7USDhOJBQkN+W7ZTPWvrOFCE3+y6MmBbFxs
aQzZmFZPxi76cEYlrf+ZPtkOzP8P/kVVCHBsgaj5PXdDLL13o+HLH1/P1VYQEOtSNtsnHys+/68j
p0jYSUotPFqu7eP6sEXujPL4b1mqnrJzHuiF5k8GkPl6BnzCe9SZDvQv7clDixJ2TTcPu1cVfwGM
VcbS2+GLT4PP0Bxm9fXI7VUkbyU/OqIqCnEQOFEUWn04XApxp1Q+pjQKnrcmr552PB960U9d00Ay
B9lJffws0/EsxVsC87jL5jfpFspwgWbQSPxDHlhHAWpSUwdAjDSfOyuXyidGKr9zeZzsi2ZHbpFX
5LkgLZ9ProPoEZtGM/8oW/cDeL5JcqQahAg6e1xDwLYkVjPrxhzvaIXlu9VdXD7bWkQxcgB+mjZE
r9yBaivat6diGJBrqgUqYEykGFJSxyaVceDngl4+NFGDyQPUSruHG5V/pIViLHkJ2Q8+d8gSvS3I
gddAjADAwBIpI0wMgFq5dfVAVg56ACP4Yoku/H0RCqwn9gw2PQLYVj60YE/0wutKspxWWkqllY69
mI5oUjDpg+lozYSJzYaWC29kCc6UJjodnTrpzoUkl1tzlMuwbGv6uBbowSFzCe/WkDW6x7UAN/Dw
OpkmiyfUh1L3CcwiY5fc8fgnhDUVbH+eOW9scEc4R4wD5oE9avYH4i36EcEYR5+lTk+GEGP0QaUT
VBOoDGtZyZqwy4mB6bCDRfic1g800Vq+/+t6TVkqHXujjTNL+ZpMpnYoDIf0HfOQb5CYJVPZRlpO
kRowvsM5yHUCPB3bjlfKQIjaVeZG1uF1TMLeBwbFR7nLuQ9tOFBmelXbQreJEYg4L5dfYXhtZIme
xAmILzyZSAyTN1Y8/wK16h3DibRFlI01Rz1QZRQ7m/JsD/9jegYpdZbRPJL+pbMsGSmtwSrGobC2
SG88jbDDpDwtB5qdRz6M7df5QurRyRgKrsVRX97jNEHytt/R0YG7dcUkfEJUCNTGahhLyf+fQOUv
eb434uMZgop7ly3NmHVqzSVMr4EaiusSNRn0Cwld/7v2ZgdRvwT3amfW9yVlh4zPnKo1SlkWwJQ7
zteZFsFZu6OAmAfmJtFr+YybeQLrRXKiwy5a2lvz/A/IafHe6ts3NTW2dJooMzCuWFzY4LhtTj5t
CsGnjiMHe+VpgeLQPPiLTyhjaLi31bXrOUSDTABY8zbnvAlzHuL4/1OeeXlJbJkQAUnjj1eTeIFW
Zu9JkthAeYdKECW4pZX20I9/nvFY4wlHmjBg8j3FOMWIk0VIJiVwnP4KTsLGcwiPpUgATaCOb/qi
iorkkrwEQCjVsc3xIOoQ5PyOY04FfN4xfQkOnx2d1E9zzJO0/Y6RU09li59pyZemTYV65ZBLM50G
ZMWvY2JYxllGsr+Bm7NVOabKXTiANA+IBcdQXvZEv1acwcj0L3kI103y0yCIynzhudnZ7ZKV8fKj
e4hSw5ltIGrjdg+NrZWcB9Yzc924BOH4ffHRn4S8Fwbwibyx2vHfNGU3gmf9gruwnz9d6asVgRin
t3morf/71cy/2RzeUgSHDThnS7tRl0yToAupAZgRvZMjTd092Sybc5fUupBnTnqR0ybpwg/d+QGb
YZVVvcacmmRxqCCSRJMzozJw3XNyd7v+g7ks0jRkNBax6x3K48l1O+60/rnaX9cZ66FqN6ujw8GB
DvDpI8LZISQ6uNevZJ89qYDaVjGMjrF8tEugjrNNIOH+adsCcI4B5+W+e8zMwHV3XX0U64aaVsXD
ElbvHf4OC5ypUkIZ3OVjIQABKDiZFi13Nhf3zCt1V3UuPTPDFh2JcsCIhuQOCs/KKfr4RQDUOJBV
NB9EYenYqsnx0XZ6Iy/nV1Hn6uh3Az5vyda4M4V8+wZ+AcOyzXmMuHvaU6FycYnD6u6P39l/JX64
Du9H5CwvaNnyoMnUFgie4w+oT3vJlsmm6pEKQ/77I3w6y/onM/tHXqvlBRem5Ef6iC//DXaNWnXj
VCquhkuY3zxiYfZZ1AaWYoiFWsjEa9p1tfgqss5K6Hy9Y6C7Apkw8IiTbj27Mr4ZmqjOaQH+aNBo
a9c2NxOKkbi3++Xs1UR6U83m86Gl9B7jKCeH6/I23m4d70F+J83HebEdWlA7+eu8obbvMw5wdYic
3cgnAcL5sCtZvqmj67ywVZBG1bKjvMBHGdSRjTFzZ3Ef90JILIEv5tPdDu7LrlWZdz7PWQ8vibPo
X6srbTkdRH83o/j9wnMURRz0w2UiLy/fCluKboqsGbjjd9GDLv+xYMBZaY53zVjVhiKQ72xOcRRh
ZY4Il4QLl7mLxfj+2pjQ7RNoKUBFiFSxgybsZg55oCQFgUBSUQ0+ZxzGz90CidDekBoOx0tW3gId
BppvJSrGYxZ95VY/XAk0Qkex+n5vqoE9L5bzV6bNqPiaJFolFc80gjdOkRfR/7LXIBvzARBpYGMc
hOLi614W1bl75KNBy0Vcayl2U45PDRN8kiIu9biQiJPo9IVwJ5u+zfdN757ab7akwRD2OjV1v1Pf
GCs1WyuxXBzndjewYAABrBKtMEM+8FDuQd73E5+0k+pjvMx58jeVwKOezsO1wkuAZpelVycLiBav
Nd1BqqSi7Ez13KtbxzFBYdQfW3795xV2QRHQXCgO0kwyGXoSjLksMHfmldFNoPrmg+6OymF2+8dp
9085TZK2E1gHES9jAHUEOgIZVqLA3q3/2EcJw+VN8xqlnaIFSbeZW+SumLNMOPQycbFuptsropET
pZqdfu3M8cCyGdAQaHT5jjoeBZ1sdkSz0Jx47y3gR4by2berLC4Gz++qD+notKpJRJniOwJ1Hwnb
o9ColnSXMB0ZPOmHSEztGTQ/ISfrbTSvFZ7bIADrRBW924DHryZGmLtgAFait4IJpuYFyOZijxHw
erU1mv0OuQ5MpqX2y3aeRl+re9zoEE5tddYwlBxzlmWHpzPeMObxmOdqxiQ+YFypOJ5I/6MrC7zT
x+Iz2ezw5axhCv3TuC/88/ZgRTW7bEMep6L2C2qAdgDhOdtUrBzhLh38In/qOZGygTfZriDRF+4C
5tN9RCTpTdoHDYW0aszpSnyTKUnGxQUPCNy22KtAZx61IkwIRZeeYN4bRnuokV9DPSiiW+voRxgV
gFLyuYSsLK4J92SrBO3g203XgokFrD1PBVMeNSUJgXbwd4+pKGSDWyaf8TFASh15hnHQzwwgjOv/
f3cmzMucpkmWklP/u5mGCkh0FhSJ4uftp+zJiQkaDEO3ozMQAzoqxwF439T5LryZxpJN3vRPxrw8
6pFLRl1R3w/Uiij1bhCAYbz5Mj9vTaHDSnY0vT3M3FD7bFStrFsrQNvlCxKgB1ZuuXJCSq+5NOyQ
nAjEA+8mmtvNdtq5piYTRSlXimZykb9kn6V0V9na9yMTejNrhYUeujlMVlG7lXVjNiA9m9K88PiV
aFhhciTBa+AJiw9qpewTCvY+ytsPRzq76EX9grx3k1yr3nTOCTNmF0rcwnDIo2l9hkdD/aNmox1+
VU88rOG+MeHDjQJ7ZZJ0dubqGA86Qzt/Co3uhaYzPdx7MyfOMkV5FXx5hA5hH0+OAV3rccqY9eOK
tf427Tk6O90gqbLbmbT5k49n1UC93qCKkVBR9vxA+V72jvXf3lgdpCK3ulO85xmj0DZmajLLn4b1
71rIub0kgngMPfLSxvwP9uq1/aST6V+CEGS5XkBsxKk8cjhE7BxsZBSRLbCcDKPrlQMucreu1AUM
eI7yKwea4BZz5FRAds7eCU4ALT0cqrJioHUn5EfPx6Sy4ndo1NZ0Q3a8dEVO2mpCkJkJLfgE8ksq
EQRtJugJsNStYS4r7nOuXbfr58HlTrg3114ENzJk6MUfeNR90f6vFl+HYKFdVBb/TLqh08uXMXFm
DolDbt2Y53fvEyIAC1Ns33htdnNva4oqoO8CPPoVE9L0rdRCEq6w+VM/fN1860NH4cEVOublZrr6
vIrW3YDrYrnddZVM/1ceLgNcMvpt3g1vOxu8bfdxhGRDbxSxkQBLnOma48HelArOpIVKBkPLwVVC
OUAM8sONqWPmYtpPN8huznPxzTLgG+nY2kqsZpd/6S92wC3mmfnBvqCfkv90HGhRMqZ2PwOGZx66
JW/I3GIC21ju/MX1+oAa9mQZcD8a1HwOU8aw9xplh1FbqjIqF1D5FUT8yu8kKJGGVo5QMRpavGpD
HMG19oB1V/R13k6qhFrdyYIlrqqruGtXoIR+Pj7voRj64ZkfSkU1EGz687LA7vLNdkbJ9fHHBWIE
0nqUUiNSZA2Hog206DsIgeelD/o2IIOMa/hfE4lgRedLeQennreSgN+J3JqutlQEhjF4o0mCXHP0
LaxY3wV/dqCI9Ozb17ryqNhC7y9T2htp3c+/GvvewpS6L8yUTWKrob6w4eFCTupOiCKl2+EQ0XEG
ytUsp63vj+PLB9y4RTntW2fvKbRM1hi4KeqnJG6x/TDMxRkm2sg4wizq6ofjJaMEbLt3LoUuHEKa
+NugL3f2R990wkl8ib6HdC7AQXQJYhRmHmkWn5N7dRS0HMR2z/KeJ8ec+LW5v/KWsHTzRPKZiTgz
ksncBZxVV5+C9VxRGRIsx+7XDtyhy33WvZh92qGxdUNu7oPAp0fYgUoihsQiaGWECNXk2tq0dQ4q
g7qYcZqqQ2tLihOOq0tIzd2XkCoWN70TbQKh0x0oAgzdJQ5cEt8xDq2IkzPI0+4BtQvVuM9zTy/B
r218YYqcahvJ1tNHFB8IqWrLMx8JjVB0y+SXXE8iIZ59Yn/RW6EGZxV0+g48JcNqwSFPuVk/bZpv
9zRhOeEu8qOlFYx2hh6HdeiRQVGP5mcm0g68uurqfBCrgUO0z3upeMkOUuSKzuggO+FTM2N1RM6w
NR5qS0ej7hWM1C8u/oFouGpp1bcpzwVH3wypIGQ3EvJvqXHf1CpPV6ignTj0XDbpKQcj4Go3Hdjv
6bc6KTvgqhwPTZCKZMylza4QS+xOVr+LYRioaHqqYiNo7oexAFpl0wr8AD8t1dhw3zZUmfFKBzb7
uVoDtc83CBI1yqtqltReBg6JOgE7KBD5wc2CSmHh/VtFnhSqW5JW+sgjgSst3hxi+3TdxR7IXAec
6TlAQaUJNjD5EfJPflUUgsJ96zFH/ddbZD3nYgZLT2VXnew5vdoX2oKD6jv4ZPb9ITkcJsEPwTjM
Vh9k2futF1pH9vEw4bvom7owkllButGoCqgsgQD2jZl7XFb4x1m2dwhpj/FS8pSMWtzRsW7AEkom
Ne2i1JLXAi0AZ4WXZVLXCvGjSIrc47fJZ8LLqcZHTrx0aQS13wbFA0P9jJulLj+fD/mNK70p9UCI
SzHQEbGsetYFb/0hUPO8f3yjZgkTjTZhEBF5mWlhCMSjtgxh5k70VBMcdjipZHn1jdePfwWEQY0j
oQ1wWwT0sGHflIHmvlHKH8fRRss+pOGn1FGNaFAoVTyWpd1ueqLZiANZUQwP99ONB4CrPdkl3tya
qOeliCLpc3I/Ogg/g7G7/YSaKq0to1ux1P1QYRUl2ssNbLs186sYQqwQGvgkgAKQJRyy5nY5w4uR
WGMArc4dNj1HMYb7vptWW6eU+KUW9DvKJGUkklhqt+QgtpbIbeN0oTwizgZQWvdfaFB1O64GV8At
X0hrVyturX11WaydVmBsFA2lCh39L3sz4rdDzjbai9Hh3XukXjA1AdSQGndAOpTPA966YqXFUF/3
wyMZ3Lj6rAPDVUEyDRrT3BtreDST+eC1I1XkzR0JHmNVzLlSXSk+YrUkAH/eclZnH7fZhrw/8Bul
pyS/zf/LxdGPuUxug7ftY3EaBNkH8u734NGvtSuij6j2XCQIwie3haMZgzkfzOxwJkJ4sHzPlTLJ
Oo/LQvCWgS5h5AqqALc5yoXMtXwfUfVwXeoHF8+x5nlhBwuPHi+tYr4vYs7y9Iw3UEEMj6FjZNmi
+TlcUbb/KjTtWZKD+Xy5OSsmhfXK+bD44cXXPt4CLineHxu1UylpC5P2OGiAqVwqBFB3tBpPb7MY
tWrwEkYC+DXjNL34LpMU7dAFfehJfQO63le8dWTK5tyRejR6eoPxgulv5CsQUjAclwhJwpARD2BB
275xUpQ9FU1996GZJ8N2tldQQLAHiVSburoQbmSIj+6kh0RTgXhc33Se2+zmmxwSoKevkTZplwGl
iMZPA2pJlekciI18JZWMkXIWSlnaxOczbJNuo+UrvwRKvGyWH/GrEI5a7r46we5nehOmyOShuWR5
7YRrfTCR+KoaPlWU6ZuO2eHYE6jjWCWbY6ofHgIhRh8POguhXzywjP14ZrozN+Bc7EF0PRpBp2Ot
RQVObb5xCFXsQILI7/FDDBg2D0a3O2oHfjYj5UlUHwOGycqAdy+xgKyjnDmtBxeEyYNtI4+kydoH
qkBf55fSbqSsq+rLpea84X57H9i2zhggtgFtKzoXX6DHQKu/sfAqRVR0z0aBHA+8dFz2t0uTp0m5
r+9iwnytGPukKxGK1LCc5fm793Xir/Xi+L99DwKYkBOauaniQFDuDxktySttoMWD0AdsKrHKFXzX
jefoeGrwZ1o9mbBkvILyUVMTO6gEcU4lWchLeoT+MZMZYCI4bNSfx/bmvdVhGCMWmTXAfMFo/LiW
alJKllsXzugRrAReQVjlqC/mdb1DKPKJ2wpflLrDeSBGBxRQje2I9pIDEg8hr831K43v+cInKACT
XC+SXUWCkhXWw4/hI7DQtdVVv0KW5Ipr85gvp+YqFhX92y1zixl1STJiB4MJqdFh+ZkOElmSwz5E
tm93S0akxpiSNANfPqds/+wHjn08bJtAkLTV41Yauy9l5to/nChNzDJKL2NQaOVJ65Axp/k2Nz0/
K7PXEv9MrAUYnscok86JqMfGDrlpFB+x9L+c4Xf21lo7Ek1M4Mcm7sU//MVSD7mzbv7ps61m/OXp
60CRPwcEraVGi2kANqLvVajWPCSz2lMjU9NLcX6H3umVdMLEHnrQZv3ghCoJ46JvtF5ES9aTpapQ
KzqOgH+AEdNLLmpqw0uDOeNaaiOIDiFJATxQU4y4cLcm3cQQearqK43MvWYkpA3+vsn/YDj+GpkY
MfCujnVb7tvRXmOtc9S2sCd4rl4RY0K5oQ9IHW+sARhhyempd4115zL4joQYmaz5UnS8NpJnAkMj
+yb7Stv064jik96XGo7hW6hKAZPTrHxMJX4AmXe9PCfZfd2QWmNBhS3IIDKYb/BL5X6yS453vCAZ
qiijoD3WwCUXMcGD1wLICEy04lQAAi7eleaD43u2ieilegknEt6z7OK1KUy88YIEbnXHecldN4E9
RRY5/9JpdJNJrdRkoYn6S9COdcP5JjITW1KssPJCgdNsIf6HTtQAj3ttALXJpuUIoTGfyI98JrFB
8S55Yi3Cpq7RaftlaBWAaREaLR29rnuLDjgl/Lg+vY+F7VqDJyCGxdkYJiSd9bJRlegDVFFlQKf6
wZQc/Cv1q3J57U3h3dIrdLR3d24mtAEcR8VOoZqx9xhZv67DoqC0p+7TOZ4+PE7a4chxqMFgKwRr
nh8Ziic1BBcVzDkeQ5l2EMRbvyDkvnF2BEUqIckFFJPLbRx3tSq/hVkaWe+gwUEp4bCWsyNR+6xv
EyEVvaNR/HYELgJzgra3h4xcl9B9WwFldQHwVTV+F2BoMLlDPfEGnfLCWEvYEsz/q1c3dKNt0ndh
Syj2lzTi3DDTfvItx1pNjcNnsBDqXK4GW9VgvgCh5Y17iqCF1C45UMDSPrSRDKJ0LO0BQOd5nEZp
IpqiANEi5Jh0d8MBEg4GgPlKXXPEK/+wEOo6AKOmg3EgmZl5muOhEElf6wEHMat3iQwSbXe4rXk8
f6vvIW8qIzRASKj3Eqz8klmavsDpNX1QPAUg2xmMNC4TZrTxeVCrw6gU95gFW2e/85LU613oyayw
7smIUZUJcEbzDoSmIBBUfgY+GFE2v9wRZDP2PFZGA40hb4PIFozvOkGPjPV9tPePgCmierhnweT5
YhW4shpFFvwG6OxuQb9EY2bYBlmYgfp5wo+zyvOBguG+lERP/l6U4LNyJ+Uv4tl2ldvXohXjiWOh
S7SsSDUr/qY7o0GmNp2D4f1UBgMKj4ZTGqO7VFZ5S8BtPyT7NL6/b3faQpizCPlqORv2S3hPho/j
1DorOq0CK65YTNI8uJmEi5/g9dgYZlOy3WVhy9tsNlyiPZ1wqkL63lsxgpsxS50ebGwj4Ep1OBg7
S3aQWSUPZEkVwn0Okip8Ea+W5CtMllwOD0zYTylcl7zpeO/ddzcwyuIidDny9voprzaIyh1whMWQ
WuWS1xsNwAOxSzXZdUyeicV4M1BQ8OHdP8WB8RtYfkmOctqyeP1WWAZY8gm14QohBWivzUXXRK5U
tGAO7kWMirMIR9y4r0ItELtQIV1W0yYgmvE+nGoD09zPdZqXaO/PoudewMlP+zvsTrg0YLbgDdo9
MbzusvqqmyNKwrcWratZc60u0dr3pEkDFEkOwLOem/NLF3+eCv21ilqDbbWW9ExaF5cgOum2Y0n3
O+gubBduLTFOLCKgk3/kec5+Ttn9TvygsGuBy9LhZsmGctBWdTCJh1Lg4EDFGokXPu0ehTSx50To
WBzP6+E0uwsj6+5MedCsH3tJRVf9o2GpOE55Dd2xBsHnt0j/KizP4WsdfBAUlJsLJFZF+tGaVfxn
2CoSLSJblP/Z9H9RX6EnWLRA7g3aqOte5iupn6TjejwHNlit4pHAMGr3EDHcnYxVNemrsQyFa+TM
Kt1LFKAlhKtH2UYMzTysF65W8xnzGRXISCqWKeFSp1a4wHaaNF3eQGJYXrbY4+W6Gzzj830IT+7Y
ET2v8HAP027kI598LhFOki4eaUBc4h6K7kzPmdUp6C9Ch9HvbY0e5A3HniKTQpFv1qax+KM0L2N1
ICKAEJ2Rp4azsQqf6Qh4p8rC9IHoE4tCZyQH9UTcyQPO3vFjAq+eAY0ByfRhJ1E2Xx6olk4eFLQR
3JZWvZR/FKvl/5srdR4s6bbFvpgzv4amBoZlGZ5sF7Ch8L7cSEazEJSN6EX4cvFDLURlLlzXTVSS
Zz99bXP888xE63ZXKQr0E0sWwwODapKS+jZj11IMsYJ6JKYQdLHuAlT5HFfGUXXxQyua9fSPdnzu
98npKUvn8wZum1fMAo+rEOwCZbJewEi3IsEdKSwRWoGcM1VT2rVwnbEhiJmXMRi3t9jHEY3bPuXE
6xFCnb9r5s6n1RXZKW15ZdrqVt8opm8pKab8uTbIISRWjImZ/bRGA+xT00/G+pVPRG7P/51Au24a
NCxypgoidxvZ5e7t1GQ5I+VoViULfUrvG0tce5w5urnfjUezgNAF+NouIMXveiRVTXww+kr7gjIV
t9ELboUpn2jUl+DnR7sb4QAYCpB22cj5lne8nnf5sQT7n0jb0CAK5F1xZNGSXJRwn8bTYM08lEvo
zkENM0swrrgtyRMw8W01kkBdliAXU3kHRhFlGeql+XASrW/O1WnI50lQC/PeqAzFvvv8qlBhXwwf
fJ/Eu2ODx0uSgKHPNehDvbivjcJt7cU2WYSrGIniSoLEy1HRmx5p0fegikEDmiDklZsiBmhBeB9M
anXaDm+mB7p7kXE1SCN1jtYB01/9jzskF3vVpvlSzJWgA4lb/UbXn/aiBrbYncDC7cwp5JKgsfIG
3E+41pAnxyf0qZ+mmo20H60xO5zxzWHFIM0D6UFNcHtQ/mdsIwFj4CYFngBOrCntfBFyJOicdiLb
fEiqc+qWjXhC9E5xauRbFR836CvfBrU2su9SWVQdxeooEMypczM9OgxE2fU3FSmuUH58yHrnKfi5
fqXkvHw7PqAp3aMxFnmIGFQ44+h4nHa13Ayp+i2KtEtDVw2nJOm1Jiuqz+01fB3CELt54/ehsSMG
ZgQH8fApKNhxrMx3aTTrRLV8yDphPOgzJgtPMtEBkx7a6iiM1SBzocaLgVkJl/avUSsH+PznIEaF
P18gZa/max8CinlC5eiP9xubWyibZWx7Zt3sMJYHgyqt8tkScWe7G8qsSnNMArg55uLbP1c2NHRj
qXMZqhm0jcuRY+9mdssPhjg0SgP8eaWwJnynvzbkeNRnZxNqFbfmDMwvgzCxEJpEqmIw9iNoSVV+
hIzwr8sSIis4BPAxOBONMjgIGfteoiLtRNyZCTP0R9boMLm0WqruiXoRIYsUJOjK00GnjSPtY1mu
9le0RXpuvlWWW1EFRH7FcKX4Ud6kTCoWw9/yENTcRwtvQX9Tax39d6k90tzgUZ7qt0b/QNw0MZo/
q6qykki3Jv73yx3l1+EQCVHlZJ7B1VpxX2aS4jy8tZdJDnvJggjBIb383fUGipG55BLU9NDV5cbI
imrosBt9Tw4QYF/GOeIffvufdaJUOs11HhhWplqtg6yARiRe3dofCYXmGUO/2OHDsvZ4M4caMO2/
u6UFcmYke+ikZhTLtCl7eY714/vkItzeoT791CGH11huXrL+5CvnaVrjqXtLBbRM5gripo3NnTLL
DyFNRARQ5oawAs7TggCVBCOw37ba2kaDPBGXLn5JCDjw5K73X/8L1lwEyAFl77TEoFrIcfEa5aox
jgtVKZld1jDEhugZzEniq5NJ9IsgC6DLU5UDTH1w44flYWIpd5JaFxHLwzi0vdTjGzkmJA8DA621
98kN/Yac3Mx0lUHxRnVdjx0dWCSBTBrCc2idWF0QDEuvqGc34yfmcxTUzBWoJFlfl1ACvBQJeLVV
UXtY7kG9GnvOzZyh6ZkpcHHoaFhkojflkwdqfzpHLx3V9KqxmWd8jeEcPknvddYaFz/r99r2YzoP
yqruLEa3pCRYFZQdWxkzqe78h5UsI762mpKmtRckV5Y8ujtXszAOgYpofeIUuWk9vkVan/iS8Vqc
7f5msYLvIqndNv5XLBmoyP5Lh6JeGNGmEnP+lAIf8z/ieq8jTbPxbUodVV2zirEjf/oAXJCG0rG7
QAEUitGcIXkLjmKZPJDKEkPzUr7rVWpYy3VShgOLVz+CDWF9YIH8Wtq4xya5H63e0kkwQxdWaWGT
Z78NmCAGN5lmAhGFV82Qlx33ZL0TK7416ZDgY3zKZ+aAev9GIoLkEQPDExhjr3DlpFM1WUsXWIXv
kWhZtssrEWcMskzr0a6aCp9f8ujRxQXojJcDzYl9UzaZP3RrRVy67dX/oGOO1lwy7maQR+lq2pXU
jKD+GbvbYQoFDFWK0pAzNgqJbfRcXbqXLZbGMISTbFtvjrqp6zdQ3J5nSUps81tC0cCGuaLpiojb
a91mt6vrfdTRo/zLCyqbD8jKJYv40lvZYXFZ6bEuhj/sW+YJjH+kCeazGUNnJrmp1roIuIcEM7VD
QodT9cztGR1AAAV2skHhV5Jc/lMx48Oxl3lLLJ7lpWpUlog4tdkJgyMdobhwwBg33XmSPM1hFnP4
Jbi7Dsf7XtGv7gLcbTzSz2r981RKKQiylkhZ+0RhH4EuuhxzEmuiX3wUg/k7S353XFSF4tUV3GkL
gn6UOlsc+dWjBV/dFafLNYZTTJIlkn9lmXrD7ZX5EKU7gYNoo/Umc2ubFO0CvKCVG9LTwtzJPDTb
2CBBWgqZJtrnAEu+ee+gOIzY9nx+BY4fQpielypdUOVHNpqnIBzTdE20BzKnJMxWwfd6bx3uSFDa
dKbLHswVAtnpHP4FcMrYVOx/0QdOeo8DTqczok1JA5WxKX33Dg1ing0Xl3o3dJyxFU/W32/Qt4RF
pRYSyyGJVEUVz0xTX3sYSo5gzi6+rECjqbCazuQ4s0nbdZGJr3ZxB+yXl9gt8bHxDnnhkSdmixHt
KOjak887p8/j5DrkgjYGsZylr8OVd/sBKYG9SF+kg9GtW57+vUibarTZ/ZYq3FlDxNZ8uDXUd2ST
kAiuEi5E+/jF58kh1K0T8DMc3ccpJ3L8/GgGKgCcNYD90J0ZY9G9sp0yvC31dcY/WKECcv+NIdcw
RWqDXLmc8Hn/9fBSLZb9KoDg1ygqA+ws5RuP5Z1MNXKFcW7PKnlUPunlIzG5Or77E7ANFtDpqlPm
e+Oul91kdxjwvAzGe4D47QlaHpj4K5ywLc0Vt2Rk2k1Wvj2+rewEFnmr8aCayT/VWrXa81yOESZh
J8Qah6cMe8oSz5LUxMkv26AKfVrriKzMGFi74+KMAsqS8+isS2ZXD1SGONFudaCkqQTr0quhZjRQ
4WOxGH9I/zCEoWtS2L4Zj04hgnk2Cyu7oeT89L6GhlvadbIMdbZKzabV9NJT/NKZ15KrAB5x+SxB
dZsLZ925V03ngk9l8TiZRmt5ptU01gmUpILVcYby4kitzUrXMQH/Wp+QFKtvB0lp5kL0aMJetvq9
AoOMGHO7xSPnOfvkwC4sXJs7A+fxTv2D273NHTBFqCJKDaKnNgH+XocJZkA0d1qvcY6EYu80XEH4
q1/qvZTHWdesH+KJn49O4fg8c8Ag20qsmc0YrBNLpKfy2BjktL/ZFevNf1ZfqC+PfDOZruoi3X7p
cCe2dHx3fMPW+fLIWT1Gx9jYQt8RuAFf7GtLZXzWXX84DMAGzOhGRioaWoz+qyzWk7n+AtTv+Ka9
4b4wtwq6dHyEHR2nz66+QxJY/swco3zISqfsIppQxZx53rkai4nlLNnTq8VD9KCND6KEfQw91hhW
BO4nxw7iSg1gkti7XUSQJoZ1RCiNCbkMh5ikfuPsvuVrJ9aSo77BAmMJCCUtVc671Hg2jdPftOxK
MkYXMpO9AOMrgqi4EfIi0mvHhX7/kGI5eJnVbr1icQ2qUi62rEOP0boWsk+ALKEJTgdGqiaRmxxs
yFXT8t8GCpu8Z+KgyaRk7mTKOzkxWEWrH1iVj+ewh3954fNbEGBXeLH6C/kuW/0Fow3y0XAzcfaf
Q482tVK8fqrClcRZo8Z3NDW8nM2YY/Ng8qW0oGyFc4kIoCrCpBDXPBb0XGPR1KNODI5uWLRkz8mW
Dq7f3fUukbgob9pwr5HVQgFh27h8DSa2LXtVhSMgOiurUS9enP3PtDO+dloTW+V0DzLmgfQwlrtr
lvLelPhmPifhJHicTfWQbZljNMy8xAyJIuoLgKXFwOLlUVXaJs9uPURGbxnIEqQz+BjY/rRNHrPM
K3/1eIP2af+n84nMVaZldLhyAT4spzrC/oYuWeOzid9rfDsIdxh9H/T5cJVBTqtmtKMPI/eoYz27
YO8K2klRVyvRu/WJsgGE/bfVvvzEXmRZdfgBWRqQDZbYl7Eyf5stJ9DfBzZbkCHeZGyCVirqq/x1
+CXgXUWrkoJzhKl6ojnOHr7HlWGhlVVG7pL9Jlgggj29yA4YTKyM/JWLsSR0Wn9qX47a3VzRNdNL
7qd5z3npL29Y/VnGlE0AQqzkt8fVwHXfKNB9MrH5rV/astzYbURspOkX9NRmSWC0Vlxis9ehJkDi
zIJRpJ7iKHoTKx9RBZ3zdFW9Fu/I0UJ5yjeLopvamm/0RPLVhwy9ZyegK62d/D4UzLEPu/FfhWzx
VC87O2ndrfUZTYzJXeJR1SdX3rXYV+wBH/R4Vr73sb3gfk7rhheldzhBX5ld9TRWjRSMQ7h1vEZ0
7lYEOD8L3zuM/+hYO60FuAiiwldZRI+76duchmFnJRsCcmUgzZ9ctYQ/pDIXousdy6FqclEFsPg9
pM+iz8A+YunSD7uSU9pZL5HwNsVNhpjUBWVIk0WbqgpuyJ75Oe9fSkqiFtNe0Smo2izsifxPlYX7
lcWQNGZwQnNOEct75F6SJ6/1U5ZyDg3fNIs45wh0ArnMpiHW6oAnmJXtlsQSNCdGdkAW7+EMkF++
GsQrERFYKck1QthG+4KYfx1gep7/S1CpOJYmlQzZ6D3DnScpSWh9GAMGD4RhrooI69ReVaCdhzTt
ijJIb2ynINiDgzJFaEC/vyPcmprX5keLPCgwlfc7b/+P5vpqzJV0nUk9iFzNRR4s1N6pS6mk8eMl
Di9sia4kOTIzQc2gEPE0IOEjkDF0RxZjncMZKk+z0rceDOnmtxsNNes71NGTjQcN1QzIIWvZ9kKn
1uZa8x1EZBfUdhCv8BfBblO7OUXeThdrKZNiOGuzd42gZ3GbPv5yQTgrhuiZncsDHwcfqPHTkwVN
Jf0H1EUf4VLx/PT3xWUns+XAavYljgejPm7WRPl9PbNLmcGNPQTQl0q5WiKcqZcGWQ1OZKZUbd3j
aRCBW4FvIdoITXbgQI/SlCA72yDxaOpViASUSbYc+9WTn00DppHqqkZ38bxAXWC3hVM+MlaMuM2s
30IvsadeJGu/IE+aAT8LQmsTRKjthmFMZTJvd/juJ0XS/xQoOIFGQD+MWZH2+8GdrdCrrpRGWy5l
Hl/jIZ6/Uw1edMoLWxiNBQv0RpQiztzNwtAY64s9ZQuqx4gH9geuSxOZ4sufqY+PVITea91M4l1F
SAw/HPPB2BRBAEM3dwSTK9ZYyMR13Vi+8dbdpWSXnwtNOegOXWrGxgJuDC3qyQ09RNGl5ah1Eppi
hFIC7cnyuwjkzEDsZAJju7ST688vvqZ9z8XTxAVGOvw5+ef1KBghbuh3qjUyGgZMSI+WFtGEC75P
tLJQXz5WQibFp3gsNwCdY4Kqay6w6BQY9T/uHOSeoxucokyCjTAb7RSOIIvmZ0BHRddevvObTg2z
J1LMezaQwWiqAZ6ZqgT94/uk+4VdWjIWXJfWA/yxEvccZAFESyPqlwD07H7LdbLje0jkWz9TRWYE
3xst4tiRzGgMegKmLr12d/8gYqlOcNrBJ2L0lrrI3Dk5wAGk16kEuWFrwe34Nn82915yYLCRyz4U
cBIaf1ScA3KgJxQt+FE/WctsC/32hBWnFyCIAv4ekTrxryDizBPb2Xfb6se+u0Wr749M0YSvdTa4
XuN4eNJVr0cK5zxX/ckZRFQPSSBOWwOvT1TwxLdejNMj6MCTzQsMdMk6iGrz/s+vSmeMF3EjvFDC
4IOF5sU26LE91B276lkJQmoaW2mqiib3q+FO6KYqVP7VWvAvf+wBEYmy+D/Ml8fAunCiovBCbdc8
QSLb8NALuaeBTiD2u1GwuetjZ29yRWjZTZuK72WzhdI0dFvCo+NjzzxpV5ZjKSUTRURbWOXSe82B
FkRriExbJ1uScwpaT0o/TFGnececeVjzeL98c7t6RAl41NxKWuKSSBrNSmUEtEgh4EW05xu6n81V
vMVvgh0V68i1+YVrmv/nVxkWMpohMf1sldmkJm7U9ErtCcWQQp377J2VCrhp9jufNhPufyEGSben
Dx7PA3vT9/KTb8bqDnfduspcY8d/ejNQvzOIOKj/tzYt3N2oaTqJZ2/8WjIfk6/F1FECT4lO8xPB
v9NzYEagRQMY2QxUsuV28B3EP3PPV+uCl/GC0SbyF/MUI1GLTPBgR/fsggkMG9u4t8IJ9IiUGnFL
1gMbNjQiiEd0VSmd6/o1HBdWih47xOfTrCk0Uh6WiYJXS6fXG/ejt98ePd6ObFuGV/6UxzZv7Ydh
qs/pmEqMCMaYw5bgShK//9Zz1dp1yg8L77MeON2bZsD/oAuzGcZc/SuftEYdObqdO+eb5T3pwo+1
MfUF7k9Sg60L34BDtmPDzT+ezQk5aeNCP4kqqa793NWASj8+rHbyOfZQ3RMdp9u9t2XG5ySZ3pGw
UXYjedEaM7Eti9IW6hDcnvWfdFwpuJ1Q+IQ3zCWfv9vLcmuqcqpv1BLvhyn1l6jHhdyJHKzM3/lo
yIuggbstZPk6HY6eFeEEL6dUUq/j6dZhrSqvmxHPPc/7OD+rPvNay1qSBteW2iH+cfNRP7/Q2KhF
iCHOHfbRmun5jX6wYhOkPl9YtHxB63zKmWNQ1T5unNRwMjzme+cZjf5dGFAk+r5IFtSiKG6tCsUY
alF7H60O855DZprHtBJMyiViUztgNFz7vsTctpGG83UVsbc08z6R3PIHs4Uz7LlW0dh+p3Vfrc7E
3LRllAhqa27dRE1s9tAClcCfLrwBkWMuCkbiW43TB49EtYwHHhTM6Q6kHTG0IMDmIu29/w2wTVx4
j0CLkx/QJa6hgbQZDdgMLrKMxZzkFy/UKfL7P03ugi3JD0WOxd8C84RhPmML1mmM8ctfbXLqJ6so
Z9XoMXh5x5YmRalS1ZmZLw5BRyb6XzVmQDwWMTZKFDP7g1k7AcXl6jQsa2QZuCWhI56A+f7LNKTW
9wExVTZX2JpR22JYnPC6uh4l45UtKD/xf9m++HQdCT7fPyIxlClBPTMDilThLyYuCnfJD8xLjpN8
GXDbrHDHgFr95sBDmQI+8uCXeBGwI5DiHtN1e+peVsuaz1o7fBdkn2VF6kdSB4a0hx5B2KzZBLRN
j7/HQUm8hWfIc0/Vp6YRMRjgvp5GRvLFEmm/CEzjk3bC4KIDVl4gZfITsaSUxi90oRko54JR9RnF
3P74ZKGKagja7eR3S77G+OknCAj4QZtL/rZcQ6B6iV7rd6ne3b0eZxlb9lqsmagvcVbhozfiX/Mq
zbOYEgOFjEShfk71zliaLsxbV2PQ4L+uf4LlSnRdRKlUldq9FFXRBCXTzybCzcdanb9j0YNQVvxA
k3nqCFDg5d2QWPLn7F6Ba3zbRoOOoH6f1j7BQbZQbxQ/c5V0rRr0zGH4INWQ6ZqHcDDsEv8dTZfR
1Auka7oXmMbX2qbTNEeZP76qDoAJAAHwiAL8tAxv/aUUgil30uNSYJLHDgnuw+9/+c/r87c7aNE2
37e+PL6O/i0kG5E+qDqpQ3Npm5vUSyYuoOsI2XZtjONsrhs9csThDxfXJkiqQ5pK6hD3rY6TmJie
OdfT5qFTxVypHTdpNO5XG8ynSMkIYd9aF90j7gszpyMSd4HjipzFZgEvpo1VSTVPfodHnz4uHU31
s+AqXipBYInU0v7Ki91pDSND3PEX3g1oE2HBBs0t6oR9HLQXjY1vR+ZIVNSypgtTPS+PmbeHVdhh
o4HIi1EZhWi03FehdfWwSpHcekWa2GqvOs+nG+y35DDMLnENCFF7aPzNb89WSaT34AcfoaUCGysw
ewU8b4KlC48hgkdkGgOUUUg9ZB+OoJGYemyFHs4jWjIOYSwj2DYH342jaja+RS5cXTKN0CMlSFg/
NNw5M2751Aqc2Qkmb0b+gG0HfBJ0AlbV7Fgxm2E2weiJ7MkDT1ibJaLXFg76Q3bAYMUNVVbs/vIe
hP063pkm2l1uPPFng+odowleiDAZwgAingVipK0TiIf5ppk/6jXN5oy3FEEyIE2kjLyo+3IaqCUf
WkeNre4gNST2DwUI3xXZKDHyXqvP88vpeJwpXqAq15mqOlFSc6RHaoH3ZCk/Xdm4H0WFlO1W+tHk
sFRKYqZwm0/yIT6qRPKEH0fdHegflRr6IQ3Gt0/zAnWt1JPVlIEHCUlHlkdlBIGZT6PIiOu6wWKx
W4rEVuloa7yc4fQ8Y8xvdJ1r7Z3kSSVq4e62gftKVhqv7U5LDaGdsPJYZvnWRSHj49TJo0xxbTKb
5tRPU7ePXKwWOktl+I/ZC+Ow19aQ/57tV9npYA+vPo0XgDnHg4JMBiPvseIlAiaZgA/V4qtol8Ju
nqAUL4mZpCiMFz08YUGQu9pN8YL9RbecwGaMH45iey0b+oz7YZtS1qPj6bpFosEEm4vtWbObxzpC
5KJVgbIcdBktnqfZ4dsfNDtaS2ct82O+agKcTiqQNsFJS7XZ+pRQyKgV2SZ7q7BLxltUMOdM2O1p
dA9LqAOb6zdRUOSEiaAIN1e3zyPPJeKpVDfDci412yhx2RMtzGGLXZwYROvPcNZyI67vbeVc6kkh
YWl0mbFcbSKxaZUHRtzhhLNZ8a15eGU2l4k6GyDxoNHuyKbMCuBfoTSNcgcNed8ugeypKMbdWm3Q
Exlyrbi0ItgbYYTSkiNdnJq5I+PrYzye2cMs3JsvWlB58X1TAD9U/qD6J4zZdG3DVCvEDt1mzCiP
bwfBscM9j/5ZYjd04pIYimcK29TUJS+Q+Y3a2H0A34Tz+LO1xQ6Dup8/vpQvNg7HNR1eLrgyPoJp
H2aLViX8d7gNyOnzXsG1Lnx+vubObD1NwqPith09WkFbjjdpENz80b7qL7ao7RXjdhv6KGx5Rent
kpliu8c+7mlHDi1q+7BZ9ENL6ZCeetD+hbzCTLhwzYQfFAgAoUPwJxtJUMOcKY9bNORfxDd8LyCA
jUpZvYSQfombQG7eQvF6fpsMELgv+U6Eoas01aJWotwQwmyWrMQ7E2FMDEOwvF6eTBV5nM4rE6yG
4RapSh7WX8dt3Ul+2HFssqLtHz9sQf0DhiR0dtKsCZsW+jLkY2tiUpvWoDtLz4kcG5TPZATn360p
Ldi73ZK8uKQN0EtaSCQk27RRGJrlQftmtfMY3WB1X3QFWq6luZns3vuIasj08PIg0Y3f0zQmdSvf
p3nLt4AXKsPHlNdLJeA95dPy10qAX5Q9NjhU83kG5EvFcyfLLA8rcWOcfFHO4kOgK4SVSdncpghs
pwvNm+z4is1jbhhPAZO5FOX6osAmcDyxfmGXGGbDgOkXCBZsnmzivHfN3+0hQguCdb0WN+fRubvD
s1Y6yDny2WKYAGJJ3qzK078ve1j9tNlueUTGiX6VWd4MTVUrUZpoCawUm9fQmyG7ZBQ1hE+Ww07s
z8yiQeIUbyZML7l7iRYmgRU2reGcpeCpy0D7P4bnPkeDmUhHWRTaRwrGepr4rnofaaQblnzKR11Z
oorU6ijppHYUYUUHo6dmykbKNULA0dPlIJ5IVILd0q0gejYapIe5K82KjjXd5XyoQI3Fnx76xPI8
/2laJ1JUcQxR+8AaM8nK1B7YHSvhpVN3qyi1A67tdS0mJfd/2R16YpHbbhLn/txyu2crI9IcZ+Yr
Xs4asBSMvc0ntOeYC119yE3tFUiRwksZy1Ag3E/ejs20e6UsLqfCh2HGaBQHLnm3DFKM7vdOJo7s
MepA/MuQ+zkhW1lLeqnptvsHdjPUOfvzpWWepCgYg5ozSCRXQhMhEKhbBmY2I5dp1LzNn8tXbI4K
FZldPKCtCPaoGFCfy6wu5UrzqR16SE96/XHFyCdw34z2Mu+SZqf2XyMzPK658AclFlSaOeltQwaf
+/shg8vwUy3u2BDyDxE1Z4pjBA8xdoSTnbsxHVA2NGchttCIt/RGRRlc+1FEsWHTn9tKezEAVjoI
iTgswsRxLPQdqDk2IKFo+GjjDIoWv1752UJ/bApJ73+H3serbfqCfG/e2z4FOST7Kz9o2lwEWGIL
3JFhnBDJvWwv6g0Wqa3+SLr0lc96qKWtOn6qh6b8jjCsabq6XZqrLunhqHTI2mwwXkCKqyZrNpSb
de6NYVCYNkrUIEHHSaPRbkI3lyVukPQC7DYqrFlBYOLfohpv6Pj9AhxPXoOt161DDZ1v5g+v1ygL
InMiBWOzrwjx/wWMTWZtoIIIwv1si58gSaUcm78vdlcbnR/wcVRB362lyWBtfEkYMSmWKM4yP7Zw
bXEqnN8JbiRJFAguvk1beu0I3QAzjiy7rBdBG3/06SJQP4sm7G5+U8V2koN+0t2gO8BTeE8NjIgm
bWY8c5+6tTJOreq8iWp/EX3fLdwBhnMqPsEo+c1lIK59CTuXHiwlnU8B9jLQHBl55ecloyYmvejx
zLohs4I5ZmH225xTYnMTLzk/aSLzm3hqt6X/77RyFFRubLgGO61D4IiKf46f5U32kfRE/7Ady+ve
UTx742s4g6IJ9tUjFFLHJ19ZOAfyXLzR09WnVcym3lzzJlE09b4co7XjvFS1bptmjom3eJHSB6Q2
5fQH6h6YIeY9U3dky07kvISrmXamSpHb67oRvlGslW9YOi9qIwGKNW1t42TziUWBxEF4K2qov7/7
LtzQNmJD04oZu5OhY/+C/7aqhiBojRuBCjJToVqnSVX8tAZZfucJPNYnVizJQ3++we23OjemCh96
FL76qz3IG5TuQuQ/+Vo03YB5lgqwGbuW9L1/RV/F5m1bmxs/eAfMTtE+xjKFioWNKdyPBheAmbOe
ZtxP8yqmjrw/tH1EZf+fU5lsKWu5T4OntgkTxdqJ8YA+7PYt+LDiKdPXMDGoliSFh67Qx8cxyqqR
h0wt3zAoeF45Md4Up3PC7+Qkf+0jhAsSO2kVX8PvoDx+Tab4g8nL1feQy168LfzNrdy1b8l8lJhC
FP05ksKKY9q1x3BU1gTdY0Uk1GSpgyK7JyhWr1quwqmBUIm62svqMNHqebzt3lddBVjTxzADEf6e
QqAKrdwrCVjKTeHFtSKrqe3Gr4UstnlijA6kXlaQkN/77I4L5KqEWBHTfsuFRJGpMywd4XnWVPyG
0qyHE76YY+OIUIMEhF3DPR99E54FE2l/h0k5zQgDV2bwOI83JsmPZo4npEyVCCVw3BOczRwGKbu5
Z/Ht/F5skZDGl4q5cO6GEMbn2JN0wyv/1c27a60VOI4Nq8ST+iZ8QER08BuK1IZcWgQvDx+HhqZf
j7eCs5X7C975pkgXksIVD+tfF7Z+/dOGu/yBycQXgHAYNqvXx88WrL/TpiZrLfTEglAlMUCLnMFS
seXWfrEWS2DLB4sbu4Er7t9gLCLznGNVFmkWo1E2s++g+KXDYzB1iCY1zQIHgRsEKyONYSM3WP8a
+ub8/Lg0VEXWNWqzk2J7RXJmJlPpaZegGqRvYcB2eRpz7X/xgrcQzEv5pKQgj8H4ogJY8Rkg/JAs
zaRc85HkoR+vI93YNIAb2+GwOXNB3lkE38Cy37W9PT0pETGCYB+5UmM8/6P+pkY6KGMNZdWWRZrK
yFRA0ZURoqYMDYyJjSVvhHsU286noDIHbzEHfbbdRlc9v1ktPWlmYI/r+MBBd3FXPb8dEZao0Nj2
2olobpymLN05zRJT8d8aY0uzb3R3DSUsI4dS3ZRmN4h/rTU6nf4XpLPArlRzFyUUvGFn6mqqNFpK
o+sIJ3m0bbNp3H3oKWukd1/kVqjjls97wuHy/DxZ+elro4+NL6dm8BBmIFNF8hsKRIBvx5AD1CK5
wYp140ULFVlQRy5T0Xfo/VW+w5sKbOPZz0dgrTjvo41O0fylxnD/39bjLXyo66kBc/UIniUuYtve
k05Oh3lOjk0ueqaZyGgy33U6Eo4scctGkBuX5YjtZK7otjKy12BITsygSE7G7V6MOXCCjn1EAsi6
AiJcCByvRrnhkllNu9iC/Qr7ssAcqg4qNAH0MqpMU3WKp7ky1XIsVK9cgpCsBLGTj4iPi6KreWz+
zRgKQSGNKpcm5pVGWwbvWfRqqmvJj1SV1GphzqTuOYENZlhp8nlPBOkTnzShjB7IZNT/d+tpgsYl
pWqU/3Lu9vg2/VkknNaZbx5Q4XL4EaQxRWPqdd0HEwPSu1QDhHoHBurYM5uWMLgvYtEIOoMDl8Cq
mAIltpPSQTSrGbJroGuMuZXnr8vPI21hOH25mk6zRYSOksqekNzOfXiRNwcRcuvo7bm+9nXwaFQh
rfhmvgYcMRk45g6EAFKlHgggYV9E5/BpmNcdJdM0n8L98wnJLo6aRIvnITvhLInycu9sj9zlEuYM
cj1uum/oUZdZFC64jzJZCxIXGEM1HHi8XiMLG/ghFEwV3WT79SKUuhDULSdmtba7ooUlLtTeBaUK
buA2AYuWxHlH6tvetBOlYbegdThn5ZCcoaTq56m/oPIRbgAB1zYY4FkS7kUgF8jp/YYzySc3fmm1
m6e9/TuryGfEE3BWgGUyg80Lm1WA8SGAzgDzLomljFtN9a/vCWUBfLlSq/5pDWgCCmTgfrNU26yA
fjTPUYA83Esh5M13gFyZ4SqKnf/JW5RpzqxOr9cZCc1UHXgIBzM3Y07ykwqr7+Pb6+vjtm1b1Osp
BHJigccOYbJTZeUSaHdxgDR1QPZ6ye52iVZPwkdlJoJQgcXip32G7zVpbUBA9Cmga8tbSh3V09XC
QcZS3JK84TlBAVy5FrdOs8Mec/q/KXYWKY/4XfeDDSQ82z2oZHaiWMIPuuhkrEi+U1mMFmpOklgH
ienN/QgCfKmkFpL8yI1VNH6+Nui+Om10t3lUHqgQfE3lWUC5WOUOW/W7Cj19h3l33BIXAsesXUdD
J/8bDLQvJAnx3cMqkEi/cuQwHMmsZVfjJP/s896KAyAd+eSoKC53t+y/abNyy6w/MJ4FuN7yf9oh
6aQqhO8pe8KPYBO1vBExemVGQDTEwL+6XgzlKbBAEN6zdqmdKekyMmZDCrgwzSXAkhYFwPApg1bj
drdC+j1vwAgdSxPlVLctdjVqv6IMAvFkERJ57e2+GdkSVC7PVwp+bAWshxnhUxGW6YXVIQqbysbz
ebMp/ja9TnCzwooUO+ucEQ9L32LvI5ZuLZIKy/niO2a2mJpE5FbDdPRpNcXj+7tg01zf93vHM7fr
fseAtvWVXWhPcaPztvysaulZuPpaC4NbrDBhAjIAA7zR78wFnvxZdx7x4ob57NfnPFa4C0v5Mx9A
ysCHmA2G/rc4ynKLBs+9IEQIJf01A5uCak32JMWKcxh1Ic4yBCrAgNH6AATXHHcXy7IT0swegiC7
aNFc3GCO15pff5vaWc7rCON0aVNVDTEdXnLxQeG+Bs60YMmjBys7HCuZR9jgjHOhVxijwHfMamRs
P5/hs3KVkGItX4LJLF9xRcPs+uAozfmzbxXbR2VOUW03lAHIhOTohMHIW8FsSS6uOvindhDpjcU5
bfjfA+P8f9SAci6fUEFXFVovP199He7GbvGXlN/qUkJC2bIuerf/TZF6JptPcUxfEWHIcTfKUMLv
GWulpoIuHxiIEmU8ulFID7as2QQexd9B6cy3Qlt+AUFYjehLshtAlry+pynx+/kcsW/qEuhk0gCY
+ryXbfUWb28vYQvwXQREeVIDjsLqiw8c0ZTlwcLzSF4UYptVYqk9FTix4hw9YsZ2cYgAF06IGkqN
cDt5D28zqzFITPjKd/ZDPRRJTLrH7rS7lvcSQ8z0WpprxE7k+WDcLNGqt9bprYnOXKL3yH0ihPFZ
1oEKXr3bI0qY1Uudpa60tZbEGj65v0sT+VkWhyQVO1jDOYwVT4FCazuNpDjnfk32cWW36IE/wThD
Bigm1oP+w57OPkuZs7D+VNF9NtwYRJbC6C8Sn9qtt8hKLgY0c0ig5VIJWaHI+ES24Gy71Q4DFIB0
nwy4nKa0/8O6fRjHUzoa0yI4gtcRNJu4spokRa7hPFxJWo8qrXGiFJlK9+n76iUsVd1w54MTEiqz
U8P+MaMmzIpvug6TcSbedUBPKS9YtF5ZGqCRTS7BmdkpM71/rcF+yvBt9rfFc8ZI+nO76mXUQPPc
fxEUQdiTp8YHx7hDjcxzTbibI7tkd+5ZIXPbaj8qljc2URB3/HM2CLS+nha55Oa7HeFmhaeG78j7
Hc5nfhe/sXug/XouA44sA23PotseJjW5OSEaiLpSQgBHzrxJBwR30XgCeOgnllh4iD3xEKA/x81R
xHqcwBYx9Luho28PXcZzmvCfS07vIgvKjj/IaSbG262wczWoyNKizrrcyhfMo+ZrN1dQR9BRTcmI
rDgA/hptNWWdzwPpo8dYlJ8VZVXXjcjes5c3kXo7UBvtG7U/707kcfHNIlWohy0dd59fcZt+Vbs7
x67Xc5qwX67uIC+3g7RowPkp53feW8/Vx1Rir2Kj2hPtF9GZlk1R6SZ0qne1rP4TnM+TkT1OUmiJ
jqEFjjx3CHJREwvRlDhSA1b09IKGsZUgZUmBxtJhI4BhsWKJLmoWomucT3zlpbh5k4McW6KnID8E
Wirs0dcdh7X36O0q4Jjc+KB04Nr2ebjzgI+m2QTwCQXI3xA5ruuPAwYGSuJqZe6EwWIlf5qAojJ0
z+9cuE2Q2T9uK/MNuxdrKlcqTUvUXlkSCTNlGAZs+2j71+rQGBS0N46z9XWh82e2RtmVe4RazhYI
jgSeaj03gzL7FceDSXj57Rn23On+ian/CPMyT7lBNA29WgxDOZOBdSWd+PgxYeCyGZPIBydU40tU
N9sz0qEZWb0OoLJECBLvDIul6GhOnqOem2bBScOrJ3X54Ex38+czkVfEJuICMXpruJoR/MXmJOaI
0k4NZhL3wgkb4j/1YKHVB/+WPy8q5Vq1CgZDdpSb9VwiQOzPxJfUZTxcbsJjyDrEWI7RyBmJAksu
eLydWs7i3NnowDtG5Prv2avTMsDoteNTRInbHQPa1ddWPR+uMlgW1oR+fS9EzFS5Mt4Ypn2SlXXj
4Khq3UywNDZf2zXW/9VTraVOMx3caAcWmO6MZWrYWMaPUM8BWD/0dkF9bOw3i6BGb5de8Klwdjt4
8212yp1whKHUGgcEbZcyPPUcXzhI8u4Tx2NdBNDqwTv00/QUIqjLLeaz2cLBye36DMd55dV532BF
3DUUGnkmheUGDXGPW74YvqKnP9kW6MXfR8k5p5t8r/26V4gNA7b+JQnm3pwEh7iA56qRa7uuVyAp
DeiVQBypPqgymXpLeaHO7WwLZklaylw6v5PO2k5Tir9aw/ywHzUcvbpCz7ePwjtFatJm0xgZWCgc
1dTx0mAvdl2nF32WsLNKkZDOEh8y9m/miyBZut7SXv6DfAs1jWPaMU10iM01kKGRsIFWOIrz98Aw
rsHflG2QXmH5XvczlfKytkIC0M8ObF0tRziupP7b7fge2ZIqRBIhUuNYCiHVBO0IkY5vHBsSI4sl
tr9Y6zJF/zqbiydJDz1J0gYX7OY5GtzISptoUVEy6e4VfxNUtDzF8BJc7r5Hb49uOktfeumHB8VW
TfRIs0myF2+rJKH+ZHYFvsFyYt90i0ub3hc7bFCFZZ7fErOJzjHwGVjm9yd7HC/YzyP8GSqJjZsR
WKVZKXsYQrBnP8+eHL05MFdoBqi7O+sNEdWbQSluOxM0dthlnrNezcIgLB9W34rE7Ihs0/Ackh8H
yMKRQNnp/CtLbKYihIlWWIb/RCBVkk8UTnuB75aiitsmVOENWnAmhWUafaR9a2r7Dzpk6sRywmp8
rP8+kIVMcQG8uxqF1hah4cxP/leBlaVlpzStjkUZjzfrLbMz/S6ad07mwdu2hNYRV6Plmswhnt7B
TfNvTtE4A+BIHyFBBCzZ5YhoC9/HkiXHB4tikHeyia2r8wbxDwr2Xsjedfy60ZtjYUfAdEyndpcK
DYFthS5AYZ3T3K2Aul36bB+XfZS3AItH8vrk/fqcnQrVCaQMA7Sdzs7ssPTRKqp+dFpgvE0EKIOB
hdgR+I6Ygc6dcjV0DgGfCfZcQzKHjl8cZTYYL0xHNnRPFNAk+mdO527neRQASK+lC5QhomyKSlZB
Xr1u0075NGjgEXVHrr05X1t2mooIY/qyvSHIcPl9Lw5TAFC29XSKWvmIqMvU+7E3fD9hyBS7c3MN
ChLLlYLW4Fc/UE8JfCyem634gl+yCKondhA32qqM1+LsctF7DroyChouZq2XeHrLBmZ7ahAOVHZ0
Pq5onYaAPN+C4ZrBBdXDlbhoTTDEv5YqB8gf4rkno43CKFF+VoLWcBfvqoxl445CZT8Pjfe0vTmY
WRhJX6yo3cWHRPuyoQtKRaO8GPGN4VIE0B9iVT4SBEzbbs4sgUCYnvpgzbBTUYKkkccihL3a9HD6
VcuV0a0FXVCA747y4ms8WgqdrpdKqYhjl1sxMdNGRVwb6lnz9+9b4/40PClZwYR/1zxGGUNFnLmB
7aKDCG52YepfsMwxdbStftbF2ACw40yeH0mu47NPLR4YKmM305XChJShgsym4OWnsb4CLjV7z/MX
N9XZUOsMUpDHtrVojjSIMjbG/nWLSLEMvtC6kn0pseKsaG+3dcIZ4QzBIzDVTXmk3vdRw68UIAFO
l2O3dWmmi+Q2moM0PJTk0et08bUizlA04+wF9cgq5RS5IbrFM/iQxBIBWK9Cl6HzpFr9M8Fb8rpn
4zIC8raM3LWsuE0bO/eEr66G+sHufJQ/+41lmPONxasTe4cblvvoH+AW4sWl953ZNKhOeyQdMLR6
ARuAPR99EWFFWW6MGcYVmnpE8yPSbQXa9s2UKQ6J0bHm0TtcvbcACCjHBGR0xSS6MdKkKYfhfjcp
2mynPHNeWjUNVtdC/cNoQohTh/J5g9vUTB06D6gaXB87BTgORr0a5MLboaYt9J7sD+ghjtUJ8ZOo
I0cIGYsuNlebBN9LvntXkX4/BFRrODdPfp3sILx5H0u8EUiggpoc4XNnuzm0XSMIecTnbA9LsgZE
r9J+frGZ52ggvMT+LMZmt080wvQLOf+boLUw/kVRjGS+BDJVCUgEEdgotB68KmIVyVBsoAll5le3
B5q2KUr5jyO+tslKEfxOorKJCMkr0XNWpUZMuv6c6475kujf4EUtudQFXZjkZz33ED1rylP+CwA3
Gy/Z6xd5zurNb07LucdwRNXaKamB47cJgHImbUnF7gB345CSvh5W1nT65FXdzr21S6bSpAokBzVc
hUj6/3ydk/aQkrJ1KGP6SmgJl8S4BIIKNzC9YVJN0UxN6wvS5kdD8EqcR1uuc+1vPDgAqJi82Ese
a5higltRdKgvJlft1N1Nr5wb4RrM2soZcAbfEgRoxqu396WBV0IeWMXWLZMnzlhYY9kym5SMsHQ5
wo5a4707yQF3iFe2r/1XKo9aRIlvtzoqkxacN35j8Sh/HFnMZQ6WLZmd0R81n6EJxsKNTguib1Sn
tt5i9slGMQV2XVNoOQDgVccN4G2tOTyfT9ChvA7MmaNEziiM7HBnc36O8SIAERT5cuqa5ij71mbA
zneOo1aRoKawrWdkmn5fZllMqsgYlLEpDzxvJ9j7rVyrwfsB2CBL5KEq+mGvNc7W98R4qFjXW868
hXLJD9KeoR9L2iF9uO0Q6HUiJ/cvNQDUBG1buo+V5HR/u+uZKHl6CBGjHB5LH8w4oSt6jSW53I1m
CSfhDH6/VfgOFX+fp/23Uvfll8HiXV6/f/ATbsqBJCM6O+7gpKXpRSU6VGFL49mZzNiFQxl4TpSd
LhCSJ56HAvJ/rvvEwGCGdIhDZUZOUGw/AtymxpcyWrEEUVGNBwnoQsfw938GaSJ1k4N9Gg8hdFJw
HpzT7ZoO4Vphsa1BvnzC+8Tg809k9Zi4YbbCiwWbVgBznCGwfP/EXU6WJwslwZ3cWDQ742cdY7qj
ka+ZYyd8Vg+i8JyWDy3kZdFkULk/QQseAVTdcOJ+sD+RY2QG75hKEqwOv5DCuUiqQYFOQUaZOerz
NmBxNqsreWzxK68ZoX0Hhpl0Q1nnfEg7GtJsNZPWWSwQccR9xIELZLM3QNtqgH5rnZk3EbvToNUy
Y+ROJQ8RHcE2u1jjSCQyDlToHzha8n4Ca6BJpJ+bpMF8HovC6Zrsx2HB8zvA+E6726C2F9k0siwY
YAiBZJ6FzUsd7rlACz7KpcKzMX0JrgBq7sZ2bpEsy+dsizjAFBTtpH1Ssg38a5fYWaGhY03+1NKl
MltgQJ3WOjC2xG+29wmimI9lIjMIrln/7onLoHomZ77eg/29aa5rNQyIDMUkN09UX7T4z4jo5yVD
uUV12OBC2yKTMYMXOXUlORTYaoxYNjbRtoileJC8dXyyHVKI2hxparn515bw310DTqIleN9a3zTz
jOp3+YsJDmVPll9SzaMWpMffBaNSx1i7llcM4izvQjSwEmxdnrmdS7Wk/hJT162f3VbwBQnWTLDY
a0wDeYS1lRFsftRZ1LGyQqPSLi8Gn/E5hivvSFt86Z1aF5aSBhzCBgI+HSM2fozhceXuAmMvQ9GQ
/BS1Q72gyxISTs+NYPy7fyNuiBLKbRM8RE4LgXveCYM5kcurRpg1ncaI1dXrV4Cw5CqOo56seQPs
nKpbDBHslrZGKu1iQFEXXfqACVY9hwGA9FEeRTreyoFwIwwUsAc4nkjmFOW5vSnMTZ6Wjz6KVHLl
EGU8T1GdCNa8T+NwkW49Zl155ScmkbiHcOh7WkL27kI6NP8AW8liSdCW0AbFlHTvDiQGAxbxd3KS
4/5bwgsSsFgKr71T/Oc3sndF78KB7K4l31sGi+MpQrI6fCXGP2JHGKJ+VztX92UOvzyYK5tasviE
NsvTDQvPSuEJrLrE/qs5YAK6ih8Bszy2uXu2XaeQUdSclLYc3BXMC6rFtpeRY8gomxyIU3K8tdm2
wL5aLIUtIkwJwv5poBSNr0iFsiFfwe0Zhlq5+TFeAotiWXbwAVpcCIosvI9hewlV3hO1zGtc1Ohm
2R+CDigO1t8Fq9XObKXPXeGAPQeJNer1dpaFO3Jzwvq4N2fAH+zOAbLx6ckX4NiYu9VwUmcWZguI
3adS/GKje+K+HPjf1U5UKXFKu+re5cHPcxIUDrrjTEsCMFLRCXN8+4sUWu9Z+OjYFsoIWyEbfnGh
O12SU50haHI4duReUekGBZvUipzByna42DFu6UTiiU35eq82W+5HFbpTfp8M5arz1/NNAkcIR2FT
4DRVeghPFjYlzWt+aziX7MBoU2x0/D7d7fiqtHG/e134U8qejzAPXfj4X/F2VdS8IR9VbDu7Uigu
RzIeejSBkWMAhRh00fsb9slFyMDCeFYxUPMc2Ew8pPHl4OAofjBrjKNWpemGzfa/gbb+emwFElFg
BU0158iouWON+g1GzMspGSoMnONkYxh+seeKf6dNbtFHzjmIcEPCbiCL0jO90uKTDHeR2pVvHr/L
RfOFB0skpNv1nkDHWOMWb84AO+5dNziI3Jn1yL+TNHf0Dr5r6mPg/iaZsyjxSKwGJPACkSF3pi6J
KjxhwOuDd0owPRYfUGcisbnFpqCU13FBrKi/2MQSL1d1Nn53BSd9/JFer3g1oPJBNoylAZ9Oj4mb
D3WsumTIS/VImJ7KzesrdomAOKDQcyFOzOyMto3yV0GVxCQyXwC4VH5HqV/GRvDnuuF7g/+zCJk+
hEbhPf7+uHpLrbY8+BHkJ4PI7SJ2tTqACEYumacOYrAS0k9QD+DWqb/I6fwHIZUg5jOJ7wBOHRIf
hwZjJERiTRC3vzdr97l+ELmB/4/9byNn8lDyWtZBw7mp9LX9HBiL0DUMQYFZm3QJBwzBtRhwIGHR
1LqfBoBsn8/IeuGCFtWN+O/DAtVaxKLkSgfxUf6YGwebQe5R0JOWjKXV9wCvEPOaJM3yui+CMgLY
EavhoC2hLEDmWUrkhtzveIdjWvjiKUkvQWXTdzcQN2Yo+aKB+D23hzV4saQ7oYN6LwsP+w6kZbZ5
SRUKmGhUrlrnOTc+Azx/tT2cVoOavAkkZQutNZynt11+nh29hkfjdoq8EFUWIboaT+MyEvd3Mfwa
iu+enSIcVZfjKOYG9gPwTyXRJfefkAMGC2YK5lhEK0WCF1a55BhjsTNd+xxl1dlEYBK30VH17t/T
Nd6qwZqR9csvTGZcNcSgF+W9bQNVPzUJ/JATFvnsvw7+6B8Px/X4KNEAQ+FuFC/+tZJB24BzEvMG
e5t3QbmLBLmfq1pDGT9drW/1ZAdQE9R6vSnoagxFqcpGy9HyQFssWeMydFw8Pkvi/mfXAyLU17HP
eXwZ5Kif7gEWmROZHfsYUwFKkbjnsbuGkxdob70oWRmLnvsIe/Ag6N+8zYT7g3n+7ny65EgoweBk
vDvILfN7JQQkyN0W4Vv7bgnJNCL8YTbbSee7SkdnW6+R+c+FupGnmXABoD5EhiedfIVKEsm9WADM
1gfkw74YfNzT4hdxg5YPraP9+pfoRx5snJ7yOYXB8Dy3AQNtZZTL7qTsBlTSOVfU2DnujCQCWXaC
vw30omCCUX8o8p56qgiZ6Rn2g+0gaaAiP4E/5b8hube+j0y3cckhe1xW7TE42B1R4MlmnXDW2ANc
p0h/tt1zhynveHTotIO8+HZBVkabEDqvxQc5X5sVAKUvpcY1bsfJOHigb7KmSXlcG+rbXsZ+YR5B
6EqcFOF7hBywz3MELusebx/F/YxUqnqVBNjct59EHoEXsyZ6f2FVh84EZKwqeUF3u4PHYf0N85tX
ktYiCoVddFUx1jxSzjAdXIRzrUsoYE1TGgHYZfPMvxuMM/T0c0HNcRMuIjYX915IdqY3TrBsVBj5
HA14QZgFbSymzIW0O2+wxmA1+Ub/Q89OErHq2yq4haq1LP7mBS0JN1PwrtSL9wmC4tKPVCphOiFg
+CAI7SkD94u10N1AeRYckdS2HN8eaxcskQEyZ2xrSXkdhoiyPbGxvz2fZUSUmSU5pBC4ZMqnWz+j
TovZSYq1oNDojnNIetqBfRC7O5K8JgFDg90qNkiKtwf9vYVMJyIXUNhAVDM6JYFmOX96siymwZA4
JK/bq2CNSjIW60/iggpsh+QMLQwgEg3CYUO6Q/uB9C+lGJ9+3YXlen3DttVpaW409qgSPxSReGL6
8CjSkX2A79+TY1m7+4cOR/anIh17Pm4zVahcnImAREjC/G5Te7hxtZXBALijBw+DXPBqjY843/nt
GB7akwvP957eFofOSjk6vFYaUcjH7HZKhIEsIhEBBaxTWntdCAXcBlpQ0txCVPzKngjKWya4qXCE
OW7pwLlg62uFqvm0r+Tf50s18g0Y8INUOC7Bjj8zS0yd3jysQUl09hMwr6RxQWfmLPoEpBLNmTev
Fa1ZH88nB965ko2au8EfQCVNPF+EzRQ2Y3qh30alXkGyyTggXuHGUvszOGA/twM7OxKBPa6l+h/m
5WyCmSJV3Mm8QBXuqOLqoCLEYLzYt4bqS1QNx22nH4pjBPj/6/uBSthiGgM9FsmdWebOua2QEb+/
I0m4TT+chW3jMYuzrMwRZGdY83M6wKyEgUVC1Kmg28UhszU/qUG53g43iFqzsOd7O6rtIfD8fJFo
TE1o6k+Cs18Fcj0JvinPKg0Q2BlSq/HYmjdG0cHaU/jnvdjnUZoECxTBGApEANVXmhOfF++m5tI2
j8asKCvMmPV+eQrKKxlZF4f7eqWaqEq+B69oK8xE4m7IQTlbzoHExFuYsEeepApcRucxMCI4P+oq
CtqLC9hfVuwKu5ERkAf1E8N+mWf3AvcpoHZtNsLMPQe3lvSKqpEG0iI/LOFmkGQ2l9SqcV+QL8j2
bFOoKfvlLwrWwr9nVsikzSaP/X80ZLog+zoIwNbS3TylkzgvCyXVTVMmkd2LEApCSdEqTixhc6SP
954cfJEYonQLZRHwDOKua4EOryrYnV39bhdl0qB0n8S7uBm5Z8rfpyQoU9gBiz512TVS25q79gMa
3W28MuukjO7Vgwqq4VttAsogMwzEKrJfng6UOf6fm9jy9FGG053XQY8XB1NeIGDrulbZxQwadSIR
Ci7mdJCEWZI23QEVbUDHzVDv7CFDYGah40MJtMYxiJq0c17Y98NP9M+hknpNQSstgFuSLplNbPWA
y2n0PJGRdx4ZydFykF991zctyXcLSGKR3LaLaPhxmzqh82wOj1Xf7phnVFX4/y0ZmZTv3U3RPK4o
JGHDFACkbmsQdPb07gXdcq7WhnO4Tz9ErPerkGfzYZIUGtg725KArNn03wWccK3eT8rkfY2qrtEA
ujFLA+j+PDY7s3o4mJe5e+7VHmZmDcdd5H338dW1BKxeanSmZuvfEjWa8XTAihserhP+YM+vo5PE
c6Ub3omeSrosdJ4A2IRxdeAXCFF5WND6sSMHyCAXkpUEVDgx3or4Uswlv9+ZMZhobpaFnm9mW3uW
7DKpLdYumKzni0sIQG41FUu46yWvKIhSvbVkccjNzW+cMiiW5fWvJ2H+6H29f2GosJf9rbWQ/OyC
Cv7Bk8SXTUhwsH+tNcrNPKMQ2oXy9UFwEeuWhr/hJylND6Lk6WxF92KANt49MxMWi9/iM8zVHIJU
rXZQCgNE758RCIDnI0j3wTD5xmr4TNj7yqtFuHXAeFcgrNMjnCkzRSF2v8/25N2Xh715l5lxBA4F
lvIdKHuzUPvFrQXVLU33Dfvyc166O8R9x/6PMMqGmji0Cv10dm8D7s3OhHceqfBUPQVoGeIUDq24
mZCMOEMdXyjXZ0ASKe3KllmF5rmEk61gWDbZbV1PYZT6To77uK+ZQvsAXb6MW7S6Zj5dHuqzsrwU
XahUgmJubjmP47POKk/YNmTMXUqwE9RBopzI9LahALIejI12940ZWHt6fiCQDtpafgnYBkvK9U48
6c3Xq//lYwPuPkyGE2GtNv9N1p0tHD3kfplZ5rBaOsuYPK7M0zlDH7E0gi0BZZTQSku9NrgHeRax
uyJas+FliXI940ixXiqF5SZa//xGME4PsZk9SbnJ7ou8G+lQBK1IppehpQZkp4VhSQf6k3UaTAst
RA9+aYdi2xmA1YaQFe5qkPnLLt93HjM+4Calr+L1Hldp6RRTvXDw2O3yETH5I5vgEjRqO3Ktk2yU
+pnsYgj+fjvshUo5AYwdobJFYO2lgXuX9WYVYSLCCFnmIjBRkCNVZMgjjt+aQh1QtV4sBK8Yq0Y/
Kn5Wj8MMPj/Z24CewnR+/QCmu2XjPFK53iSettUk9r9pauK2us8GJmBV9wmbynaUm1DAWL0yCH1l
8OjOfqn0WLm19R1iSJN+0m3Uitai+rXVt+Zjw12Sss0nI93pbJxJ+j0iwkll1QcOoXUWisKr0cRK
02rLrvEnEBoh1ergH7sDwfXe8BFLUMC4eeEBOzDuR2wZFheQU5fT0UPmgm573xHoWLzLS2ZfhrCO
tiyVqoDFAP1etBEjYdIZMFDlpFAYPbAztbETmL4jXO9a4+e4L/LT4cJULZC07qs4PL7PK5jU2Q4w
4CkAiPVir4z1nC35bWgOKTNUEOvJVdYL96dGaAIAxFFO1iLjIYOWkJ5UB9IQdrVKFfhzl8GC8ON6
Y3rTlbB9gg7UIDEL4tfE8NsrZL/CKepH6p+E4I8UYeohmmXGPaXh5vrtQ3xwTSP+SpDr9Dig0dDC
zXQflrwOFvW+izer9R2IN3hP0FbYGMh6c80+OtTMkn6AohcVqyVG34XqrEn/lEB6vk6+iEKU4EJU
x61rBkluA3df5TOYHDZYDQqkBV/67/ESdN7L1ujRPf+4KE5XOl/HDfyONjwfhPftX8TxYtT3N/ev
Ir9Q1DFxMmBgZwzwm4AgAlSr6V72Z8M25OLKLdZesnv4MQqePBFw1qKyw2XVKO/alsiELNBk2vv6
EXsaiIkyWKGEilRxxTM1jvWIrEHRbYv1TJmmZSJW8huBPNyUxaGw/PY/gyGP63YMnAFxaCCXfcRR
DxpDIBSA+FjKgym33BWB/0hX7ZCKhnHb/WRYCLB7z2Qxvjs/wdeD9ZBTZbQ9UqwJxngphwK+MupK
VesvIlUtEEhUfuq5vnlhXEBSRRXkhDAZFcz2o7oNik+5cQZ546gZO+xpskSsINo41+71SNC0kaQJ
/BoLcnEB8qQzkWWfhJMVnA+PDaFELl2JarXXJmfygI+ChuYFCVGz3GAhOtdlydzTGfjBVNaMS8c6
wVQVaix0Y11F0e6PEmqEIjFwyOZhkKv/OvobS5cyxqo2c5n+mYKPUH6mSFl+LQsdH8jt8Xakayt9
6rp7fpXCHRBkDB1+umYP68+UGJgdhfdRi6bXLNUOsEeo3/co7cGLFx+N8u2I2JMSoHgnNkoZhfN8
XkDcLsqO+cNL5Y38sBgbREUbWtxNoE6P9XXzx2wj14lSoiCZAaFXL4WOhsggwdXGnNjvBmMkHYj4
EIk4i/vkvCskTtr1Y45PEVBU1D/F4EdBnn1t6c8qbFrLeiurajOp4K4ERg8bKuwY4xM4w1gvq/fP
hS8oBr4YEKpjcvvEeV8RIHL7f2rhHnJ6PKAkszUYuOBjeKPjzyQxMoDpQS1Ix1Es7JhxWNsfICBX
1506HksxWfohfC4lEu0LAcvYEVXSUwdjfWNR3J8uY/ktuxNYqp49VxeaDUVebvsecOc7PU9SxTFd
x38L8c0ORii4i8OLBFne99L01MGPgIlJgJw61xvTi5A2mqlonLFr1TeKR5g2476cEdlvFya2JAGU
xllzVXqBqMG32aqRhbbcZVyU6zrCDmQx3cDwXkfzMgZNrYoS3V3Lr1akjyuAMB/+GwMEA/GR+LFz
l4076zYAFoiu5AIBegLfGQuIKhEpTMiHNgxWvNggXCpLUbg61BH9w/BbvE7DIoSNQ2+9ex8/VlMk
U49Vke27c+gT3T/Cq1DHHyCja4/UiUhHxNwW6iIuEUyzcwB8x4ekHgR56bI/hV0yI/NwntE6umu2
C2sS3XK2RGgu5oel7EG/u6T5s9AvC/EkI1WgHtqGaUScRvaq9jw6cYKkc1HDgcW8YfuSFT6/ET6/
GbxwxYRxJbmKetwAUeB8uDEj1ONgP3sLqw0MidTRHgXqJAiPerGbEARcP+8D1GlpzF4Ur83XwvMI
B+AnvKVIRwC8do1y21gmOTNQX1OiorChY4oDBq7Vu3OP3o2XmRK8SmLSy0V1/zz3WpBi4jsHCiyE
/ywchjUm1pZjis4pJRSZKd2YiySLIEqqdo/xEwbgZDhLURDIvfC8MhiRWbkHZCMMyKEuRDwIOJHZ
6q52OZ232Jj2YJK4T5JqwLzFidYVvp7J/pVIxsnI6alLHWdNTG2eWwAjJWLH4LTlWrD/wEXzDxD6
qxgVHoF25Zn+QTD9TPGaEOEzLfQkSzblJKD5nXdxrypffb0OR7BYItnrZnBEO2s91+n9D/OTCMCA
bImRUUft25vTcfoGY2ZZRDcyzmMDnARbVmxzTG2HFKYMH2No3rGqhiosVjC63VBBqZTGyg6n9L3l
7+cAqfmzJVDD3GD3uOrv6jTXECbtV/tKS+wN6dQ3XaT5FNQImXO5QmISo0QtoV3NtlP5zHYgVDtB
cu5tQeNaKLpdDmMrJAqDOuWAtZOfSSZUbBE+ISDra+9iALIDmpECc5VmjJPBRFAviWTjDryvZInU
8GJx5I3g0rpDYq33bmWC32a5fyjzKHZoVOwqIlntrFkBUcGcUHTO3X/wXUYjILqWyQ5+BBb0wYC9
z+hzir+O9nsJ/F0mPV3pEgIonDwKgMB4fND+5Urj4iyepJsyhxq0KFXKtV9d80KH8eXlyrOxh1Dm
NLgiXe0gq6b9Ze3hFyDzu+Jpzby2eKGlYx8Bz/Y9dW9BrvCaCK+KFW5FsK0xGvDoWvao7AZodt2Y
ySIhAbN3lIwpbCpGKvqw5M0bJBHXCA4qUs4Yfv2zk43XYAT2snWiiZMpjbePpI3RSnT3u+ie+8N/
c0MvXRuBX7+eLZMsbMlF/M57KTXxSGciUgQzu5Pv/wY8oOVKCsBaUGWSdrevbjCUD5yHpf7QiYPE
71O58StzvOA/MFRMbT5rElHkYTu8YZ0Fa6mIonvkT18lcB8FHIOM9MgQmPeTJDrjgP1FaEDry596
9NdNJwgvnL2Krlkx8JRkH4J2toaYThNsHhtsjA5Idhltc32/wH+i8/8TF6DGRNMgZzHZ0Glo3qcx
9Zuhv15JwobjIkJgKf1ysr7kYagsvH5WaRscjAG+wMfFSMBytVJhQjs0lyTdL4hZPPKyeSeY2fv9
Ncf+51RpiHTEqiEjRNOy+2RK3XX1zoy9WHrMo6FCFS/E5az11/3LHNPz/auVSiwxOiLyhuEHWppv
AmsJB/lAlTKg3B0wSFYwnxXpv1acLBPxVG3q3+gXINObA05JosR9l+WZ4ygHHHv4p/gKm0I1btX0
lWLToTqiDmCr2lnSGq44xX4cgIWgVHL8sU+ErmuRTz/F0QGitsvLKoCgmcjiIRyqU8kQJyED5dEW
Sq3iStgRsgWCId+yYbtlzn63B3JjAgWuxYWSWdK5wjkdbrE2Z1ixQ5fKAVH8H83fwf2AhJq+CfqJ
guDTuJxBsP4+5wS/Pv/LFnCk4FNBhBu+eKD6Fae0ajiKucoaPPAR8Bs34RrFFzy1Gvw91CSO99qp
mAPZ/rFLtVC1aWIiDNdwXQ98RYwbD6eV/zfVuPxilSegOscjWt8IqaoawzYI6bSwxO52IRrR8UEm
pOAGf0+zQu4P0cKdGTC+V/7F02Qp8I2qgbVQWlca/pKUb3pCTCN2tfWlIJMOXgl6w+UH3FPhExYD
lFjR39TXIX9poyuzFRlMY+iciIBcymXbcW7uBBT2Cd2rEU657GbA/VdaHqTf9LUbvIZaEZgbWivt
MHH6+wtpBQHW8wwEPi7aD0b+5qei/yE/7v4IMicU7mNQjD5p77p+vGspnHTlNI+206GSt7amrNZ1
asEFwy8N8fyjY44wTfLDTrVeIdq+9BMy3sH/Bi/BB+H3rP6d1n01BId0sWyDcnN73II8xpUrkyPE
sNojqQgkSHYLugMe9dW9bictlKD2+13d5YVG1LASCEBeH8dQXydMIhYif1LK8qiH74d8OQzDPTL/
9NCl9v7wLG0jS4li0Lm21ZIClIofuHWQB6VU/JaXTJ5foy3ckiscsxZyjyQxdavKHuoa20ALjXVS
fEzd/0k6PTWvJCiL5ZDSWRkcC/HsPztm6L5+GhxdzTfHbWJhL5wvMN4a2roFr/76Pa9m/hWZ2AZZ
zn2esVhYywEIgOu0raZM9MyXiM1Qb4o3gNdNzu4/arLlLwrAYkBZjCsxjhl3/S7RNZg2fND13JFl
W0UK/55WiKnaRX2DvegLPHmtgPOUMarinWkZ17WOk16t6Ba4m6vvXsrGkRoUQjSvI0jNPkFWdLb7
zsjHNvjbzpFEenyQ+ZWB8m1eVVCWQCJiT7u8LRo14eJQMDP6XLYi6rk6Jv0mNhzf4Ab0dHQsKopN
edJHir9rltcgzZCeEDwmmtZZQxD/e5LYs+Ft3d33+DRbc5zy7HQlvU9R1DZZsbAmYF87mrvXZImV
CCX91RenJKGVBAQDGeyhbfGPd/577d420IO2nQ+1g8RzInVjkUP03dYsAn6b2E6+HbmI4fypCU7v
9lu6g+xE+I1L35P9fBO57VkKcbaGTPgETZiJrRtkW6eC8WQj9bW8NE5UxShFnZASJixRKmUkkA10
ocU1yYPL7iorun5hNYUzMR7W/P6Lch7mCUEnA+xcG1Ybf+UYqKzYAK9GtiTPzJfJKHzhaboXIPyg
34aEQjrujwRMb1g75UNKD3ns9AYsd7daglpeareDzJDgXK9PgAKCOR3KYAx2eoHyK9TslDthRR/x
Sr2+upu7irKD5L7uhqKE6aOcOp2DiO43zHc6s5YFy0xeNJvXsvI556r+bUmhw/B3dZK+SwytRQiI
oZ6+YkXeDoFd/rSC6f0BgT5J1Ihqyq1vhVXENS65IHxi3Ps4vKfSLArsQoN8qpo5cXxqGnXIe/Mg
hMWNWknjUSzBg8a1n2ZAsyj9aHiaWs0RuYaGPYwSoVgPGB3RKIj8+Ekl5Mqr4pdph2I2WBon7MIe
4j+MApEldiocMLTuYOaxZ2Rx7VPAWV1IjpAHPYp9WvwKpC8vXc+ZqIc+Hmk+5r6DdptW9ab6HTnb
mSybOgJjtkvyiZIcJAumL4PjaO3vwEHIamwZuCpYWu1a5Vt/IBMyGgPGoay2rz3GZ2GhpG71gwDQ
8vFwZOIubWn6gs72irA8u2bJtFT6vnWlaZ1C+5/RqQsFAiGzQsWxFmXY6N9oOWujDPl+YObXbeuz
T2x0PX4QYIR73waPNWRvLBwWiHLmTrMZk5UdYDZMaQp7oq71kWiq+bOpjalKXaYaMSoa47+Mq0Zj
LAt5qOunIa34KOEkPyUTrd+hHphPBH8djHrWWoGjTMPEvt3X7LcaVRuPrpCE/cnqaUtNRd7BR5vC
MnYOP+RvFBPTVcrf3BQI7L5WsVn0nvTCz9dsyZQ0coIfaLJ3tIAIqpwnL7OqoNEiFbYuEqL3cjJL
AJv+i/G2upqYFpHt2eWfC8etF3XtqlhgsK+KHxmaQ0mwTBGpc2sPg3MlVjjQlkmFWRPeOSwg/oal
R1v0HII1ezaFlbAICwLJY5z8NgG66Q/Pj7CpncJyW3d+qlT/VLOo4RULqcNMsV7iFghYRf6h/jRd
CZzHySS5zn2SyxIqmKBD2n5ngvBXL6/R1CRGLWoLkkZ6w1VVmbdOXSnDin0MplJnVU3z6FMIYJka
WoiYAYp/J3FPTiCN13j28Fc6DC1FiUNSuVeF9W6KH+b8N2Z0aKySvy0VNaPuaTSO94xft3TwnpNd
4um04c8hN5oqxKJeSrxVlyBFOkd+kFHshbv7tTIu8L5n8t+cilGEdDl3RxWwBHhKK6xP6ZgdPDoS
MH20twDK4Mqrp9lWZt8Hb3AGwM4DMZTLmwaPdeZNYbCeI8yYsfdu95qvKmI3Bn+RKjmj422YAqk1
GQZjlHTO0sIbv1crG8wM+S0jM6OgvLL/sE8x2aFGihd41tO2JvY2vNbvXJtZwPu3WXs/11WPEilv
yN/Rcb9q4s3A62IfqMYhPlfFtWcD7uDyRU0MCDL+QXPfAsXFpfcvW7aHpF2j6HIX5Gz2I8bIeQk3
aNmk7vwX5yaYy+NVYDD07p666K6w7syP6FC7eJnIvzC2wEiteYNpw/BHU+fBY6fTuXWpDeDjUIj/
b4vqfGu0No9RmhaHUWnJ6UVgxBE9Y5LjwhqsR/X2rEHaI9t/UkPYC4cmfQdKHnHjXaG96o4W5UD3
gCwYfXNEDFIkZl9qzxgGEoUdPFQMKhqbgloVfFTiOsMriuoZ2CrxRwfDn+YDbaDH1mnk4ZOGklMP
OnFDxJdJYrtRLuzKdqvdk4uIxYLVjSBv+O4DkexAJg8sRCJ8u9THr/1Tw3aiME8SsxmNySYOQRIg
yuev8Q7AiAAzR2jSPURzmzZc7HiGeLYM43NbHOE4qb1jrz7KHae4L3kDupyw54/8USRO+pObB3CP
a1296++2zBRp+27xONmVXndduYkS2SZn7aOre1KSUdwh6fkjXDbJcgHb6ugIpvH0jmz12dy/xn7J
lkki5C6SinxqHnvAe+3lJbh0meKbL1t0UgaNufx/gno7hCNRULJxXpd6wOWd17UQDEmRU4bdQZUC
CwWVLuijghiM2K8/EdfFSMieS1Hu8D7MF29I+bi/MRsUCFzms8RmNYzv4i9U1PtB3Bu3bJhRHCEk
0FcjD2zREdk2PepwG7Ze+jVSScbOCI7lx3q2hncAjZ5nyhtUWfXbVvKQjCNTDOBv2kcCpS3tC5Tu
aB9J7p2SzjvdX8yrjC3HGyVmW68M0fkVdXRF+Rj1cSDMfywPAWA7DBop3GcJ7368PAZoqw7srTvb
MlJHi3IO5Vul5gRFsLwxelpAvclwp5zyax1PSARP2JGv6dbMMOcG7w7L5A2qcHRkQMh3zL+hf9ps
dmkytsYIh1VOW/NPobXp0+ecuNYefBzJdlg8fzpECz5fx3hMH/z9oh+EOFXxvrLgkGJAMB2+Ra6u
pdt9ByZ76zy3aB5PP/HuaKuMM7nxNABjtJZ7Yd8qaV1hY/FTa/3vr0b9991gEMLBdfG6s/ZNM8/4
lSWvBJcD2u+ebJJ92DpMqkAwmqivgfjHKAfvOnpMKP3BPrKK1LCtuW5WGoJQeZOMhb8tXGSeoX4w
OKUohBCVIssqTcain3BcInsPyquUnWY8jCi8LJG9Qduq9Bt3S6c071zWEEpT31ieDjXTHQbr646F
VKkXb6ytagh68SJoiAgYxoTYYALTxBiOV/peg/LQmQmYj1GjLyfCRPc5HgltUPSxKMEr3khtI4U7
uUsMbVJdN9HYhritUcgEv+hP383uTYO+2MCxPKMlk5JdHfF4Thtt4/MSEUa6+Zex8tQmItY8PHs9
Y2Z/PAJdoqi2sy+3rk8/1g5xksH2Q1QU9kHC/LHYt8tNs4GKCzGzQegc3sm4EOMmtT7lGMoGh3d3
igPREyW3Q9+wTs7+iECJQT+Y/YYCZTNlr4bJ1eOQtTyMc8XSJv/cP0vqpCylb6yBG+XHAthtlWn+
dTthZs40/+uG9iknkxdShVGBQhPFFZdqqiDeeA6TcUcrW44ymemVWQz5kE/se8rvnDg2bizDndpk
l3EkIpo2fihwhw8krRvdSo/uWOIjtC6Vt7r+mWLb8YuexxrQ43eLezX2cgZV97IQLheadmOqg5tO
8IBMIqV6t9Sv3FjjQ5hQ1YT7PHZ94KP9D1dSIln9oUuTC8OiCj31bwX0xxsvf1rhK7/XN60VlJVw
KG6JF+DIvEvUmHOVHKP9EFcv4PqwTLWXNlAAIpVc/e+BjyxvpjEU+lGvFuHsnQUJDedIdVDZTxg6
Em99JSQl9hogJ+9qAS8hq84j6EHkjDW7HEMuMdKpxhvc39qX/YUgNDxm4vLVmDIC21U/yq3iS4Mx
MHgOM6NdB4qalS74yJkREyvBmtP4PBpROJB2+UROogX4wxx6x8nMOyAsTsJob4b7vpWgdS2JEkJu
Q0r7qIfp0AYQhdvsXBuHCVEcBgaNbFiHIpkPwfKyBbhb6xLqNRl2E9668F+jTGib74QyMVCAPgp4
0PcEBT6/XCpNxVxX7DqSntamCdok0dFDLFHa27oKd7TUwwV2m/K1S92x39nlZ7TvyS2PAWfYBGl2
U43c/kcPYrp3ThLi1u7sS+JitlsicPrlwkypxSUg2h0o6SwlQjeJvTecDyPI6EVn7NtNLnyvGqmK
Sq8zfn/Bw2Bci0GBqIbB9ur0Rgy7fkrndOgAN8eNeYsn0jtqoYJQByy+zIc40F2WVsL1uMoGQI2O
SRtF8SX7Bxt9KUQp43mOAESw8mkO2mT789VyAWf4u6ZLBOJmDUoDNTcN1YOMrr7jLVDT7U8fmGJ8
zRw6UhBZZbCHzITSitk665AQa5orsCSEd9NviMa/tjvZPbFHORbWGWCJFv+txEJX2s7UGyHINfzY
nzH18QcZADGgDIv4synfKuXjKlILQc2RmXu4iirV9FCXsehLj6W7fdQQO4dpZgBmcPE2o+Vc1aKE
FK7pyrkFWPUQT8ToMm8UYbPKMpe78TUKO4SzwbUo6BL5891LairouhQVb9kgx3LG9FgGaBlTrCOE
s0HZ1S8mS1dirxODH3jYuTu1pW9+/0m61R5f7nfz/IuIaWEUtkp+hJNYbOUzr7lcp1TPGkmP8ct1
YQX6ghgJojThB78G4HhI+c2TYwSoouFrP5zzX/2vgXLSelBJ1wUScz8wdFZXZhzYN+DK6hMudNV+
+5TdDhjlrBK4w7r6uoo86taoPjTBPJlX2VjDGj5FG2r2F/dntkkXDmDMzRWroskU/iwBd9YhK6wV
u5gcaGScSrAA9CqiB2KjYTtuMJtpb2OTjk/oyFJuS63OuXmJ/LCsnf7snsE239Bsrz1haOufXt4M
3v4aJuL5YusOmyzip2+Pe73ralw+R6fN2fDQBCzS5kxuePUCAXzGMgOJoBq4DQUrtkcmZcrlIOto
3Yc/fl8sYlIgHZ0B1mdInPh6uKg9tNEZguoih5HPLqrEbBiW4xTmMik49vZIfpnIaiV4P8jM2xpM
oh+L+Y54IzeuCIKjn6+L1CWUuvMMIBYE7lK5NHHfAlkDe+naxHYdtH0PB100w8uW2mW6k8nzvtMZ
7BY0vMzmk0/0COX+czLX2QxGMItEbUHA0zQFSfJ8TmsV7yOpjUsaOld0cfAYWlwnk1q9HbtfebuN
X4EvR7wgop/+xeZ1yVvtrCB53k9Pn9X/DkoWmwa0MR3Lf4QVWY4KpeomSMoB/LdFG29Ezpso5GuX
eKzkkQIVgJHbjNohdGNa0qm0ymvT42KEEWL3Vz5geeP1NSsNyM6TD/uNuu4PkEZ8IPyuqMxVv2/C
+4KupwIie/hNuQ2/aHm8LuCpkKGlSLDatKfg2FIlukHkwDKgK8uAoAQWOFb79VeyjH/bNR653TD+
xfzC9YdUrraiLzFO++vVXBgX2kp46qKJVlm0Vu8S9Rfo1DhdsxgPdOuo4gpgmzDeEAv0c6ykgj/5
OWOK49i5+ngw0KFBgqRiUXeTeb8Uwk0inRr0tRLymLr2bXLiRS8vo6rZCtAaIY4ElHEyJa5VjRaR
mQNlsF/KveSIK8hl5VWcOPK3gaYtcmAVT5DMkROX+HCtyVRySBwndcZUuKCMbRbRtGPm8GHWg16G
6Xj21ZgXalfpGkgfeJiiFlbOI66DY1XUCtmd/cLSHu2TcjL4mVdFHBxgrFTH0uPaUMQg44HE8tfc
h0423iZPGKs1Cje32qkz0GBdlSNN1Gu/EVgZoN/lCoDEiJOZJfiHR+3oEbonFWGj+/Bg1iOVsyUL
d0tzeC3hK/g3RmboJDHMcfYNFbFw151tpzUjr9kT3uxUObPhPtPiX6s+6/UkotoTE6D4f1HpVUzl
lYQ7PMXZsSt2VXVESwc6HDBo2e5Tzk9l4DY3A4FKpLmKyxyx/TN0KiUZFvxy4l4wO5NtSqfcmVhX
9IOQ8UcEd9+fEH+/vQ/0rJ0OpP4P89TFP4HcDluIKq9FyTQrXk671RzDL5XQqCAPOww3vXu4e2op
GqX4K+8TljMdqsYDdAM+ZNNsWxQA+EnzpTrmf4bF/12qzOVWbikyIl5UmbWLm4BodrzOstzAed9f
CCt2swYFoMENvx2DRlIfxGNtE02O7AHyVDMtkTRMlb9hTeA2mezyHdaIX8lp/u4k4hIiGcpp0Wu1
1w+rcxwtHnkXREidAn7/WXaZ6I92X2dEWTbM3EsI/g5xkTOh6y3iYVyPU3YB9J42gQyejXwHpzkJ
UBNwIAYW3yDrpRJmNMGlGWx2OH02V8SKL0Ra1GphjRyt6xq+XQ30HBUdoD5WiRTtlNaadRbUVXro
xFZxGujB8caVF+2diFQ2VPWQCV9PHd7SVmo2H/JUITRHocumnJN1QoWemSz7B+lH0o8ZjHHTETvW
C3V1WiX8zyKIk87uvd8eToBiG6KD5t+iOgudS0O3Qn8Vew4D00nyPr4CGJJ1ukwn/C1Zpy3jJAYP
B0KKqe+QB3ifC/fQeDET57xRP0jQM2PCX9LJZa6L3a1PCM1x9Y3XNX7/Pd/Qt3Yrl8aOJZbd0PKA
178299l7uoX0wLY3cM69n8/Z9bJJp8Pc98UvSi4mQKymliKVircbUQrcmtq3h0R4a62cYAal7fr0
jdxGqLpmq+ONVeNpwRU36COqBRVkybOGvESfOdVJLFgcJmju3glCjuodrlIreJ7kxdwDBIgCjupt
lkJf0CejgxcZobA38P8ZRiiDWrjIMOLqf4Uv9jryOvYsvP9tvVV155oZ/ORWFD32FLwPm4xXBISv
K24mufv3fMb+qIZN7CAAdOGwwJb5Wwec4B/O0XGYqyEuquGS/AAI1/UBkhPKO8AIRgDSAptiOFzz
Es9e0iuDhvPSifc49xuqgnVtWuK0Fwxypf45MYemFmctl+C3flSB2yD4gKiYoYv9PYGOrVnrmbho
lvce6cwC46cdzAaOlSBi2AuXoAnZg0none4VWtECW/eBtK8UyzaddKjESNK3/mTFd8fKVPBIL8Tx
O7vxDxym8ZuvSi1ysdaHpAkyg/IN7HdvcHofSHdLeTJkiLG1oqBOsVMOmqt4um7Z/BMSONA08/65
GHfw3oDDxpoI2NczxjQpWgPPJ57xTq4nD85Y3poc/ykjX4esOI5japCeofrOcuUxqdYna0yPvzcI
8SS6DSNqrud1dimI8TbrJt8HKIhFZQcADoaCkxRsVgQd0m+hwvNgSfPToVtcYvKg6G1PgNKJaOfV
MI1y+TVVhmuXIJyZ7VdJYBIxVh4FDJRJ+K80fvQdCMEysRtuOY4Y3Wmv7mwMhg1TVVp91NfqhOoB
lU1eZ3+w2hy8fA51+H9bUP5H4/fzUtx151SlPuVyNcbSZDIjuGVy5HitA9ZUMVOIth6hCaaY3SPU
mR9dK2slIJVN7VjwpMH2WKN1W//KhfnsVXnInd7G6NzpXVUuHbKGK8Qy7McCe8tBWF4Pt8rCB8zZ
tvuUKl1UI2rcDUmg7ATw4Tu7/piVaH8rU+XEwTt1DcW5moBHZm5M64H0txZYWUEkOaR4UXi6ZZj9
rDHkh/NNONDutvZJBy1sxecm7CcbUkKY65JGAg0vWiw4dt9njBWM52rjLCi6uEDZRomchLqtXqNo
c2RIl5nTlj+2wFGDnOHKMk/w7ZuUN+JW/ydVjdJ3/toeYi+FT3Ov5QXyZcGALjXq2unSwA4WOJTF
FSNm0e2fnazA49kP367019GWn+VX4dCnDpAVHrb7vo8AK2Gmqgc/5wrUXINWZtrOvxD47GZpnPM/
E9ayQv8NJsAjhD7eUccgE8j1quY0Z4ggEeskfs+WHdx4cdO8CQXjHCBa2lBIBOyq+xtxKSEfh8tR
UryJNP4PR2nVCcPto5mta3VYbPCvqFyo6RZMmzugDAwq29vkWjirQSNQ25Rkyn/o4LOMsD7n2hFG
df28GjkJTZv+zvQbAV9ZUqPi1HlPMV5Cdhg79zCZIZi2Yc9sN0EiYUYeOhr5ZTa5yqwzWQrKWVIf
w2FNC23WinIwT9xFlud/PobD4MR8PXocomSqLprtTH0NM51HEYTfz0ltqCJBvADdpLwIYvbwvq/k
bGJfoB8HTKhrrurCSGZvctOMKg1nrNrGmvJ7BNzR1UJpplLdQkX8IjTej0uhzdg+WmqlfcNAcnF2
u1BVVl14BKfr2N3xlkd/nf3tkT+Mbx7INy61LVIFdRPpIb9kh9ec0CysJTSV39Do+9/pKYzCrgHe
pW/cuDInm8uiXS6gJOwWFe+aZ1oUC/H6D4L6VjmO3fo/1heQPtBEC8LYrhWJDB/MRW+yh584gBLW
v2ChLCaRSmehhTm+o4NwiC5NvG3Ey2RZIQS67H/T8nADtt1t9QoyhCMnmXif2qHdnSe2jO3MF3vY
heMRC2kqDcm5bAc7U23FvryCMjnZQUP6wCHWp5fGgMpUpHl107cvBomdITpmPyIxIo9QbtVK5Hr7
YDPVGinqm5zDYRPvkqWWyyE7UZGsseuvuCkxJFuytvbelBRlJuDBRzkBpnhOOlL0J4H3V7B7bjHo
lz8i0iHA+GP4OjMN1CtbQc9oH6w3iZapRdk9uKZlf19lgCWLLO/nGGAawlmI48KNqqa/y4lSXkan
aQ+pzmiZe1LzxRQj/ULBz5NWPQm2n993MnPsExDBRnwMJ37yifTVI8tNBn13Or7opFhT/G2NgFX3
1eIUW7NbjcSF85GrBsprBYWnYHdGvlhtxewHe90/tHm6w0fcGzr/hFfR1O7FbQkSqkmCM0crrVab
QsWXMadH0tkgXSaTnHaB++Z/3kje5pM+Amdv/0xwrzqf6QO3MkkUSP9FbQ84IKdJzuS30iQZhhir
NwynLL5eSDBVi44KQODUtJ2UG4lx7EIUQw3x7oWJ28sjDC6Ze54oKVBymLdB+Sw65CZWzMsUK6hR
PKs/0l4DH2oJJC8KW8lIpj1rTpCzzs1kAAsdHwgzsGrNL1mK5+YpLnR615zuteSupTe0RpPgMRlH
el4gm8+pNY9br8KGMzacSs2g3iiRh61BcDzr1n7XqT5fWO/z2UyLW+RE4ZBLuwjyr0JYeywfmt0H
5B51+3NhXIsuD38nDLUtPcTSUGCh9C2DCga2efID3cI+RHbBJ06d473fGzNVXMsUBY6rBCxQe5DS
L727cfpzIgKj5L7ntVcHizEy+pb1HHSfor1iNT/IEl+FHilS61HbEOj9Pf35+frQeggYaifwClop
nfdLA27gEUUjQk5pbx4mAmZuSZSuxFEBCx+rYtjXyUiYcDiXu5ygUn16u6j+oUnJ3gb7b0MQxK+M
FzuIkybKuzlu3PxfYKtbPH5ulbD2uBSK23HaQTgBi5IzW8o+j6Wn8hQ3noKEedwEx6P2e8Zce0mU
OGzUeyPSKa51No1m1YT/YuHaq80NSN6GUcIlTMmbe8gWvN77WzMtVAqs1huXsFqyM3+5+09bB8eU
X5HttTuMMkvx8e6KLSMGgtCTpjuIx6yYKmw5TKOdirAQsivjL3PfRx9JqvgcS41pNXbnYvBbRZMl
rF3blvLKquQv/bNy/O/5Y9VRuxLL7+UkBXGyhub0xsFmQh+fgKn6LhMUY7v57bBFUMSDQ3yCBf5y
aTuqhzHkoJZlLJfLTnvgTfwhCDOzbd67/7vNSmp9dy2wkmcyySSmJlM23Pt+vBPrIhlWDUcueI5q
YKnChf4lUT0HW79khQj/IoyCHYbCxNTvYe7oy7d/T2nxSwOvMlO0LbJCUt6It+d21P95gwPj5s+z
1Kn5eHAQb1Hqvvc5BmAiwpWTgpz4nJjSnC8yiyyCiGsGI4bUwb483SW86GqTZLbE451STBcNleLP
WuuKx/z31w1jZDHh5xH3spOzIpSojJSLSVIVJyhgDc9nGfT3oqD4Dx2NXl7CcfNlmm+OI+IcmoIR
xtTszP0t0E0GSfrLODw5MZR7m3obMyK/jFp6I8qiDyFNmTyHsdbKjlUAH9FA+fBcYJcZS4kfbyw8
y/nQNsFEdKQ25fxMcfhTyz1+QQdiThjhN2ZtwnN4PiyyG7lV8n5exMkwI7pOAfS4I2fYan0XnPQH
Wu5KDZrX0aiA7um7GRqZbnp550cBjT3koDF9iq+Cbu/0jx9s3bjTp1ZbEfYRGuTnh0sa6Sc+QpFZ
G10s0xdtTuJMIQ13UkUJ2f7dAqK0/JNqKb66Di5GzBQ6/fLxKX3/QDHJHe4TpZS3RHutmqfjni00
fLocRtIj7d/6gHDwJ8TpimJpjh0YO4H0gKmKhgxVypDxQ8ibb08DNJEx1hzHMyYnmYI2z/bBypx+
YdXbyCXA8RjjJcDghGLYN8YkB6pxuUawg0fjAjEr2ii1juCyG081ZsaxL5LBn1GjWP7k8sdgRHzz
k0wytGpv25+9IPNjEQU09VScL1B9IOmIMoAbruq24ohpYYlw+LLjj+FWAtPtlQ88Q6dd6WPAjkc1
YG5vnhbG9G2w3wZKO+JpWByYsIDplXR8V4kRCS7uS3xkZQMOHvrIYt6OIJCRTSfACECDKqjWMSYg
pggepVhQzhV38h3qQ5hwZ4Stms9oW/inVxpGli2d41i7wheySFrCG7hlZsDQZ2bit3Hbwp7PwJ3V
Z65xeaxncytvezmmaDyDiXU/cuq3+Mye306IIjgpfBMxG6S9wmZ+umksL7wR27qRW9/JUDZ3QGjE
LeJzMmGHeIc9PHXRMhADFl4NYsPLMdG7QjUgoG9hvWh/2/yrovuBymKIyZ8Nn+BRZfngKhBAy1TG
/JbKxA61gg/cMEl3nsRUY3R8oE9WZuWry+rNDMlTwvWH3TdxI5oji6E3RAxFS+ofhDD4Hn9xOHBS
vUUrIzvol5aJW2hvgyZF8uv+yrrGOqt0HRlFyf250eGCA4yeHO45nim0pob3jfhVcyMBuhE/rlw/
+wvzwjqVzDwkU/wFzU8f9SGvzG0J+5AxsJ3F0SgYs3uE71Ke9AFgW5IJKZwRLjJ0xBsQGZnJegh4
SaYP9ZwbbfLukq1tjLh29Y5MwNYSLopt7DL5Ux/1f7w9cf7E7aww5OgtqGHP+gtggeRYwJ1FPpx2
F1prFeqU/9YaivmpH3nhRinZ4fPar4FBv49RVk6bjpF32LCXRSLJK/U9H1+qOT7DMa9WmHBHRjPn
jGN1xehKbFIro/FQ7ms7//XofXOI8S91gzco7Ca3Hnni6zv9Eymh6SboV6qrRb47M5e5afeYEi6g
XYs4o0Cs5D/hXwdxGiZsha2mlm3Ihjrp5X76ucHgYHbxwWn+IFasL8hql1OLR6r+D/Rd3bzH+rWU
upmWQgs6nZFT8Bp3FKJSLASCXBEvh0EfqSv0mSlYAdP70zxj2qhpkA1nmkh8etL1ogorwaQWqsPk
9JIzhIgE5j7lfTp2TiLM2qZ/wZ9jzkn79N2LSB6UjGu35WEfU55yOgiMTwh87gUnWXddBucS8/Il
YENERX6qQtYUO/n7OifbAWSDwg1DHKRN3wOE4udaxgpfXyNpGbHqtlj9f2rP1Unuhqj9zGPDD8WX
Mk7siAec3kzNXaCYRWYHgvELjlrVCeUPFes2Uuq1lgtJ0sQsI9+Jdbr+trqOadq16Hb9gHXHd4SB
+23Xhjgoj2e3HyuIVwyc5wRDOLULT8r3q3K/fiVhb/z3BYZx+YFYInQkAAvb3V/Vg8OAC6URGsuY
+kst8tQzwtwFsp4Jvi/Z1q2wWLzjG4YaspLZ/5X2AnJkkRgZqMBLcJ9pknqYLmpsvU7BtRI3+Rq2
tzCwXLQ2+hWFetaBKqbFOEQpxRFofjsFJzkmoZsjzzHQEymk6cYV12lHg+IoKqXASJi0bFpURBOc
CM/ipArxJlLtKvBifIKdaqGacuXhBEpoO8EUgJ89TnOv4D0Z+n6X2WQH6gCbUBTZvmuKAl9ws+ug
1TeFr/WD+tVTedW+SAJYWiUyZjs+d3JlMojvw68oWtEVfu5IoxBzUp+dunahxMqfdXnDYfruBguW
OyrqRJDJLU77qvEsW7Ym5NZjo6szgUO+FD7y225d64jtD1rKSc5fOQJGYRRkPwVteco8i5a5qTFH
YB4JSYJxnU3NBOtJNsqW8VAoAkJxgvtb/7k2tImL4YueHa34Rfxm+Y98QrLdimuo7m3NLr1J62cJ
bTg+JaLZKgflPvXnwcsXAzrQeSB6ryZuG/HhiCs+0pOEOH9z3GOyQrIzXs3rsxkgka0OiV04cRy3
IPPp6SvvY2v2x85Da/U1pSiMy4gT0fzhn2uui00FOta4fFQLmoAlaUxbqb4/HF702Hnp15mPuLQw
RwPdqtaUQuWv5pNJ94+NEPlU5BO2H8e5pPvVCEklDQIEM2HbBWqcGG+I/9y721eUrYGrz600xbqJ
w2tPCnORgPNBFlEPa2bkjwZA0kCgzsikpWGE/fO5wvp8rvznfbMts/KNdfL8Jdo9Ytgeu2dlR01i
/IgVO0JOWHYLOqpEvt/y0x4oPDj7u9KXgXfYgJxnLdkYVI2RDwhHqsrqqRpFi7sdVH2mpbGhfoWU
hCON8hVE9C8Bqguw2T8Ne1keqm2HspzP88ufsCLG4AaK1OFY/ioQZ2pVt/N+GcnI1cZQhZmw98oJ
amDT4G9HLPHApW6zJylgHs3/mO+mRzwDSHprT8/ehRyan9E9uTSARz3ZVBBj75Ysm/QdK5WmrMVR
UPjEN7fdnbPJJTFWM5LF6AbTMKJacJQrwqScZTWPU3p6HZ/pUsTyFWajYe2xRHBschrpcpLZzW9P
U6QTzaIwdDqxSC5tUc9W6s9tgqjqcGt8NaWU7PYab/b/77PS4AdBKhqzeVPt9eotz9W7zkaJiubW
cC8+EKxsNVT1e1nS2PZYp0jJw+Hd803G00oPC17AU3s16eObrw+kTzlUQsezw0MYItAF7h2jvT4X
y+AIiXttVYOzDRwol3cGAVvaXkTgi2YYYnfd/zg2P/xjNB1vQme2V3cdqijScKj+T/KwbJydnI8j
CQt8yIuTtXQNmK45GGvseRIo0/VcxqXIPNdb1EHPddj17YD8Hk2+nLxKkzt/iuCXScL6KybiaHGs
48UgwHEEdCsrVX8Owyw8agwVFTWOvg3/6/lRF+/Gwij17HpUDtkT/ddSwyh35SVBPMbpCvYQqwqi
0xc7lnihn3cRqAWVSDbKxXEukXei2PTvOiUJtgUEDyW9rAWP815bS15sm2IlaM0LBXQ9o0tKwSnd
73jG3IMlJzzN7UjL3+YqVAgCInQfETuxzfW4URal2Nd7vBbGXE+7Vqa1s7mdChBIa5dulsEzEccJ
SA3v7L3vRZqqPuxIFvgIqr/jfaw2TkCshiTcEb2f+4V+vMdVk+YK7QlqOT0mpJxQ/Ni+yb24Lbwg
Z4eLKoA5fF3rh82YttuFPkWawR6r+JyM+IOmJeXZPabuwGlZQ2hpdyqq0CvjP+O6sa+FV+D1a3+c
68UGZoRegSTPwijkK7DtS/xNJ7Usi/qAUWhg0lmqPT5x3MWwaolqf8fJjKsxRnU7CNGFPDG6m2zS
sV+9PuEpaZFeRtYfAGNXU3FjFyuqZPtqvx9j4Ul8MKZm/0Ae2QTfTWCEzNKH5SeFGDjMqVRGWzvK
y8Hy3xm9doYS8IowaSGMqUUGzKs9RL4+B71ZGlsRV3fULIatCljUwcMHpHL5QYJLNnM6m2j3tM8w
lENG7yVALMsCkc4EueKvrO+6PrPosERipMaB7+yTAGxVsvtqT/t50rbCnqISCeB3XxfGm6Vzmczz
0jToVykKUBmFejVU77WWUEZU5DS89xAK5p19oGcxOfr9gXUwbEQcKTwoMOzYYTxGq1m447FepI/O
iOZ/Wy90auGaU12Q6eF1CFz3eWvSSZqu5ChwamEbMgRtdjYlBiej1SJaG9eL9pmehFb+ROnnTKBp
jOu22CqcqDl0SvlIQyiTbNRfv1GAl+Ha3O8SjLsYfxrHDPhq0T0rB2w+YSY7ho84bMd7tFauviPy
6GKvFCZ5QPc2by7T7SwABhmFyAB5WG2o/vuDMfYWj+Jum3bOK0yonus5JVAufb0TnKyGv8CLw85/
M1UaVcynkWEaWlWjUQWCOHwN0aDxHhfXJgkimxDqvtavaRZc/ZIE7o/Z4exdqvrjusasWFI0G3ji
xLMMMOJAH2pQ2P2xYTTdRBVggIXYq5M9Mo7//UFqMUd/3FYJKM7z40PK/hxmYStciJLCUueF0WH/
Zct8Xoe4jsMqwTQxHmLh79qLNQgqJZeMCz/W94dtsR2WiVr8ZPKBK//44rW9Pf5ySWFOfKx43CM4
/rU5zyK9MQb5FQ+lGKxQrW/7q9P23TP8YaQTdhtMuc1jsPDvvPZxw13NGP76qnDDqvypVsadyVoO
TZ5GRvGH0FLHANZMNOm8x3VHsmwR2Qz7WlCSTtQsuGzkNT8dl1vMhnGNAKx4RvILZ+GxMWuHr7VC
zTfSDUBHtLt5vwIO68IowX1USXQXoyCm+DTcAyiCyav2ulP+dgs/WGtj4zem3v/TrtGl/98yeEtc
B3zoDsXapjhU0wL2pna/8KXpS1ruLOjOBNjPJQ8KABa9HehX4DndV6ARebZYGCXcv4DHqpicw5y0
hwwgxMqaoAkWswJGwxfcWZDxKqAGAcdpKn1+YWjqI73IZwDR/hCgA/MkglPkeO3XABNlRoRNKsXW
rugCOQ1JEKuimtoyfJgzndKAXnJkfHwQ/MM9pHRg/z3O41P0qx3wR7JzOpSWp+M0AxPPwD94UnJj
8w73FiHhWBrlft8oE2dspHPZqzjLHGco1s9Bp9B1OFLnNwRCjdVYMyqvdQvtSTcOJ+067Nsjs+DV
RA7X/0D4SDR3JzB08LKJSXuBSSqU81QCA44o2xINyrMQhIIeAzaHaXHSYf59MgjB9mz9W8tIV6Jl
2W+9NgSFciWtHN9cFYE6rH4WW8nxQA2FTzr3XCOOgiucas2ATxIFYi/19RFRMBVGxwaLq9JvLY9D
nMFW6MoFEgh0TIeXa80AgLARiPqzvCKyae4j6bQi9ye1ch+o6NvvUy+eXWgxveJ7wRuXj5g1eoq9
IbjEYLhnAKrLMqHtqaxvscCV+Xa7lWa4zl5V4UxDFxOgWRlBhve446DxrAZpP1Y8hvnDFeuRBvNg
/LMVefrkxk34I1/SPeS6nw+w1LYuYeUMspwfXDKL4kp0k4JYdb1wArtlF8Lgty2PXmC9d4gJPS7L
bPIQ9CFL1kWevaEuLRGqeZOf0RuAbE8MJ6OGD9foVQ+QkA5FEzW7gmKlcGAo1lMGOJ9sYdcCY7zD
EuutbAvzingjLhj6xNs7aRuuO1PY9e6U0wL6FvcYzv3uM+8GUNdAzqtn1C9nAkhSCzvBC+5lezcR
wM9i/OljIa9TtWj831IqK5HgZCxIvJAs8SJ9NQDwL607RF7y+pmpJaixEoYA1M08aiQpAMdA8SNK
HW2d0OQTUTMxCfikt0yTdvbr+ZxmYfFbcgqsUw3unEMOLzqYzqhaWLaT19nimahAZkDA6KBfAO/P
kX7w50HrPHw34bV8/6+73XsdhU2bOau0bDmAUyBJ0gp0N/7u0WshbAmVIMKPmMyA7w9VjDgxApcO
B90HkI7Y0aURJw+Sw2hiOv0xFGaKVrP+a1y+jAz4PJtkOk0tXQ0gHpcHq6X5lrHWy+loNXIQBkVJ
N6cNUGcfqqOBasRKScpfO18aVIjFJivIr4x3EvJreVScVZN832ILDYFGfKlMZMAYaxwzniRhMTPW
CFt/BlWdgO4WMdx4tUVD5f6TzaaGAGt1qRKbId7Q6S1PutrDOwWR9rkveex+aR+GmL86nl3K9W7F
7rhRxchu/poX+URUHuMH60k2vLpNzSe2758I2E+4RO2acYgyX+H0NH6XmE/g6eqqWLRhdgw/t66B
yJgQgHqMIDzt38DYgYryOgHxHEPBWhU2GOeEMPs+yOmaiuMYLqA/ve0SOKycZ1sXVxQX/8RyARiv
GBO5ahWwDWZbo1CYLZLnEFoZbs17TtreSKb/45b5rGz5AV1zgexGfWz3zrftbX23TxA6SljXsOKf
dS0dNiHZ0jtd9+xhdxput2ECHn1H6Uhe27Der6ApLME5V4y1UVJT9rgS5iNy5jnwaRrTGaSgf5T/
ouHwBHOZQwFXr+QKI37qS3mtFOexs+EAqnVSqvg/UJ9ReCSigW9485NK/r9oGcL4mV4//upL+sPD
/uq6nLJoXkmhA8APn2RBN3ZPlxmFdKkqzRECC0tHMrm3SrNSXKrlKvVMru+tycQam/BmXHFL17VA
/kRd1deRDG37RpydxOKG95yJSjFU9EOFuomrsvPFNkJ2JKTJFw6huiSyuF1h/6zwC/7pb7XKUbNg
2Ugyzin6mkdnt835t3PPFwrQee21Gt7oLriibHg9kvPPjUXhj71BswS8wNeKkfQcadSH1Vv2DkGe
/ueDpihxpXKiiJBqnjNMwf46FOIjt6EBA04iab9C2fsE1DIBnPaepEjF8LRPO3PHRLBKSubNWwBC
Xceg9epsvYDS5lPi/wLqH7jsHF+jhcYmU8DCxLzNGxEiBp6G70IuA2HRbBNqp/ZnTWkOvrsXdqht
bh/hfT/tmvLiEE41jjiEW+6bd6XEMf89IPpEJwqlFZcNbEJ5QA78YtIK9A6wko2VfzuQg85QPCyZ
csHINcjC5OJdPx9xxcU82btevCZqyzugOKrPZxWMEg8C6TNajjX6rzKuvP/kl20aLu9H2no6cyjw
fMcmrW88pi8bJa5rTC3htbB+n5GSkcnCozVrTqZ2gkXD8PgMONiJRBhmx+EVs2f8TcoygbVfX9BT
rg8/gl4vs/WP3Ik8tGH0nDfXSaP0A3DFoRofn11ACxMeDM175SE7yk4d46BSlrN0jVGRATWziktp
HakhwZeTO1yU33DJlTJ9i0Si79Istkx1ZF/h+uUWjBWmTOtLcK4jASEMuS/Icp44LQzI10oEbrOT
UlIY50sYY6H+ZUAG4tKPr5SbhO88Vb7/+quxHtIsNwGamHK7w3IB3n2wSe9SIF2zsVSp5e21iaHT
wbMNwGegfgfiYaBopf4a6frfM071lK4XEcnDbb+SmDRMd1Or8pWm8FRwAE5X+YNBRxX92uYaOwVX
jvGPdcDiwcmLsB4LCcmhMwxNEb4GFw85CNX1FbTeb4T0WsrEmJKI9YBfDTMfUTvG2O0GGEGrSLMJ
6AwK7F3fQ46pSY3XDWQ/FKlm6UfKZhJfSRmT1cygbg0mm6JflShAlEI6wqUE8eS02ZmM0Bv7EDQp
HWNF6jZ93ZxQB4w76MD7nPpA4lEdNOljXWI4I8bYXMRap0b/7DSRW+2vTvPPKh8JyiNr9aDBQkNB
/FQHrWJxV+/evxvZQ/ZALyWwLfi6lD+c+SOiFJFzHN6NPcpNglnmf2Srb4O8+GLORWntMo4V7MJk
k0UG6z8xEIL4dJ8/97FQJ4l4d07Y3rHqB165QyIxxJQkPkYtF8Jy6cwlPk0RspMYY8P/XPJBi9D4
IUptudx49ctF8ex2xpDplNF5ymOrHmGc3fwa86Ft7XL/zTKySBfCqyFDQkV8aQOufuljtPrOFFHI
qE1V3LghZfQ64e/a9XHDVZhoBL6nEllFVArnLzNJBNg7+Q8TGjCRcNvB6SbWKjcNIkuZX2bwjIcT
LWGAOZAb0cCf2XW8O1UNSC6DOH8WbKBjux+CBHWyAzk7FjlW8ksepvEi3GM6Py4S1/8LTshyd+El
R8R5lJY5VtDKpPWKl8Fvn5mCH9ydVj7fD9ol195uWCsgymFnqQrZvl9b9WUrtHAu+Y8Wu7ZVQBkv
130AM71ahkkb4lGQt8rkvf7/nNwqXHYthd9OLkZXEkY57DMnDYixzLO92r+M540jQEB1fnt51aGj
R/htlQ5bNAnSWUrfLQtTJzDZ3O1sZFn3ISBeo67w/jtKAkgkV3RYMvavaWAe3qBfQnWFIRnSjO+7
+RyB+qLP8lpt88XufdsnHmLISxXarnmHBpAlrN58vjkLsP6tP4KaF7U5cOLzOw5mEZwJouMYez0w
o86YUrcqqzLeomxVon0WCSu+Eow/GujjJ94ydHa4HUfT/sQhd+GjZ6DLfbaZaKQBLStyyhHPb4Dn
QaDfEMmZFF+B8mm2msiFdgXP0yFempQBBmbJzeHbSH2C3uSc5AWoYdnpyjmASmJnLd/5kkZC6xNf
CHxrSd8rkWAawSsFko8ziEIlPaFs5YVnsU14F2In+doM2RdAcSnw0J+XrGOHLSazgNPu+HS6HhU9
ocoQcwjSVwfH8XD+5bYok3xmY05cI4RJlJqT+1bSjvsW5utRRS5RcIk9lw4NTby4Zws+8PfOZPEH
QwhePchO8FTPGGX9BoGNLmMg/MqnI5s7I4+nhIeljSwB905MKnqMZVygZvnxXMa8SYNbGccsqeyL
tj/FAQgHZQ3PC5hur+rj+sb/68OV8Xxv3AXrkLK5pPhkDc8EjSQPrZVdo9128eJgGsuHhdS+QITZ
u6pPddjSX9PaXRvOUhv9689atYDjeGvcJ6d5aTJzncU9peTnN9g8+TXVxkg4bI3peadkRItgckqz
vy5tqnJdgj4TZND37yzATcinndi4HUnAN4ga41Yhpl+A0FeunRIilTAKFgwvDBIX1Wu+rMtev5LC
Gl1Utp471xEjwMbCNZjAFBKSU0v83Smxn1jIBnjnqDy122fqW6aWzvLVjqoqRiVxUnxx1RqwAn12
bR1OobjfRoyPjM+L6TnOw1nBXkltAZ7Da11gA4CEwmzH5E2SNL9RmZ2DgrGFhEM9NNrGD8yWcJfz
bACIwx0uNnLG2JEVMLAbbVZ7HCjTB88Sso3aFNmjiLDtyumJZLFwK9G9aKKopWg7vylT4mHvwaQ/
NePAfpdTQiI9wtEyokCeKCGJ4jHF6kMxL/2bDOhoavTemODn+rdlgW7bj4hk6023PtZoY/7+WutZ
Q16135Ee7KUyJopryi5kxgJc/CuKNA8PBTbdd0Dru9chR82aALUbehRyo5/1gDIHkfjpx0new2HM
LK63tEAjLbT+8Ng4D2f76ajx/Gfm9AejgTCHJwrViOP98bcz7heIlqOsROOjULw7BWGdiwwf3oNi
uX62fXYPypuGvOEwrNxp6GdnhrpULXsOHKjl1lkJMOy6Wy6VM2MyHjYJynrCbkqg63yF1zQNJiim
pBz2iz9qdam80rZWwV4cAzPtTgpZN9oODyUD5LvB+I1rvTHWwNWWRmOTY9kG9kibaJb3ZCmJX6EY
vf2fba1RwyF2c932cMzNIv8c+fe0m3OBMzgOHnxK5Tf9E41+h1xtA3pzyzY0+wKNrr5GyzkUNy2U
v2+cDtkS8GXqvt8seqQkOF3DrAIgyEXpWnRRqM+i2xzeJvJ/dNvLAM88+WmW6QdF/CmJvgWHKOYR
xvfuursYA1qJUiY+xmRUpdAZxDVR7mUUQgvSYFfaiHH4FAPQuC4uw/nWIUoFIkuQeHSuQ2MSXlqE
s47RdH166PyYnot92/jCu2efImvC3+weiEWZOi5JKM9/mEFbz4cjX7hM2RJdnxyFEC6nDoZlJQSp
dXsjSA3lySeZcFyGvtQtBWrVenOzrymnzCXRqXXRinVSCMqv1mibf7sz/VllY34ZV7npJU2rt21t
cq87O4ZYjiDcGverNZ4xD8ogHC4AxSdHLVhcx0LCkdtglQGZxBWpdH/rVGZ2P6mawmrVd+Bh1K5O
fIFGNtX7PC2Lh4KNyzqjBXhYtW7USiOSWUX3yj2ztT8OPxWW3K61PDr5d4hjfz+Nx/a5vaMThjbl
XTUvoOjLbn1GA7MA+LB/vm13AVKbGQoWdg0oGAz5jlLdiayFkiDLnzVRvlZuEtnWuLNeqxlKSjZ0
tRAFkfCimaNbS1gIbXOL97R+BbyImIdtalZ7Vq93X3KVwhJ6J4d6ieVRfW82267zqaOShoE4CdV3
Em+aFujzcuDdUH65rQw+RTY/w0l72MCR7WJsS3dnQnZbOJaCE/DtZ6WrjfNVnVcqJ/zeMGGsIEzd
fe+IwYLykf4YMUZdV5qJ9iaMkWu62Hnt9m1DdZimzi6XVIX7n8a/Es8dCIrZQK1y74gYtqNu1jDq
XKsHUBOPXesBjk6nyqB1vY/sOTb87FHYIyVYuBPom1EDWCvsiJGWvTVW8tEDHgQpyQF40izzCaty
O1WxS+3yroW8NQa349Fkf/VDqnAKOJnvCtSmuwaRk/3c2sscatRkdTNIYkDCxLScHHeU6hcucLcA
5QMxoPL1c7mW1jEwzpm8lGryMHmz+RiGnN13L/VeQ05a84Ks9quAD+ZTXGn4GOcwiGigfXPrNePI
qtsNjKgo2U8200mbFdSrrPnFPjU1ajMXO6WNODlf4hfWI7d63dDT+ic8yprSka1k6xIgqIP2q7Gj
YRWxFuIaH1PABo4G/eusfdGH82NG4BEtQpKutTRgSq5TxaEa7UsK+pkJweddGrN1J9LZ8/XGFqtr
e63jGs28cE16Kro1nm8EOYTGvFFXO4QLQxaSXuzB17+dqGbTgdLjAZGlnWOAv5SFUlwvgGqnNZVV
q+QclpmvbpVs21driAIc5ZEh5cF+0s7ciRXvOjtFatBEVt6D3JhsZf2HOApuTdYhPeFYVIhVO0gB
i5DGcw7767G/ZJxNWVtw3c1VExyo9t8J15Vsamjw4X80sO2pbdkrPA3Q+CINNJGDcaA45BSGnYAM
fo93zvHMuC2XyD2/WcjhFzi9673fCXpPLNMQCsk1DH1q7DDmNp3+g825iKpHT5ECZjfZuLI0DlVn
6R3E/IE1A1UMVf0aK0ljWvQEw613tQavd11e0SbZuCFOO30v7XtrrKaR2PdeJspyuaB76xunVQ6S
BunRdTsVTZ8EbCNCQ5X9ypzkfyYQYXzthfAu4Xnq1z2ya2j8+rY8k54NSEnd7pz5eBqB/k6HIIBk
SnTk7rVC9mDDse4IkeJHeF3zTItEtmoWacfCG08ksEEY74doA0CqQfHh97uQzBV+uawaTKHCSB/1
kq4UFoYe5xJp7Vak+47/mwbx62Xm1tcllp14of7G/CsTcwiA4W+9wXNcBng3sdOVnW44YlAcv3+D
UCvIKDAktDJMkqO9JDoP9dt/kz2mX7LZHeUMS/RvXHqr8JdmSf/Wt0E/CnwkyZQnR56Uj1JMmLZA
LpBLYnm3XSF6c8iLO7gpqn3RKvBtM1OQ/KfV4RgLpOnpJCy/isa/VlKgg644GDdpLw/zIX63sdka
DA0uaL0E0+9VfEHltTyVNc8HwAqE5x6b6DSnoXeX6BX4FF+XEl05w9MyvNh5hrKti/dzC/dFF/NW
ogvCodhIbKTCwTAABq+OSb7LOVoAKP1elqf2XXkeg6v98WoovdDYyQByUsixUxfvtQAd3Fpqrlvf
47SJdJHuyvuJy8+QNy+MemTdqgdnzeoczLVl5A9uBpgeORqhEW09/meMU0MsYLgMcuq9nbJySWWO
yGGM0FjImHvULDH7m0Nzc7RkrBQXEx4aY/agLeVxOWKCPLEKaoojR7+aBTK3RKV5AqqKSKeVPQuu
6ikka0nT4CK+DTx9jxWOCs6hO+zyKYzKq8MLKdt1iXuDnGVGZF3vEGpoC3jwrOUQnFSb38qDpCBp
Vir+mlehH1eUY0Ta7AitzIlhPtQyjOlWzWioeLCj08dt2DNmZXN/mSAAF9s/9eYahAaa7MJiNByj
/+fQiKtKVjsvsBlZG8FFBW+G2oJKN5HIWCf/WoCamKtQu4PPAOdtGJocmyQOjL8J1y+NzDP2i9xu
RL7g/hc2wd5w8SDnNHjVN4dzJRoUnrFK3S9Out7pPa+RGJG2D3ZoasCQbV/oUihuWZJh9cBhIghV
rL/cq+JbcZosn2qgwAFKzOnQmZDRjcgMPzJX0uWt3B0Nn+QaeQh34Av3M4ctlY7dZN6opzJL2Sjs
KRgW7ZF669W4zWmoMxeVIAEzKunNNbm8f4UNbvUv/2aNlbCFl2hzugUQPfqqnV1kr7LGJ/1X4jDP
54omWO2sMc/ecd8DoWwuQ2d3/zEHxVHo5eCJ4qAJlQ2jnoHC37rbxX6y2+Pomb6Dyz0s1fkgKqdy
wI83Yk1HWsVuJrHABNex/mkLQpo7pv3nOEQY5t8paZBSYjjM69TwJVA5KLg4Rl8iAFQugok8q1Tb
thVHqhgCI01RpEgTZuYS+7GMci8YTYD2TI9kb4a1Ry8uqWz137nveLSzWon53aK1jisTbZPvvwpU
s/H2+jXGuK+pnxY/QYEPGUonvN5EVDbf85Mpc+IQ1T1mvgyKbpflR95XxXurL9mWK0WoW7iaea0L
jgJm3vZW44xLT40Vi/Vu8MMdjlZxWkp0ocVV4jBmQNOyP65K59gwVbyHDYQV0DHjzMFDvXo50Fcl
/JUdssgkkstBeeIZCERKG0f1asoi18Ap8sbfswT3dmCPAk9k5v2YCJx9CtxRLcP/xIkmnxwhC/+C
WmEVgaSE8Yu2QiEH81dfTt/rh3NzBiQJVwVIXFlYZxBsG8ku8X6yoofd9bGu7JWlqBco7yoVLngb
SFyKZan3fQBpPkNJnpJ1+7voGCMLkz1QygIlvZHTkbM/YXzi53w/ab9ngkvv/sBGRPCQqy2YDLaB
mCJFotCxRMqE0jImn3r5bV/q6HhFdRKujxmPXAsa5urbwK91pxBQy2thfpCRttC5TJD4B4oDx904
5y3rqtYJmWTcTlNR98yqRxSoARDU4Clzz7osHk9OIGcBzNEOSZhCQcxsZ1xFqmfonEMmfCl6m4dP
KHjfSDYqbR3boZSUdZ6vAHL5v/UiA8J5wdDrG5VMgDeSw4EHUFkTdsaSJtJQq9MY7ebaoW2JKSIq
Ck6l8Yp82rDvJ24qxPAMP0r9wJ2nIYAoOQlrWT6dNNTbY5wsxOszGTMk65miVqxQxhNwMYRAGyT3
Q6/QTiivrc5TjWbaPdg5ihsl1TVZOCquHid16EF+7r3vmtZvMC+bKPU3ndYbtWo7U4jYqDczIi4W
UfQp4xvwOovZoYsRXp0jQPXOJ4i2z5pOK8r/1gDrbmmkCJnM/uWAwiwu8/w5NSteCL2tn5eB3h7F
ABBXXn7qk5WS3/20GFZJFBOcbSOX/ioAIpKuC6GccVFBZvj8Vb+AgiUee0mcl22p7Ek8OVMKagkk
Awg0oynnbpzlMY/6mPs9575w/Cxu1jQc5pK0IZrOsOU6DCHViDvVTIj+0OJqGc4qjsFX2rmwkMCu
80o2FdFzLu8k4Of0FtGi/h61juKP2e8IMLzhywxnY+KRbCmQvEmre//aOeSAADEw6QnoIdyRuSNz
1OW57kUfc9FfKoyDtN+Vlwu85IfNE/7A5qvJONtBWriQBSzRAAzxVSIM9VlhoylCbfaZcgiM9mJp
1HdGVDXszkDBXjpkozubr6BXgSJvv/qPIF6i8nuHPF01PGowJcLEj5uS9cLvtoeNbHlDJOwiYCsY
y1HXNKv+9RRdpCra7nGpLbyPsh12HVAtkGq88sED0VQwTMgDCeBqU5vxwvKvHtRce9qhWnC9IaAl
22lYDoiT9VPBp2LUA0f5OYTZg5oOrtMWnZ7nclWP8ROEJlUBkVMG75Yn/2BNShEYohzaR2qpniGB
ePl6dWTDgpSoBq7A+8LyEVFSEQPueOwbODYZypEIvqAHM7NnMx1Pzp3jW2Z/u7cmfsbRKQTi1gGB
v0lOj/haYt1qxLtZpDZ3xlvGcBKXydf9/1YpjMAMcMV7tmUsnB33FD4JAAvwH68HYPTxY89GI2SN
bg3vz49MRWp89JbFMLarIH58J+Zp3Ei5yjoeAi9og2sKhSN1Y9ZaKRJHZdxs1aJpy3xf86vn/5wL
PKlfqBTcGVbe931QyUc1wWzgZnD6N1ZKllPuDK1mp0PH9w1NLfbE4i5FeT8GT1JufySdZtEbJloA
NZ1HGMAokR23UjhzUQt+WEsqIs6EIcC29821lT/deDsFkwLvJ+vONAgyBLGyl98BZdTeM2uGZVsH
rm/Hx641XpY5F3tdRB5rPDnJCRTMDNLEBpO3tvs1YyiIicePtSNHNXumW6aiqj18IKi7agxZWjs5
Fes1tIoa39bCOm6d+46h4bnM1dTdWohXJE4KsPqqJkOAiCzog83YF4uv4QhSlFUmrUeXlf1OrKC3
wx3cidDk1wm+/ZzGHkYa9IWQ7pQMmBGR2JxZJ12YmPgWCsi8Am1aXro8/8XKssJ6sHvc4DBJFT46
wxBcaLQyxar2hianaFD7C3Er6+hJxzD1WV9jex8idODD++Tz6MjN+GzsjYNkqVEapX785jzs28OD
IdB4hRByJlsCVU83fnUsVBjnc4ue6HLi87/2U30qXnxZ1tXeEte8wt5qXzXbAoBaAkRd12CCBLch
Ufc3ukMwa5PgD+w0ekzDUiRMzNq7D6VhexbpmuGikCqghz10Lkqw3UlxhQ7ZCAB+ne0pCHFstwef
5pPz0iQXxog+o5rmv8cbHEy6VjaYfN62fB6nkvQHmtiLzxJTJ0icwNaQ79fekqsyB4r+STq3xRnJ
QK6F4kr5g9MCxf1oYncJ7MqonKz0s33oTBZOya3dO72XpLT65pgVBO5naEhEQNyDvuuxkg/dcLMH
xdezUP5RcWXLC/00Vh8bcsh3RPbng55ZYvA27r54e97fOxG6/W4Y1HUtLe+PEPDTIRUEodtFISkz
oSFWNe2IbMsQKVQJdQ6U+GTPN1L/oimxx/PCu+HxIaMReD9l9dJgTtyQpPYBRIcu6K87aPgrerCi
fibtExpak5zeWWYIdkyXyynNLP96sUpCrACJxtjNuIRKzX74eIxNr5M2vdCeuXglrUxAoQ8T0TyE
zZrK0RiUH3Oe3S7nmSdiWLSiXreE9SCpACIbJGq6gGlRQlIS3GLk8gTbX8m0oYs2smHNx8QjmoLx
PTWHZjqwbQ32+pl5TSrnjgCpI4jtsUyOoScebF1SpP05M2msEYqKegjob2SbD0fv1xnJO8hMUmA+
O5vnBWIq3dwh2ytHj8RsP2tz5NRSFS3nPxOXhjI1Uu6hMnoXl4XGI3rjXkXnlF5NBFf1xGRP7aZr
q/XNwBuBVEThsJ7AluEm0AcLKCCmw4eB5/IKzEEEH7ArrGBkUhybfYRlLxBpvVsrO4VGqfGGjzfK
Wor3G3mOHRFcjyqeJhNEkWVPK9x/9JFStEZwn46XV8nYFgKIrf1gGaOTMPoUu77MCUUHZyNPorGH
+/gqCAQjAJe5NjawrHBZC0r51htRAO1/kqN4twZ9qP10gJdgLkd+d2RrGdiY7wg1XvjMej9ytKTb
q7bzNpkR9Fxs6szNyuKkOj9/eddFUDIGBPkGL3i21dELd+jSTZ8fmjJkxdoA87v4IbHW9olIKZCe
7DYRzrTN346XqPWzKwJUdj5nUKVdLzz3RsprmpGnn3+kNb8lQIa7IznxhpB3EkeT8hFvKd7wO4BQ
HWIKmel1762DH18ejgbf8c8PQTpTb039qlbQJ5QzKfHPn41aZje/mQxTkb0KvBtghRpaRjAI8QM3
odIoWqRjllQxiNwsZbYMZulEPKdJta0ip1wF75pIUGeomwDBh3UnbNHvF54BRRyzMvmri3QzqTGv
4048b8zm+CXBQM3myB8ikL4Ghy/fpfuu5rGmp3ZEPNVOfvG8+Qz15Lxja6A/NcqPRQERSDkYQ3Mu
Xy8ySDNjj+TFJMXK3QjkCEb6ABAw6LYNYeLQC9Pl63XIceqpxo1YVxsA505lLlMbpDIge6JM6cmk
9bfdSld/tXMWl0/uy8q/0OwUh8BYFPMRlabTNtSpJXWLaOOhRj+xoXXmSgW1sd6m4Zap5tMYHqWi
XwF+DxDF+hM/XYGnJ6SKvm3ICTtPGnf/9AFEzAPZ7BbNETbku1QwLZAchloMaAH4OxkrjukXKVBH
HLNfJklqy+i5RHvDwcJXNyOYaqKjogbP6F8SOjJbX3ZoQceSmGjUOcMvtQBkNEu4X7Zlvz6D1p1c
VYR40oF0FXFJBfBRKdWuiqBdByDbq7h+aSboKLZzSrimWMZaPatmnV+MWFLTkYOFjuEAefbV9PkT
q+rFWCQX+FkhC8O9qVmqrtgeKTAJ+wK1uhlF68XGqih+4Pkd31nsRTUC5wXgA7n/wz1Ey8E2tdKF
tVOVRNlzT5OttppF0HFfmZUI2vXtjD1dUvoeR1JSQnltDuSzyWfwjw2ECw2dSKJXLGHz1Yk6tqYa
LghOkdbyYPOoYXVSb0NXbHxfr19Zz7v89bsbdZNupM2qyTNRh9M6RnJAP4kuB9Y1YFr/OxEYXP5K
MOTdu9ShzPaHhXGHXr5Ly+y2bCNIGa7AFg5MKm0AJx4tGIg6SXnbBgFete2nOPhUAvrwnj7Tey9i
FdqlLYWmyplLc5m5F6bAoZW0ix1Ql8+xik/f//P0oHiDZSJEKnQEpzZxDC+nhO28MLbGe0KKVItv
/oHObYb6xE29U8quadMJTRk5LQYVYoOt9ywyBj8wWx/qPu3N7Bt7ebVNUtjsr/zXj3j7OUSBhkLW
Qa7jLrYLJYlB2rMzWiJatazZQCYPh/cCNIkkB4j0HZyrGef/CaJRPpdWQdK3vCuOGfogc00gTKey
riZt/FaBzyptK/O0WB1BF7V5ZYO9UwhslzXgSrO2nDHk4hSKEMH1j8CZ9WddhenyRv/T5Jea1lqZ
AYEqYyzwarVsHKMTNgSVdLzM+45h4qP+YIaQSIX9yxjXPfiUYbnNvHlJbX4KS+xTNVp8vfjynAsH
2JkU0BsK2qTozEFVJyygMcW/donBTIpCRSLZGw0Yv88fJGFd125YxtBiUV3Q7PY+8oyQHqe9jA5E
Z7kFXYgqpIW+PXQBWKma1qUP/C3JvD88WRxRkFDisfqXhkTFh3c3q4PGYtmi75AJkHZfJWT4KRmA
e6B1giUpHMGdnieQwjhnNquad2D5jsq+LbevvML/d6ryW7aSbLxoGonsliJdFDfL0hhj78TUWrTE
V83fND8fs53HHVp/MhaFaxR0SMGofT/A4J/KakJBgLloGANiGc32ON9GELF/1HbsAaVLTLsKAekd
Mhl12T27NZgP/yLOoZ/1MEoZWZVDTKUzh8U8S9YSd355RxiW+vLVkTkTgmvfj6EZFk6ZDCuX7Vm0
Z8El2j/suH6xjUbK8BoIFDVhKKTL1T83z4+sxnoyJFrMTM1LiqHGnXXp8yLQsFnIUoe6nds3o0fo
3T6DP5tQYAhg3okwMMJE/R7Q0ZG3ozHc5xqzmbKZIY51u2XZyz+lvMtKe/Otk0hlP5yGY56waksb
+ao2VR9Ge3iVoVCh4WpH+yi1UaQccclaM4yxbZADPzhSycTmB7+AhOr/2haadzXOD+WmpDH85Elc
A8I9kSapHqyO68c1c7KJCmzQ1N1EFkaqo7ywWlc7K4gMX1CcqcRyFsaRCRge2FyLijW9Tt6lr/z8
5k/uKVSLV3va1d9nl1DZK6nQMjYgdXuCS75Gz2Uk22F7RzZaxjRGyrMVv82Hc5Ha/C/u8kwRQrhE
gg6DQx9HJnlGsMmRheIB9JCqq9l2PWbftAYotUgVs/uc6IdIsEivSqpcZS3k9jMpjUTTMtKmUI9s
ncVYqDZWTEdgrHtvyN3jEFBxt56Iud3dMAD0eIvF03ZGDD5f008QhT3wxsOOWPVx8YTBhNPbljvW
/iUaiG/h+GutObpb9dw9H/IXqGPjUCeTCQCIQ/UXqcC5+Ik0f9+FXDwbn73+CEbcrFtSjEY21OYb
7Rhn9PX4hImy0rCmj33mimpmFXpe5DE5aosyTXQ5PilZZtJlvf7lzYsxTScbPLyaIHX8ts85Lm80
i/K0kwqxBAGY9uEdyvlBWGxuICKcR/c/e8FeMsnqTHNUztKgHhIVy7QBs0TIMs+5jW8Phf1w9ERO
894Db4fUTTfp7wvNFaSplyyh3xP5Pji5F74MHBYHJUid7nKnByloMbJrh8uZWCnBl2H1gbELeiGD
cCG0GdlN+5hQyZFbBVgbIOXHFUVtLDqgw0iIZPf1RSqo1PnolL64F8P4tr2nTcMnsfrkWGqiuBAd
rwFG+SluLiedaMNzY4ISngTi3+yLyLFnzdIiM1Vmg4dqegfcfu4CCyDNkV3CNwyz6mra6MCYGEbX
qzYzdCxbMPq3YnTLRPswvmYyJBtDfmGsRLFfBoJl3gpW2ogCVBwEgqUlkqLiwKUw+loBrXdBJhaA
VrHJz+jxBHoa32OswX1KIOe9BTpfGLBlR+SJaLYaZm+PqAGoNk56UWC5nAKci0zpd0GgxB/Iedlh
diog4l1ylZ/gbawpTjfw4V53pT4aRjN/cZN55WwQitrV1CB92Ffqk38apqRfpYO+6GL9YBvCIz+Q
Wv+xw0Miaun/yMVtyakI99tOl38jd3YbMH3ScmMe99Lb0dw6ocHd88sTHA2SLck1y9eUXymO8LcU
MMNTWaUDc5uMhcC3iAMhwGW5h69SyAZJv4Zdde7aYE0EYItNUZooEH9TJDMNJtzGwBcZkAcGrUqC
+TSvRHm17xKYh4hWzcmbm567cbSJuBg8eEZR+1y8fwtcz5rilkY6z/uHyDrwU2oe1GtYd9A8sj5B
9IM1+tPixpkMFbt2lyk8fP/1XaGoJA0Qr87BFftnZzJfD6aBonxL/MMFp080kcy6keycedv5E1Hf
qF5xgtd1cSbSmw4pD/osNfGxQd4zpv54jsuAzYGIrjESiwIKM3klcr4m3DbmNRIBMNEeEUelZ/HQ
TZiYX2saA4Ewd8iLTEndgAiL4xMNnMCBxpRXVXIgkWO9172IKDuvM7H+BHJxcfOtqH2WSkAMs6oi
8H+S5Ypd+AJ3LrQd1ZeJRdYZ+upbnJTFaAg0iSONz59Nrx5FTTlrNiijoq7meTW6bdftF2wj7OyT
wnSLQ4PsZlU2mr1Izj2oqhTGLMei0SUX+JjR5SKia98IvzriOo8inTyUq6kg+gsRkgsO0LtKpXar
QRLEAmPFSEgZCt8pHEDSEANHuCZvuScYrN07DeplYu5nBqs6q0eiWwS9k2cxCq7Yx3gMn5v1+GmN
L4wcZIVx3O+d/1rtVoVcq6us7LhaP3gXkrFp0Z//annM0hI+0+fIdmShSKZgo6e8r3WGlJTIB8yd
a87SDhkmGTmZTnGM5u/fZY0M2eopVsQAXzbe0NkaaQVjAbZXoW0suq7p/oUm3cO6oKUmUq8kZcbn
JFUaYcaAQS0Uivk2Znqcexl40xZ4TtTtcw5LbOGog6hrrz1CVxtEZHtH4SMGFxLAgbvvKKn5UHD/
fmCctV6qgdIYvSjVmNbqRkx6iaOASdJCzbkF2FtLaFkPk/tuSOhINYz9U5JHu6YkWiL9vqK5EzG0
xZJe0mpon4xVI4PIX2xNTsPT/G4k9doMJI+/IcIuNlrVpVnU/gqW0TM8SOtfxIEOKhEgabPJgMj2
b9mGL80ykctd6AkHzB6LH9GWS2qWNWNy81zFiDu8uRsJdLDJiTX+0fYhQXJv8o75aLTKgvjw/fos
HldrbxLFSIWtslnCdBU+qdrBcfwjX751DU/2v1+4xnwjwro3+OGbcOTNu1kRNMzkCEQdDaIXvdDN
DKDiBf89zkwCt1dI8dtntxO8EuemQv25/++IjYSKdNnlwjIMquALA518LftwIba4OpGeHsVwvVRm
gkxnOpdwP3SATcNz192TAJff3tEapjtu4eZdtcjCMcEQdK36++PxEbeSbDFccfgcLWr1OnvjavEH
9eAOwL8iJuhJHZNBAcJiF5zZ/GJWew0kmeNFBE1DNPmr9WUltCUvXI8JPXz1vQmrzdSaIa/DM8MD
FQzhHDCXnSpEaaW69WRlwUqB9R54clUx6SKox6ASjCTo4KiP0ismmTl8u6LtTbzAeu5djK5LyqPg
vB0Gp6fzoskNQ8KQtBqvoPh8Rqt7L1xJ9e84taW/M72xDT86Y3BqvXfc3Kv/2U1K9foz0k7oWDlO
7apbEN6tyM//KcwWlRQpLnGHD9gjozBt6thjQjZAXj9YOE+a8Vz7Jk9D2r6ntf0Ehl1I2EH+YOBw
K30O1/r9gAnVmq7RTY3gZvL73ZrNfzTzM7/xOyKsndScZ5pvDRXEOBAGr5r7krxffNnYclE+TjKp
PzBXcghhsJrMXUohhH026IU/XbcMiylAocnBkhH7wrbG0IR79f3Tvlh92nTWM/NvjfyExXigAaEE
A1Y9ReXIke7M+MjmANtnJImfJeGbtb0YtM3xcEmzx2LupyTpJHtR/XPo38IAcchgP7iwDpqwPN+2
drALJ/AutAtFtnCB2zrROxxZ/QDFLJN1NXv7NBZaxdJ0OymbQ7aWt+wAzo/2xBI95ocFWdVrklvE
uk1U+1GXExfseJQQS/DZl9gpVO0BKocfEG8v8esaoCeAVIwkVBsht2voWbjNUQPTxeb/nETnr8LJ
dkiautIbYD/Fuq7U26R2MIrBh6evpXPLXY9C9MQky7vZIVVYAmYapl4yHCeVEfLh+ZKIg70+a7eS
+quWyBoxDZc1cM2Lm22v5nZLaeUmukqMRjBgSejlZAhBHXQOGy54Mzqz21Xv/H9yLpUwJwd/E5pU
l6IXnCaJkwyIRy2LJ7JtSecJ6Pw+w4VUEY8AHhVoZfRy20tw0UJ/4lIbOfOlTVhQjKgIXv7p06G7
0kbrWBjURyySwOaYk9y/aWy+RhpdPuMeuvUNRj7zJze71XcwvISd+PY4JuonAyn2qwcS2mp0qlqZ
YGgR2h9wTyCnnb8C2hpuUdJGFWHYHiqpPN7K5e/uV9bo8pJbfIVpHsBt3M5XWrmteFbdrYX0tsiY
6wwx5p7B2PFy7uff6AYoPL9l28JjvG0Ub0l9MMksPqGgK9pJTuU/fPJ2SB5rUa1+QhTROwUhOUrO
drk7Se9SOcScJvbu5lgosntCwjgB8MHVUGoskCje3/NKYCbqtEO6N5zrZukRsnPyqQVJheoYUSFP
NJzQ5g8U4DwU+zDjpZwp3BaE1QJXPMlyYpHpCQqTwbPerDwU8hi52GDHNmdZHFD7Zn4RCms9PjSp
G88Jzgnz6co9Or+ViccghFjQh/YIhFuk2HxzOeLSwBTNFaXBrdQ1UPmTiMp8GsozIB0g0LBZJz0Q
W685DD0LFLXiGrorYKzH/eRQB57xfmE5QmH3F4W0HZxT5d+WYebxyvFOW6/cAyRgtmlpLIVDRtub
g5LJvXF0NruVRDhXPETlFkJpYTqzmg3cFYCWi4DhjNXPugSZUI1aftmuZ9i+AOcwYMRuKSTGR1tQ
oXfICJLHrwldCHAsRofrESXCD9+p5RSsa7f5IttlOip/5toW6A/nN4zJadgpg03qXtpf3QmccVYJ
dJFKDpf72kqH7gGP1xaZtYebXPiTQt9Y31pJlrjYEkLLY6Pz6La83q3lhTmwpmmSkWyJOaLk4gUL
UeOlhRXm/AFps95M3YEYScJrrzfc2O4akXcQObIjJF9eMHx5tjLVv4UJqdT7q9F0amdD4bTaSRS3
cyeszWxch0cLcObGy1+hCxrvEx21h+HJkIadHeGR6YB9h+SCOIYJh5u7W2+I+xc7hP1U9C3hpOur
IYWampBln3YoEA8B0ns1pLHowtPBsXZ++jwY3bcMsDkplZuZooXHNO9X8MJFOxfO8TO6RdehW5W6
tvZhnwqKYLtaOuYnSELlDiBIR4dKExO5TUWV0wnEntCSQ+FrljJpF8P+Go6xC89a/4r0Rltx8jmq
Mk05EO5bF9ox4ghH24hqPKANq8p6VMEnrfIfFPw8DHbDSiW6qguaJcyLJKuqwwYgMpdJ8fTyDU7d
y7aEaHy84QOfzoCrKwmHfhr5eILul2toZfRp6a8LuD8RAptLTAf4B0ixHEFKH6ynaFbhcFwPvAvt
DalVXynzIvuYMWthi+5C3CyVdzyfNFOo8o9mId7wYmmwD6WuDQelAezqadHsWNITnXVvTVFgYX50
ziICsrUWJWsVcpAs0L2sVOZ+fQryttZyN5nOiBbM+KNi46l+4MGqhHRp6vf+vKQOmJbqF0wiiH30
YW360qtH9Rd0fKjegdR74XrWw1po43CFwOiWYNf9UCVdHyskJZr8lKggoRgcrcV8aw/yUMIBF4/K
lxVrKWdLQiF9cBTbi8d9INQKM1AnCPpobEtCqiLd13ugeWwGW60ZJYzRv4LjhqDlJ3bEbG/sdtu8
fvkl+UZa8BH8fZSFofkniOzM511zeXbf3neMQlKPX8zBAPjKkWAl30tQIVJvJWMeagmT8UyXGjdP
lCwSN1EfN8NLlj6c+XHPxSto7VkFNAGtE3A1EsdsKxu01If8AFeuXGvjxgaJ5QE70RnsbyR7spAg
TIBjj7h2n298GMY2nlOVV5+k9+kH5jBX7J+mWjhTFY3+rfI0Pslk7C1S5qWb8eoN5VmJ8XwBKe6v
dfzawHALwhRFk/SJtGVSrf0I3xIX4cxmTQL3mbav5R+DPQGk2dTAzxz8WqQ8jguUeQFdJBuI/XDi
HnrcwxbQ8onRnHAyB3n/YkIWEtI+Kzj9m50fTsa8jJBC+AULyLhbtlOR0LV6qOctJ2IroMUDlT//
j1GU9MKtdEGVw2qG6cfM/r8RlbCM0NrudQ+LS9gcvr3NjCQ3FT+y8L1eCp+aLAdye4gnO+mJZgv6
wafsDWorTGHwVX43/XnOMQ9lliYF3P2Q6iMC10tiALO5+C+rved5KQr5J1XvgAZEvg4TUfF2ukyu
HKYNkkQDmG655MVL1LwhdcNuSnuOfeWkMJgxszagk8hXDJ1uuT1Z379nEYboL9kX4/q0Dd361oIX
/swU/YYdUXetOgCg9hkZNSirx2G7mkor2m8qg9JIo/iGIsySEnJhy3gfkIdXkAWjx69JRInyeB7m
mYTxet92y2pxqXfvzrM252+qeN9H+FaPpvQGkvYk+bpe9xnsOQbxym/+hhsDy+rFabijzauJOPXb
1Yk8WVUbEwC+nI0WmGoDpf/Ua839Vs27MBnQcKTfDm9YVFvXWIp0yVVV7FpOGVcKRvvj6324neYG
/ysqSZg7Rhncjr14GL6EUfV4cmb/CY9b3B56QSQ4FGAQvjHE2AJf/TMcDHEd/TfOiRnMLb0QoUpm
viLzGoc3k2FvX+HIZzBPWSu93fe2OjOnUxv/34bm2pU7bi8tg3/LS35+GYOf2wbfG7VUs4z0o289
bbxHy5Lp3wYtCI5N6IBIMkz+VeTJWzzEXledqMSCIrkPhZRYr4OZdx/Z/uJPYKQiQRvZXXhn0AOu
deDNX05JYAXMwkN7/bkb43Z1M67SHQxTJdEN/6IDBW7DqOhpgLHiENqwNZQIMowcBTiyxoE1PSib
DnVCaVHwB7OvCEBGSN2Fce7+EHERCeKsHsjjSQsfOpjMpsWqbd98I2NGag1PUb+L7DqOzB23bEuh
9lSM67qXy4knHRJjUbJyJv2GHRxINagzIPJkk3xSPQGr0IzcACT3xRAMzSUhAdIt8ddMBT8jQYK1
1fzNL+WHKqciFnbewfvBbc3YE5Or3n0me5NqNjhkyDlDGrbaSvJ04wA7A/hwTJlcszHPd0hEzJnz
5uloLGf+4ZAnpfQniUkITZA7Iu1cH/ayzlqvKh2e5xbrhMxIilKn1Bm3LzgdcSUuo6DPNFaeWCRn
1Kn9dK7BZPXBMbB2RpkIvWl9Epn9Mb2KTy2rKoxmV6kGhrnAcOnYlhJ0KYh15tyRO2ewnS/X08Bd
tp/QrlSkX1vv4xlpUriPgCtqrLtLOdF6Mw/1EaTMZVQQqJrRK5l1fPTsIN+L3Ttokmf6LyOmJR5b
7HjNHFqxpR61RcMoNa+qhv7XCQhI6trtaeR73Kx5nkuI5Knup8TD1J+pe/LHLlNm96Tn5Dn0uFQ/
NCwvM/RyR0LS3isa5d5TRGns1hPv/QBf8nnyP8sigXO9PstCEM80N+uWImY5Ngf/45qUGBaFZ8G0
lCJhYhACLRyILAC9GMF90AeYDL4ZClI38OnPdbJW0VWcVdjSQMvbHLHpHmaspIFd26GRuj9Xy/dR
ULZtSt7+Db3RncTm+44KBOgAhpx662rNqJ8caKY1D2U7lNfNumeGVveODxTb4iLE1r+AOGrzqZnt
Nqhqz6iC5wT4MdmotXulhZOCMTqoB9UyixHkNaEQ4BXMY13Hm6u/mhQ5pDvfz0qHV+SmGeV0q7fc
ZmxRSVMtLq/0LD0qOwuuqrOrOB+yzpBJaOzKAMv67IC57qT4CeFBPOV7EpJnU2HFnmAzWemmTqNs
GDh7fXSgz44iJ2ghu8azCrY0e7f1E/tDFuENPnT/YaLI58Z53BERjcycXjCtuIIUd+nVDzY+mnoJ
jfq4wd7ALhOvuo3unBXuB7KLHa5EKYzkjBBfeOzq8FQjM7qL4p2yL5KM44Ecwdu1g4Sq5k0pfG7Z
j3Sm4Rwl5EZMixU+vMaRLpCJcPuogKFoeHxnuTq8rQGPNQ1T5PyDAtR4mPPaG9mrdTQz9NVDSKkd
rYTSxU68SkX3hRHKzoieU3R/HkQlzdoGrLSKc0eJ95/8qZize5ZOoFlya2iGAoKZAIHCjfbVbBtM
FDk14AC7ufOuL0MCYuCg20QThgABEanbanP0Kg0BFGwvh5o5ubXvUomMFH4nPxOvxusJGG7Hl3x6
dZ+XsYmaGGIT/pdi7HbXcA/zc6/dcd6/2c2mqYZcPBjf19D/qUs/ZLhikFDRtmQd3a0QXjfFJWEp
IDB/jL5mpiNvQzkhUrBhY4lgg0AFPglBa8IqbFTiZ6dqx7TIa+DpKja1GLyTlQwwL9F9YWKH7DDl
wOBNb8t12BGBOpfWWSer15A1McjIPSRmQJi4D6AWj0kARviH2dZJbV6tqjCh6EDgxA+rddbfaBwj
JnudjsrTjr8bAWSSq0Yot0xi9KHFT6mgqq+dOACYIFSr/VWbk9ZZ2a8JGkULGg7fp1FXwdBm98yl
xsYjHnthCVM1o5NWFE5oI7tvl7q29tlvYMEsAvFDhIO16D014H/hLbHhpYGJeRpOFpzqmNE9G+VS
E1K27S6Ewk4tNoqJLgLyAiWkwr4+rWg8mYlkj9of1gx7MwwIEhgDNsJ8YR/w0/muQtq8xTKtXqW5
0EAJ43F++Q3cNvMMR6KwL8YO8OK9+awy/ZwPgYSFuJr9eoT7DUnioYVRp3721EZ9u/Rf7N8QGONh
IR28f2HZbans1BTcpcIAPuvlosnMxEh9EDKA8i7VefWkYqhKTzLkPD+fHmBzm8xbHXfj8mHNXkiL
HAu9ye6GsTGTfZtKi89s5UYuHHkwKMrrnVQAXaD5Bp2uBsu3zB08wkQQusvaCWrQcfYFlIwMsSio
cQGDT/tSyYWpm3/BgUA+GTe4AZkocTwPNflWSam0fFc3oyvH8vC+2pWleG9lCAf2IB8Nh2qOgE7Q
FciWObRtJ+Sgv4Ol1+0EtmvcwPu2S2TjUYHXJMUGmP+pJH3VZHdZ56ctznUzQxVlMSH4MpBMvvqg
zjJUDIdJ0CTGh0zDDMjVhJ8pctCIcnVbHw5UlW5brM0JtnlP1GwC4mUzzAGkDOumnHK4tN/6lOLv
Gt9jc8QxCaqpMlass8xHvlEWdyOcNQmO8LomvyZfRDBt8HjrJezi0AGaiMyRi78egBaIK5kbrv4J
5nmOlC6FV8DUEdm7nL1PnqJ8aWqn7YYNugxbLzS35Jhpk7vXthyLz6BNOx7Wxx6vcYrLHestKgPf
J5c0dGRbAa9tVzr/XtJsXrO/0FKZ9XEYG5oWVJ/urF7Viay9ADyd6PNXBbwnVYlsGemtvkmuGBny
amP/pceZ1KxAG1fjpZg/vsvuTejSwQYMHGk7Vdy97caeir1YKRcDJ3581GZ7wNoxYJOly5G12pnd
eYk5uV5B6x2Yt8YtJf/VElB2AHka88bjEZqYZxwn+YvpH6MyYCPDhWvBnjncaN72+TRiTdbiXx2B
oYZs76R+uvhcuN4D4uxIC51k6QYrYeXwpD95JPLgQMHxoRUdDo1rNVyuWQJAAgZ34SWMmdutKI/F
kNDLOcRHlFKJCDBlwtvwfIfaMR8FRyUDRkCEiB7VBGyhaS/EJ6xQuq1a+in6GomaaRNmu4kWhNGO
ntcj/jMALLXt3wrnGIvEeuK70QX05jltCzwu6HMySwhlz/1iTdWoyx1OHBLUkI+nQmGfG00wQGBY
ZSpU9PIUIdvxq00z4WwVN8SB/dkY180T+8Ol1tk4LM3f2qvVWTxqcqbmcJnEOhUKvbcMboKMdbFh
plU55zqyII2UO8k8Ob7jdf2PB5uyoqWqWdgTp4UqgXCnZfzo30xU8AsmThlyWySxZURDlK2uWNjZ
BNyrFu/BbmSTduQa/ASfZPX1gXbv1WYFZ14Wi1WeR13/eeWtzHWVCiyA3HsNOjbzdo2lykQNNZCG
EVVDaDrBa3eq+1gjLkhqibfq5iTENXh8G5jrxR/7bm5ZMW5bIgtO7LU+NWHYaGFkreAbJfyOLYCG
SDTslBrL+u34ExIvjRkzpcdv4Bzs97MaDcVTLpDWAbWxXsUmkwmfB7R7y4M6EngzJB6viWACqk0r
SwZs7gHSOHhCLIMLRuNb8PQiGCHc+3s+cypkLvLOe6ucy6WufCKRTh9x2v0lyJYgGObmYLLIDPPF
KY+KUGB/lAr8zC/OqZqAwE53MdMQocEbK33FI9GFXj7Is800eCf5WhYrIEGlcpyR63wV8hBE7Tt7
Fi+XuvWe1mu5eUxrS+gCgACod4XQOScytcTu4bk/wGByD7GN9wmdxNuiBl89+5KcRtPp8qJ50iIt
IJfyodh12sfpV5foZ/4d+AhoUvkHw7c4+oeyeDyD9JhChvaQ7UvaF477FcBNZHVCk4F1RkLC6WRw
QvyvBuaxmho8j1NldvfgbHI+Ne1+7t41qTG8Phb8YgCwZmQLElK8O5tGexaUSbiCiR3cXk3v0lXg
u1LCwdVX4MbA6uz8e4lYlQfkm/xAzXP39F9Ej/Qs5/66SBXrL2CQCCun+yYfiL5SexQ18Hb80VfR
Xefayovly6mPHQjeEHob0ANKsI+nWKisgAX5tV6e7ZAAKHbncnRxtwCLywuulge3lZb9r3bAo38z
ZS1rSKFLWp2tk/oWNx6GxUjcGtBdbnozERlLfwj19oE8qZFvRApC7JDdkmbSFhT1V8js8WHtV/qm
mufsdf1qE6MZArMhpC/Dkr2qIfwKuyiJ0XyXa0sUkbO0rCXGA3hsK3oK+aRDLqoRLqqM0kGCUMOv
EibsX8dibm6+bIhVmXw65cCjaWDE7KExRicTaoZGnCpIhczgWzPAZOf8eZBJi0ZDiMJ0xj2DXxGX
G4BgYmM7SGNIJeHSBSLno6XV7jo+iEyNvjMe7DZQv6z3UfZYsZWBYYcprNZw+z4AyHApA8pbVrWv
rGByk9EL8WCGD5UA7mu5ytsGUIzWoyBWAWP/ly2o2kBNMEaVJ5fV+kz5lDAvy/oBdzuQEB8jpYd0
sSKWBl061Y9yIiZZ2RuYS2xSTw/y04s9qoXx2sbfdbj+BHHTaFPDGsFn/B/RTKsdS71ycYZfzGzB
6NuyzzbCpt5bNkKCCaGM+7diEgij8oCLHsKBcCoODzyxXJl6fxdAdFwat0/i5z8T3VkZYYTgPVk5
yV2m0v72mVW4gHoJ3dNwOWL5rsex/2WMJPB+s52956BcRB8kX7QWGfcDfSK415pL39jKk/0sVVQw
U25cc2mjvYa0eYBNvY7HR9jAYt8KoMgbrj1ohYW5bC5ERPx98cRnNzLCKjpTAXdmFIp6ausRmn5o
bjOYkA1WBPaX/7gShyCUXzbEuyjfzI71fwU2NmOd/nFFwQ3fUUAG9J9vmVBmMBDQ8aOWlIzmGRn6
rN/Kse82UwvOMl0mhgfiztBwE7aEtscUGCn1dTVoFnF1BNMkDENAMDUqXXgugCwSF3qiOlNPropL
3N+aXQ8PR73Dt5B6V1iKF/dVzlKEVGIP/UNpOZGxS6R9zXJ9b6zIRTRrMLLbexuQ9/ucNthxkyzE
xseeTJ8yGMaSFPTK1LxW+8s9+m1x4TRMftIi5TsNJq0k3A5UFqwVsUl41kScdhiYJfuo/W2yk+oF
YqbQ9K75IdNUuxqXAJJZQieSxFyfMerktdarX+EsMe9CEznQKA2dZl1WfGw0l23Wtcfm4I5Ki6Z1
+n6JEeOuWTGnriAWX3oKzIf0ZJWHZwa/RWng68tDIm1mTirRC6D2Cw1Hwd0fkOZfkf4bgmmSF/ji
uPmFQw860IUN7YDR1fWFm9AoHgs72AvUrG8dYc1DiuMxcr/jJrNcBa6v3z2RRwvO7UZz642lB3Yr
Sjl3yaXzKoiwTd7WxMO4mKDWRy9Jd4x7fOFGFSBYOE8xUvmzLYsuynHJf50j68c8xGWVRP6+SSQ5
51QuD//kyrjzH2yTAlWyLHDESCTMBil3iMe3ClBgug91ain9kem8zPDP4KLpHMipqmf2qUcmd60X
yUJchqmjtLYJK76nQtLCUDrO7EymYxxRyQH6dutraUhrjc8AzJogNFP1BmfG3It4FdZkVSF0rR5J
GHcBMIgNi9kfKnL316R87IZZRNJ5qQu6t0P01i/q52aTcYdKoazd3i3DMVEPPUeyhBojY/gxDYSC
uKn3rWdyeMBzvDdmnc4vvLQCF2HEvXUUa+p0C0yBaVKgs2ErPjFJYI3o0wLHKB4F+fs/uBnhMFco
UDxeH2Jvx8LsdCLRSbItl1buCQ2Hnt9F/Ew/H1cKsDS05FduaRp05moFQLrv6IbBQ9KzbuqrvgWE
crJlQYKEIC3JyQ7ikQIpTdpcyouarGsqhEkCYc8orCanEqz2KrIDywr0gDqfgCCFVQBqnbzdjVjW
KCdYwbxxWh4tQv/L5AvOqcH9Y9JEGTVk8QTzPsub2kujW/SmBgcfjOAZghmm1SFQgSj9TTrrwfF7
L5U7EdIL8TVMqy2Ycvsq+S3S/xteBNUI8/SRCvhBdwA4ND4M1jzyT/fGOKBvwenVz5z8gHPureFD
ZKlioD1Oq1XUhJDdfQkFfPm87n8CCMyH3DBbXC1XIqv6Ow0MXZ9Br3JIuZiQ8oIAlr9dSaBEKP+q
1p/df/bddSUh7VZEAH2lHn7IXUb4OwU5Oi+IMnNW8euzHvsizrdDKyTFRlZ3x9gbzEtvZUkN/Ynh
Y1TQ6nGAcG2zG4FYKXt5SBn9FAT/Z9/Ki0gCXehcFEEY8uLiWPfkHl+otyQ4ls1eMR54FGSiBWyl
ittDOlXuA8U2bvKLYJ0R84Xgiamj2zEu/RB6HxvOdcqoYRbLobaO/5Ge/K0KlIZ4eD/vUQCJs2yy
RikQI0zM+CUrfs4uH1hed35x9xltIWS5ntyt8MY6ihELIoP729ieWHH2YjoqDF2lwgIJijN0LhZc
8/zTOi84ld8VOxH6vrNNLa+RZfJZAK2Ca5Vs7rJM53Jsb7u89yXZkHLTMi9aN9uSAtLiIkZEscen
ziKfxjnt0/XNLECSwISV4x/upDnwHzpaDxlE6UyX7D3e1Qrt+wNilJiCkyDUtit8hU2CVw6mnfrl
4aCZBH8U8LsMocCXVrC5vbIK1n9wiVqxV8IBR3DFcJ+8yviOdPhaBk17KAAmVBgVjCd4Cu8tIONo
RYr97hY86IMHqEQB2vsy86p3Eipjm1O43+mdgAquuFeyP30iGy6kRc56q8+JaAb+H/m++mWBhsus
FIxbjoG/cIjvtUqk6ZcrSaNVtX8dxQ79qqtgNp48/sg2F0pfCZ5rRfaApD6fb5Sgo+3u47DqI+x1
KIQ/hCCuH9zuD1MgG9ZbsQOIomqJ+R8kQNovw8Lpuvucf7qlNmIzRbRyLaE8dnfg9gxZPYvP57Cn
jpWURjYjwk6mA2FRF84lKpWdQj+VMjq9GBXAY8e2oeQfa3+HetsMFaQGF8roFYOFFT31yVZIIp0A
ez/Yf0Bcg37sM4uUkIJdufxbkJ2pXn9x9HdUutlwyi92t5UgrYcANnyS4RURcijdk94594XR/p8W
CDnRHqay3J9xKmaVUpcBftOBA0rbNdkbIU5ENrXpSy8e6J3N5voXie/4D87II4TgUVNqyUuHADgs
kYA748i9KaHUL1UOydPi5z/GppwGf1IhpYPze0MCU67npvHhxAC0ECaxExdHZpdw0YXKjBubra+R
Wkl/lcZJDfCBhC0qrPzGUQrfpeVV3L/h4DkjbiXR3HofAFnyhYkV/5gFHUr41J2fw/ahMijSxGaJ
o0PN3ck7LlvDjvMbYu1LIlk7YM03ipbaXitHZvEHNfzvirKsYr3RMjyyei1nLAMHrhcVXJGvmz22
TZnYKvrbEK50zlE61Su0thG6zOvsGuKD0KEp1gTt7xpjtbBSZNuecA987JkLAQmsHUULF3mhiVf2
mEH1oLh5axsR2Hdh9+kJ1Q2gVGz8ydse9Ge0J+gytYWnyP9RB3W/vyWdfqesRIj2EGHUOnp90/xJ
nY2popkoqZCkJX/G+zsE63KIyRUeYpJfSFK656/zAKJY+JTNz42FA13zDE/ezKeiVhtMHU4Yi9kO
dtGSx6Hxtc8luHBoJ5ZQg4elxriL9WcvTUox2bTM54ulsaAp48pPn18PgVnOhOfsumjkFcIK8lLY
wQnxQmb3vef5NzWtkucFPGOSetMM4Vf7z2yr77Zl3AE86tSYHXPyll6D6DIDm/cJ5mJZYjnaNvxZ
9cte3gJs4V8X/FOciKKf0DNLS0HQBaMTm9wdrSIWOCC3gDx5Nbdv7Eb55nX8pIm7s7CqAP3Oxe2O
nWWNfNk+PrQW61ioXrZKTdpGwmQlTtnEncpETIDng0etAYfSadMHKzaCTBn8gip57tbnKk116aIV
QsegaxNyJVXGZ/LhAFvQd37PH9mDrxHt2idWcfuhJ/Zz/7o1qbcRc8qIWGn47aNmYiT2ONFncmhW
PUB0VhIASNHYQ1fbP0s0f2VSzJAu4lzQv0fNVUMxnTh82O2nuug8mU/Egz0iqNxD6sFxICAeUKUT
AZmXxHpqncpESXG7OQe+2cW0HdhTEYM47AYXogMLn06jHIDc71WToLcm3+gglG2axWP+lEfm/bLr
EK1oWjsfZU5tyrVkmKv+qtmpNTJkgezbiptzImcUEMa/dKX7poa/9ivosiSA0gHuM/gkLYerOSIf
HJjNgHDr7/IWDqIZTsA4NaEP5WnUwQYhanYUSmcyD5FYiHoZP94ACzmDBa9W74+PsANtYUfOBCVm
BxIQbF+UDqfkAQkMvaQujakZ3kerS1RfSrZI8/4Su5Ymbz37ajoIkuPP0TnJX64dOhFy6619plp5
8IAyx2XxLQvD1N8kQOGIqvXaCs6ON2qjS2VB1rpyAAjUvU/d8NyMIILrZJSWMqAJLCeW1d0dO1OJ
om3smFIoOgpW+xiwVIK6RYhYF39zLf8pyfLhVeB9UuzUyu1yVwFkeB1ebx2fDN7SpH7jbuVJR3ZV
dqO4lfv5kxoSiKOijnELjo4+I61zjvvXbAcreqgSPV6TLYRV/rczd49+qk5YGEo2mAihqdg/Mqzo
Vkgu7RSjIGa0pRJlZ7NE6S+uT1hnVY6PiFamjONr8f469laQZGDuXiZDkcs8N5v957yTnRgEDduG
D947P0BKaitsC8b9xpA3t01husogfDH0ARsc/oZkdgVHuDHbw8FfD1OICOyH9fXbQlI8yaUzU8mf
6PZLJQJFYVsJMbx3Lec50ypA91hELC6rmcdY86Ph79Omsdnid7zhc+geiNvhahFM1MXv+YGQQKdd
lHA/HHhVOQrgI3psqy9f026aoN2NvAnHI1gQlgzlK1rk9OthgZvCHuBIi55J7OJkQwe2I6TSDnPR
Js5rBN65VEWrbYJsAbtn0JVGyMxsnI+ZFX1Q3Fv3o6W9S9hYTsrCFXuCmHJfgzFJKRURVnwHiZTi
KEHFY34Lv+5lTYIbd1jAhwXp7Naf63BNxl+n8Rq3MNv0i/TWQ2ieKCA7zzio+9EQlGjwuYvStHdL
bdVRG2dZMfSXaBx0uuArWRIrYaf3wfC6TCdVMmdOTTlnP6AHFlFi6LV8fFIlgNwhHcCiyxmuOO+B
DbruJXimHvpccyNaNmtqKA0TqB1ZDCltVNJyy2/Cr8qCD0nZMeRPEYnAVBPPa2Rym+A22z3wbjvg
r5GNl57UypstgVznYz6STlotIU33ZbAqvzhXBameTZedvMQAjfp+2n0IPTAyzYsMpnYU8jRYuztM
v0C0m8ajAyjurqJQY788LDb8tZaLFQ5TKK3OGYc+EFt9LCa4nZcQWOMJlh8inNvK+kpEXN+lP1db
9NO+bPefUWe7UyIh6Q04ltWBPqPY2dIA2cr0s5YKhnx8eidgHLlnjSFjn5ihTmPyquNaNrPln/Bl
MnsVDhcHLx0qWt46GsDGFQf7r5NodaXUMTHPk+5R0XjD4iBjAo7D8CpIIgraEJA8pd6H+fNNJJ6z
WqgAlkpUUzYa8ekPh8MvCfNVRcPTG6ryzEjfuG+CEBDA+TJhIiLfqKVDvIUwrnmR7bLpaMuxEULn
+xwmt7F9aZY3e3QFnbZsDBgdLHQdWAcqxwoR7j7jvuK0t+MjbFE6GOpbWRBUPojDo3IX+fkk5GE6
ofL3OYplwn0is7qno8Y7CkQriENdxXFmajReR1ygS8x/wfygiaMl0lu+588SbyYyrKF0VB42OGLy
hAOZVfGaVYUhkh2Zw3aytRGTpHLwUJPz3DbNJhBCiqZjhLDMD4VW81KvD+FOo/3C83O/rtPrqWRC
CM5SBbw2MYRVDBDEwgYUC89lYBnmUv4MkI6W05oTiTTZoQ82JwIcoUtFffiUySL3QMwuFST2Mdbe
CByBftj96X4AIXxQlUcfbjpWEkupNh77ttyFdcMoszUjMMSpsFhOtexdyHTi7EXEXGooXw3KgH7O
9fPMmMN+DR9vqe6D23UXEBWOX14jASieuzS/HVuljByckGh4eAWrsIBTxWJEpo51QiJsu9Ap13Yj
MgBlqgGxMonsnpYxddNsz817jSQ66IuhDDrYNb3NTqfZw/j/JsPB5+Qc7Qv9S04TQEHMtUF9K/Jn
AQyFXmrfvKrDXimsKV+looFpAMsXI7wSEVC+fpDo+gHiNO/gF0VrGXj3YYFnmihBZAABlPn2Abq5
zIicvXsZDeJ/wUhKkf37MpQhLPk5oRQPUOECQ4MsVyzuVy+J7dilB7ppCQ16fMY+iJi18+YOLgt+
V9R+lKa9Ip8hRIjLWLBKOAWWb1aad0Jxsk/DRJIjxni6U1e9E9zuceB7wskxeGWkOPLpOoFAeO+I
1i9iCbAMcHRQAnmxUNYf+EnTPMC7l7+SJg46qTcUX4DTqkwdbvzIzvjYEYnF/ybrMiniPiTqHHKP
uKEB2Hpo6UZZyF8doYICjanFMps5oU87IoClrjPRgpd4CEsLZF2Q3+EU7XRgL5PldvUkhc4VwKn1
wW438uzkfdRyvl9ItSFveOASzzO6yC5Piv76aAbb7d/30xTNNhUkEdyctG4iEzHAfGOSGSKA3b+V
2VKRv1RfeKwzmLD4lJ7xpnmNpAgU1wgaNxE5Q8wvyhm4Nc3/eWZxvomOuusSW+GUZWTMwHYesLen
BI9pwTAzmAlYBcfTQFr/H3ukKZR+wv3nleLdVDSOdOCSw+pFwGISnSdki+cOm3jZcSb+ONf1CNin
EtIYMefR28fAIFub70Pq0Ajd7tk5TVfqA1zEZgOvEIpYiEh43hPC87mPQs0j2b5AQkXt8RsyRCob
cZwGMPPTBFWjP3IavV3YfdlOYnbKrdnBV1jbzBR9gx4UMF74Q3KjCRjkpew5v3ldclXapH3Z+acK
kqZ+XGZnoSNVTGF8Oz0nGvrukfw8uND/DfVyOs9GW3fC7SPO49GFKy26qrbMzNDWcUURdKnbNL3n
ZwkgaZ57q4RL9N9KR1b7FswST2oAgGBTGgxv/4RKHBu/l87cW6d1JFbgtfTYkyIbitrXOjV79R5M
4r4Az7iyCm8mrPicikLSPpuIMFmuq/GNbo9GCI06jeqnVm+e6fFOptuiSIHkO8j4IQKufAh3k8ZV
OV7bayMdo5mQyVjFDquQP8wecPwLxE7Oj8EVkAf7B4D4bR5r8PoJFI48Xo06pEqbvjafeiMsP9ml
wYp5QMCK496+6CwLSeemhM+XfH2EIWyW5WJArCpHq3yxcTkFlBWp8T7eMsNRTRmnvax+6XC3Zr/5
0ZwX9TSp/6NADEpU38B5DRi+KX6pSxXZd0aWfPZ4Us1JPjoxvkWTyM3DAwoQF80XU0LXMQ4dO0DF
bnbv+dl5e8YXHXYNv11nUMU/VPK9s57wq6j3QrA3xo4dzoXEl60/Zy9NGx8R/JwXT/m+nQzpbYdt
N73+zcBv4/YX9u4clphTv2HkNbl006Jgr8rLPRTWbn/Bqex7X8LcmBel+AGd0BMDUXYlpQpBJ8H/
Rg0vNMAhBWi4InUTI3Z4QOUO0k0zoQp8UGlkNsDwvTohW6ALmcc6ZEaOUAdVWOr8F5Yc8dMpCKMw
kpLcEhIWkn+3yZ6LAzpUTv94v1BThFOQHqL10B+cavmMKvJxfei57H1Zf1C4yzPBcyfT83RRCUFt
pm88tdI0w23oIs9+c8Cn9E7kK+TKFaS/N9bYzqWqulxhm0Nkz4ccnLWq/ihptt1Jk45MHi3c1D8S
4yJjSyIsQZoQeFxp3Uins05Fosw7XqvfUPdEdA0Fl6RQDDDfuSVr1Q90wNJCtSjaYnuHNsfwgp7A
IOHAOiZ6zZ1TuP37jpJyIZXCJ8o7pSNgXrHX+opFVKK6b8I2uEtW7Tq6wopUftmo8zxsup6qRCrC
kIpQ6w1NJenQId+EaxeoXdChlo2AXugtOHDW9t6nPgSHlivG6370KPCTdNpjrYu2iXMBpv3D4qgW
WDNMhv26lJYRbRxH2nURDAcM0RgD42hKa5r19/FbkfwRrvon5+s7+U+qIasao6L+x09KgNVqKjQr
HmSncuiJzNEhwl302nv4xSECmp/EmASbvdOq4ShyiOPa7+BfnBDVUctBFDy5bWxxPSFd6Rb7P0Vf
sfy3qj5JhzM4wQjW5N1J5S1aN5BglALsmfG95trdoyz/fmHmPgUZnhw2ScjwSq0zIBYlRWtzn+mt
fdIpT2IZt4ZQraqlwndm5uV4JJZ17XEves6G0aVKt7OGkxm6ktCZaKg+sE1I9FvC9nnSD1xkohCm
Vx7M09y1czRPGDHb0Gq7bKU7N3mDnn/KBiBw5O2B/doj6E7P1bpdMLKI/Vonq4ZOMP9cov0PQTWU
HNMNLiQdjBIQZyWbwAqS/8UUPVWF/TswjU3ccgQCDNhJAiVGZN/4UiWsCVCWtUo130LLlsGITr1a
Q4iF+NKQDjRyQpqKMEdnjvmvzbl25d2QAH6IJ5jGiEUnxaBP5b/BIaBmfaekL417RvQYfV9yDQAU
U4yqhu21kMc3X040LEKI8ZWWwPQIpEpw9LC2fl/DTo8Tyr/qsZziPuwhSaGLdPz1Aqz0SBi6qLmK
k/IsbN9sXC5eccHziPG5vtNQhITkfl8w75Yl/0NUe6UX0WjL25ujh3W9jP04A+tt01g8upSxs7a0
mCzIZr2+PBFnj51eWuvtjn/VA/0AFi4C9etMirq6fgBt5eHt47iFfAM444PAQkdXLpyaH4JqvnkR
y9tKfmqQk7EdJrLDNJkYfdeqUWpmkiCOND4mHdp7+2HwGtADWdGJwKKMyGvAponrYzqpJZdf80W5
ixfUQ40uzLguv8gh8K/XEUrJYP+qRejH433TdA5YsdJGPNBGhCxGa0owMvRJLa8WDZ31t+ZmnT+i
WcPrQ0LBx1fMcn5ckyg56y/XqGYA9oJF0Dul2S8hfc7cbfYRDj+fmVFPgp2lqs2TKoWpy4OEajmY
oEQa6p2eV7q0QAWBXDi3DMxEtXIKYGyYmO4FZqZFDKCP3K2deGdUzBv6prD0nnZ3DZNc7ii/7eHX
mxkiVg6iy5OJ2KjLYEFTBz5g5T7pdh8oXz6ApCvRViGunUmJ1w0bxR7E2no+BwNLE5loNJ56gp96
sDawKswL/cm1cvECPGuj4f1tc6AX4W58gLKMO2+46Uvr5+zUyYkzJ6PqOUVQXZt/0frub/SDjYh0
U+1BN3SJkQdO8OZU/hm0sS3Y4gZwVztQZCgA+UNcJIjyjXpHTvysSe7iUoeHqce90eNYkr04o8f3
UzTOI7rvN/d9WVGqmcUXE/aeogZgcGmTq7S5HCFBOGoZsUlrvAnnV2NMA+GdjMulpkCCjPg4vVri
CFXPFEH8KzCoeEiPaAD2WpVOAIv2hDf6Al0n4+sRsjWAI19BdYtW/Z3pAk6AMWcEIWNQfOT8v3Gg
JxHobwvJtDt3+LCDbQhQDmWfEvb71s+FAZyM7P8zH0SIEagxFxmOoKFT/jJXe64yZlOB0eRmb/cA
IHunylnFXicBovh2oPHrunfT207FnuIertIpGzErQBl7LvHRCpxWpPUuiY5F/N7JOo8Xn1Cso44e
n1Zs0KJSNoQJ/YmUlcjjyULJZjzo9EJb75T5tN2TlimPrbQ5hBTkQeoQvov8FWqZVYAEKdTPzwwM
rvSqQQP5aZfvaimXWwPuOvYhjkPp1YKsUUudfsVA0AEwIVCNjQ4otqf9bMEVJsIC8cf2F5HkvuSo
4vf0mKfDLIVJ3gYNs8EJ01PmQpXX1OO/QWmhQp+Gf2OV7LkARSzidZ0jyng4Ss7yTiSNBq6JlPJ+
54yiBf53eTpZDqCR7lSbXh+YX+gGd6phhnJ9N86xjvtJREYd2TEzYEwGH7DTO50t5qy3TfXM2h9j
+JHylxovImVdR2rfRIYoqtibPKevNQnDYlS9+sSOEvmz13Yx45q1tWfRWYCQ7Niw+XuTIZOlpahC
j7z7djWcFY+eto1AOJVuvjHxt3L+pV/qs7kEvezhmnp/3QXkq+5UnoQI664iy1taB7awNCkfzVud
hlv58evMvkH8J/6ff00m3jZfuA+pCG0+2MlRZK1V/WYMNA1f+QZ4GDzg4x1Q73/iWuHGg9qhmU4S
f+zOWU3IfGGfPCBDFKvzjVjNtly9r3Csg/1OEHz0ZSNhSlfhiXduzfMCPJLHymI6QtSaC9lrMx4O
gonF3GCVS5eckOpLAXoEeXQI7zLKN4Pcy+8DbRnGqOvGE6QWM6AchKMrV/6nmUEVAaVduLJ0/pMp
GqHt7PUzQ9uQ2XpSTDZrubl0SdbyMMdQDoMHmterK8lgj1q7bO5hfCvrhcxQvXyby4uyHX+9OlgH
1Cvgx1+agnuG8RHeKKI42HvGcwyIofP+klEWAq1dZjVjrA1jlp5vrXSVYvfKv8woqP2XJJ8AIRGR
i1ECgmsZy4vSwZgEbk1BIthsH21c5JaRtC8JpS4dPSnLY0lJfworrBx1KS+8d6w/S08jUbuUNMv+
/1Pkkig/gEaFhgwRJLTJ5N3msQ2/6VQWSLk47zptClPOen8LxymGJKeiKKvQ6ZJZdbAJloJXdr8k
rwQC7L7tHoN2V997fO0VnU4MBJ5nhFaBYEU0DaEo3DLOtM198c+rjim8X5dJMBRDarltKqaDzS/+
pfwZxiMdbEyIKBP1gxnDdGa2U8BstYiHw3JaiE2Z/z49WGSYlblp38p/Hjm4QBmPSWZdgpBSzSjJ
QkAPv0xpJB5UsBV9ygYi//atIzVg3VQFDY/QbX0eBcgNhy6XH6QS0RoyKvbwgM6u7IPlOJT9U0Ux
JO2FkqYPm45u0D9BZCLnpUKTD1AaHAM/nBgfIPYniQwGW7DyZcHeMUPiZnjMWMMMLt4gDoab3W+J
6i1P/vR1yyXHaxvxUiPDGB6q/0Jw+GIEg717fgcZxraJz+0hvi35yQLuBFZt2m1VPLdjCFjIVgkq
lc6gZ7Kat2Oj7sHoDXvsjFTp4ZCEaOFjXCH2zQPi1fe/cm90QC8K1YMZfgl8EGgsVk7aq0EJhxsj
x1xHBUZ6krRMNa1Qu1UdWR1Lzt4nQI8ajWPqEFJqqv+FhYalchnwmd7EsMoEZ8wnF1tx6xD4IzTV
keIbQXvZKPm9Sql55YtXKD+PuCCtwOx8LoN0fAt71RDfrXR+Ffli5UUuQz2KTXNyWLHuIvg2A6Zw
vTupsJhuP19en2gLV8o8prpaje7wBk81XohYkCcVE4J4aJaUTLIQzyloIiYIZIDXMn7DbFi+BklW
/Oh5/zAUi8RxSEuZAiLU1PqlTm867G5MYLmD2vUpdGEuw2C7PPemddxHSCVICLk+MevFWiYa4AF+
E7e7EnqPh6HeFPt8xSe8KGlLDmuAdiL5QGGSifilyQmcezcT5/ik8GBBuWlYPog70CdbGr8EJqtW
j3RSgEYxS8n+lsARC62hwmpwRbE3pmJNMa03heLQtEwia9BRnLarA3ZUIBd7bO6rLeWCa9BP3qiT
h3cDJgh+iZP+CPxoQd1ORVjVoFK7EBJfW/+Lm8E6eInGMDNM6lfGD1TIKtEHKed/cWMDS58RuYSN
iPBnL3nfI2kekIRcdZYbv0sYeO8/y/px/cwE5Rf5tU120xi+V7metzXObEK7p61YhupikUeL1T5M
hm03yxYGd3z8MblYcBsDt8J+uz4QDFDV6x6p5+4A5dJ5Dh/qINm3GYv5NPMScaq4aCO13jk+LjuO
f6PzcbTXoN+cfXQKWz+VIvU/XbulaU7NRcx5vD8URrbjRfGTYhaxe5GsMLvvjTlGLImTpOxkbn/o
bCOJ3rVkb10aTcexqJinhhDDL8DBFWslPwS9D0Ve7rU2w03ULlgWp6UhTsLBDnvtmBRh8AQYb6xO
rr4s1IAsGfkOXPWuv3YemDR39Nia14VwTPVXfvru5QV1CZDUFYvH7Tfc1EXM6oLXOUZYQMBhVMzK
rGA9E8ZSdn9jqpebrbpgQzhcYmWETp/RpL47YnfiuXxTo/4zDPhYGO1RWMA56D01To0flhlWlsyi
3BAFkJsRI7hpK4ZMTJashbtuPJ9tttwaEKUxjk4AbshYzN6Qka/QcsgbRefswYB3Lc8MAbkoL6lo
/ajsQ17V2X3on+pXnTWVxx0lI4NRK4ymxes0TEwlMlkgg8teETp3DvHiT0trudBzT8pi9VXPMLse
cJyawOXpf28AKhLQCW1HPX7nMSZJCE/jpvFY1ul8P9vbNszM28LS7+hIdFlu9NpN+V6mW8MO8f0j
beZUm9TTY0x314Gzl0Cau0qJSCDh+u8aIvCYV2r2hq3gcj+AQ7tBAXZoTbx1myW4KO88naGgFBBP
sxJSI+XANM4XrHP03Ykp7ew/qHmbb7oHPVMmnobLNUpxkjxCoCezXzA9aFPS5KSbOaoTqmBX8d9a
rDpyBz68PvaoK40lgfPklXq/784U6pOe1JNjx5m8pbLIGILdTDAJAGMNXHkzHEUj4hPCxBKwRleG
z/MIDoExkJrEEtrq0JpQGSlPlzIkpLxGOhOlJH596GOfzYzZy0x20+EZiDlPqhkwa4nmsfAjcmOy
exgMXauz+PiVwnkspdmLbus4BANPmrE/NoD1nvNYkveqNaX6MiDAL8d8d+aUrsyNC0rh8ODFMGhm
/wO/dFPEGpQ1jWClfFT4nonCTrSG135VPUmd8ON9AUYb2Q7Bgb2J9ElUEX0mPjx3p+IolqELE3fG
NOj56eQ9YNYTUPlzkHhW2iPU1YN33ut2WXIDOyh3+s/NtmKTvgta0QUtFdtKBWGQ18ik6t3F4inn
vpQKLBKSauWqmziiHXLBtjoa+nyytnY61elB5wFn+WBOZfpxeAl/IiUQtQurxSqHyv0hoMLUjMzE
0yYKho0J9cH0ftoHZoWD7iSb64SAq/oiCg9pBA1YGgmjXHZuRgzQP825VZHkp0I71ZVUXuMAze9r
DS393H5EiGZFPBp/tAugiXS5qAuWl62TuxQykKKW66F4RhTO52iQb9s1utVq1nfA16GPshdLFIjr
IfHqeyL+GWYr1R0wY1QIK4dcuhMzGm8CFUmdJW5V00z4hky1hZRiCDh/Og+CYccSItOhzrpbmFqP
tYato7Q9+VNrFHF6CmlAWrTKuO/PC+sdZQhCJvUnv62ArG20YthaiFh1n74tozFJP9hnRJXqfyoe
BCYIdpbzCUesAr+bi/sUVNKqmRpFyFLbL70RNeC+YbTHg3xCYc2KJzPWcjXYcW9IH91m/wdJ3YwJ
s659SfPv+VvbGqwzRCN++QotHCoDbVhMrVxeyyiYnttuJ1egSMLgvYZ7SVSWXw9hDFLULs+E6BfO
gK66O/+GOfXrACQeCIik98KKPMUpEUezroWscrWpLBWB/Eh/zbwh3P81POBNzl0piHSd5CWZGQeH
Mxjawi/Bao4SCdcXHTcZN5GYoZc9KaQHX54Lgi7jG93opBwXXMUMIDG0lv29+bwA8m7nI/jeggv1
czY2DGA9Ikh37JJ37hC1ICtFmsQW45Gn8AzBbQ6B7el/pR0DQeFW1AQwfrBmlTScjnPhsCy0d5sa
l8qJGIkBHDOPC9Nx1+C5o6Je5oy0lcBtA8f/AtCL+DvNQJCyQvkVnJwFzxRPV6qpiJb5EwTDfus8
gL7SyaJvvc8v0/98zNBQG46gjeMf3lHUfqsu/swLlyF8KwrFZxPWRNpBrgthGi5bkXs+o0J4DZ4M
DmjCDb0XClQHcyWykzxpqodCe5jyE7dJHy4fgXc0iMS8RghMwOCTY1tMbLH0SdPTcMA8Z1yr22YJ
YbTszlgbuJy4tLuLq6wbbFdhPJ1AALA425wrd8yMItsZyWyHqQ2aKxDwS/sgpVCs1eiAm33DvW5F
Pm29eVo2h1qpu6vx8ZOeGdQc/FSh/KCsiQSxtsV8hv/Q2GXbha1TnND1Befu9DKejfNfSCLxbzNM
4kAhoNT84uilO2UwPXhEmPTcvjZJlV1o+YHxKe+b1UvlGnsNKzrmNyRLXEZE1bQnhdRjafWXRU4v
s1VCq/y8qK1KpYa94fxP5q9DWKcUMwlsS18VmdkMRykTYPqN90ivlpyP0FtNnnVS9ofTqNW2nK9r
psy6WfbTG2fOB41qad+9jEb9VzUIHX0pgHw0ymBEWbHBYdYGJoJ0+743lJhuOcxaI/xkMnYRz2xY
Osv0XBm3S/YQkLDXpREm1MAmzcaY5BA7VUTTTHPkA16Jn5byo48BAgHnfmNlTMTgd7U3a2Fbo7Qi
no0OkJcPC4nyX31X2GuNLs31S+Fli2C2hE+50XVamsevre6R1FWHBrzrdVL773wIZEgWbCiwDth/
ouWLFgPE1ecitxdmMWnPez3NTVy+IfHYmo5n9QPDQCQ+PJyI8uuuNHEFgGql9Y3rdeJMnO2fWY0e
AQvUPC2DBCwuIg9eZSbO3+AoAr+rvSgmS9a+nOVqLA/dnR+PsjMMPJMUoejyTZwwoUSTOPs2uNfO
PrJXOqj4llMQcAo3+WkGrrPExcBIwT4tC2YX1mlg1X+8Uesg822O7TgIfXt8L7R0wNjaw5asMt7q
ztc5Bg/SC/bl+39o8MSU0ZfjmRVkvLHzSZaTR2sFPdUfy2YcHIWKAviNJaQmwglKAT954Y1pnoqx
wD7zjUaeamsaxoNyPz+eSRIGo4kleasY89REKx5QPFjc0BzmV/wGTr3xbyOm06HFNjb+v4UY2CIS
xvH+r+SFfIwmTlPmnFN63PT1r61+vML3//qSok1BKRu5ZqpiylmUwWyFhcpyzFX96SU8kzN+FCs4
0hzZA+RvQYPokO8INcHvJXkyMy5Ch4tCQRKqDYaW/1H+N+Mnss4Y38yt6Z77ZybLnyCEIrS1fjAg
XXc2nLTg77U4yGXOy4PE9WSdrQ2/LxQy0nUDocUxTx7R1I73OVh8SoGzOd03QlYsPvl/9TwfaljZ
j57q/KtW3aGOLqgJy46/n3FqLI1QyWBHAv347EnTuzINg6xYzkBGehGbXE12XDSapL5L+SwCsvBT
Z6HWHCyYx9IY1XvXSWziNJFIaQ8Bh7jWwBk3U2Bb5lYfHOLZfaihBX2mVvewk4VYaUW2XHozHdos
eRQ3CSO7zf5fS2EcNkBYQP59ZFeCN/q8tPXiF7cvX94vzTKLsAKfoDJ+Cp7yiOGaeOmdA27wxvhg
hmtCed6J8hWWGXa9svhUwig5LV3rINUQ+MqZaIEdXN6yKX1FMDv6iETsibaHhqjbUYpem14UmBQ+
SOyOkYwU30AYzIdtB/mZlwqkGIwoK2DE+crYe+Fw1wcqUUZrAhUuPkoo1+JUDiZDlAX+bcgtN0/e
YMvb4jJLE9KgD8nuvmZy6U2gmGJ1MY+Hc+MF3pe/B98fwccEJYf3RTqUcRFpY0QixIWzh6oVziu8
hIA7Yk2Oe3tSIT8Wk9qOXtzIijSOiF1YqJJ/LNJA2g+I0h2h+2Usxh2jPLzCHRvDlmHkfcDAy/7Z
D8uno6hKViKntcqDCLUtBARCQhpBt57VrEgaaKv/sYrIE2SP149aMFHPzqcKZIBBFcFw7MuCr/LV
g3TZ0EO9v7i/L07yyYNaSqMiJAXMPdCux4maC5rUTNs9GoH47Revd1d/JjFVLP1KvnhMDyADw+XP
Ep5nxyv+P7HluHkv5lgf5hye9pz/NF3R4FoVtf58BZBqclVLWfuCfTGb20JrR05UHLJMXwQUP7yd
GHkIPKo1iyvKuywEaM2x/an3KVGAejJrX38zAdT9nqa0hPNyxFVCo4MomuMdxMNMXYE7OylVGXki
SAVxkSjdQSiKXz3C2abSqtUz9NMFuAgGEwgE6wYXmqFB++O5RbYjLrSVhAIbfv2UkzU1Vuk/PUwn
eUTXNd44Pf4tVM4jjrbuiEzN8gNRvJOAIV7O7eJeE8KqXRtwp23rGsQrJBW3ZdWqTBliSfaGN1uK
GXNJv5im5kMskTxqeUhgA5pejs1WIbe9/IEwQV9/qWi5N12ppJeyvt9KO7h38Mm5Ypzktq5pB2+K
5M35OmViawiJt4hv+4P4eod8+7l/h0bICJYKX+GuOoBd5xq1yzMxq940yft14njKpn0zb/9t3QeG
U1KaBm19pwk4P67QY++RiIpGkIHfhb6MySZdDXu9eAA5v04tUBQZleiUIViNyobzG1vnNjBMOgep
bfP5T1AUuwUTHVcjyrKs3+26veOaTOc01kv1n5UjWp5jjZW3lkW6rNSXT9vI9l0WuuGs/MFtmyAc
EIQElLw3cdE5ZmAZa2eIO0KvcXZFML9YaWsZsUrvUb5Xq8vxVXE3e4hm2I8Nn6NRDUQ82oJ8dKuU
Zkey8Sc7frGtDI07IfBHbdyBYGdhj1yKdYynCPW8WDezSt2sd8tCMwMGwSaXSArgFkzdKyWRHmVr
mYqDEDATyZZomo7ZVsVRd1jUiNK2edvANa8OTlY4gM9zUoSrWK0P15uA3OENT2akA3kBaFYiJoDo
yaltVNJOJ/yPzLFAS8ZszBgXgfsjVOUTz28zvVuseM9ZxU6E7NyqbFJW09tjUhpCyumQuryVK+9N
2eVA9KFRwAQ4mxkK431XfzntQJWLt2+HI4mh/j2zhrklmgsnozuJYB77nVjHjpqg3L+zshPzzstl
V6MH5J+VwyggxZOqPGzMdmDBkztD0wqbfZKpeo1/sowugvn8sOymicaM/qTmSn1hsCxPR8v43Nbp
mrxC5P8IJ9AYnQXOVGrzczF5+2Fsur6cziKy3tLPgZnLxrg2G18mwUirtYA6qiB9eRNA4xEQPKr+
qMkaKSq+tx2XdS46MhkCXOxJNJSy/pyICtMPyYnF2LzjMoT653hGV5AJbkVAdipf4Y7NUSVWlCNF
w8yeQ1nGNrnexDQtyllC5OF9WFm9AifK7qIxaBHFNr6jkp1hSIDklHqSkTg2KawQGpNb+0xwuJsu
G87vSOZiywLO8nIk7xhKcgldjSJ14ZiVTFoCp8NpeDwENnDKluXRFFOOfsFEbyik87Kl1QxIl401
3L6mQXmOeXkC0oMuQjGEd9OXmda/TfbGY44dfV3NZWhzHh0yL7uyJefH2GNDnKNO1MXN4SquAKB0
eCksopWCKBF9wZFJoSscFMAtwAJpUHYs+YcCFg1hESS2d9utKtpln+2uLsQQTKsvTlRU01lx6xse
tTS3+0NTfbZNjInRH0XFemKRcGs5/iCnmTe9XYyW9by6TJYINhhcfGDLEDvxp8qnmkiMTHGFImiH
1KLnOfR/lv7aQbJYuVHjPPzwfcHtvqpm881Tw7r8s0euonfsS3rQvLHrOJeQzY2CobsHF3CMSLvI
pVQwxw1AqZw4toJLkW4CD8WIM7wGuGSlE9TNW6CWVXXkJIl7x0/yBdxx5Hn/J/BaxBf4VcWcXD4B
+mNSi2sdgGywTXnqvE0G7RWRBkfzrHpOemv/vz/aJ32pJ+Knq7BIznfTGmbLTr1mp9jeSwpx0b3Y
R7yDrF5J1jSZQNVv7Rs9NPUPkEES1dRngr2RFP6DNgZtRAb7syod5zmr4VRNImSAgrmWTtFhcy+s
50hmDob/S4ajSHagj0w2xgjSEqPpt89QsIlyuq0PQ2iw0GQvpAuohvggFnqym9nrtZtdRjIdOENK
3kMPM0pju0DAmWoRLIpgmI18G1zvgAXznbt6mYpeNl9EHbPHaifwahA24wCGiXny2Xv3+euvyGIo
IK0nmE9um1SHvE5bLblgZfYXHt73laPnYFhag2o2iMVusjmIdatR+qrtjBedn55gROL7jX1U5hOO
oNCwl5BQWz84FqsN8OSf0Nxv/l3z02bADwCdwFJDt07MULWIA4nE1HFfxj0tFLoUIab29q20U7J0
GVFF/C6s33x8lf1HIpMJ2EWKXe2YKUruebnR4FyIr8YogwPc+UJztc70Y9J4U1WlN7Kps+y9rVos
ahisBtfP7wiyEo/be1SO3718IJ9MG4vviqq0Bg9WY7YN+5zreX+mtz/ybRAMmvsD46Wton1UGhad
Z+Sw8exyqxzHg6sGfxPd0zWqzv/bQjNeEATMSG8fDGMKV9mhnS0W9jqF+ug5msnXAM9TF8JxPvzX
WuNRATwa83E08A/cIR6QXLmyFHMPvcu3Ut//ZtTM1a+sNwJ4Ve+RmGRbKunmY9Eo0mDBq3JQCsXf
m2iBEtdifRBHGJel6KVevfDp4DFkS/hDeHiU8ZF97KB2Dp+IjMSC0GlFcP6WUIbLf9W8IVnzueES
/FvwY8uyYSLbvApzpSjWWWExpGOsI0y2Q08yUac+9WENWFoVjFBZJ2XDC062OMa95dstpsuCOJN7
pbOwOv4VupTJRoYW5cHMYitB1r26ykOKa/2ljTqnuRSxmaH80B3M+W4AilWNpAH+Zi1bcKivgFZ1
BDN5AJXKta8LqfIqI5VAU3BkOs4Z8csRPBLY7bymhOPE4uSCOfB/VLSfA2F8VBn9KPVEfQo4HmzA
G3SgZZVlXZMdK0ByfYFexaPv8SSSk0QGd2XI69wolLSej4l4/PBoAUzR24bUCgrg94EaTWOnrQ5y
rAICWmR6M7bsbw+ZsUjxzNk7cXfiIvfXthg1gHaoTOaEMBabznIMUYNGQ6ky97COvQRAz0h5LjO4
Z0uwbTWXyaqGiZXYeVfxlqVnw3dbgkem3Z5ZizKZcEe6ueEAmduV/2F9/FD6s+OS75X6lMRH8vJg
NGssNvAZ7IErXMVfIeqLfrSJ3VWGccVpTsTXOaYviCIxbIopU4tNVGjLWbiAUtM8+kxUHxazy2Wa
4er54Ey79uP90ISabrFTAZmuJt1R8vYmhUwLnDrdLdjY6Ui5pltxCW27Mv4Kd52U12JXq4+tC/vB
gGqarwOhPYisnlMf8lsxddHfgbA6CWpMMhks8rpg3n74fSAX5dwonS0ES8Tha2y6kXm5Lgmu6l44
b/PfQxGp7XGIkk8Mb9BGRyvXRDq+Ju/3DhYuGWgePuoLwyeVlSX/CZb0cqiwwDdM3TUCEN2UuLu3
5ali9vNXQcfudM2giMH7dCyCnRpp/FrwRDRRrNLKpt4bWkW00nA/N2Vr754bxgAFGNEs8QKG8ekr
ccqZx177i2MKFGAzLC+1FuA/xSyodYvS/JBUTpdfM8ZLbqXrrhHKy4N6pYflRT/BRaRKuVYE6lN5
nfJXa8+McL40MUzXV1r2pF4vxBM0VGRxFy5KFp/qoiRhFxIimqAnDhtCF0/zq79rO8YYrI7GCuTS
zy7MtssR95nctjXxzMrdkuBWhrtyeOUZLTBYfiLgTa4MKb1h6XWXghDMaLJXCNSSwthCEc1nCJdG
a2JX0wuAoYDIKV40ubYT/TL8Z1XqGnZGZr4WczO9uGnFD6aGmnOi3F2MLM+O515PYBBDyfR6Itk2
vvR5FO3UxHUlSIxFNfXXSfD8aPH1sfbVM6K15Uci3JTzhl30aRq0zKa/zUaNMsLIHIezQGLJOtom
oRHpqIGSKgyERgFDjjbdGxu+HWH2m1ATo7xxip9JgySsPS7pN5wLLlhEjLsGJfcVp3WCajOX0aXT
cWP6l7UD0iPSCkBL+vTqBJKjqQ1rziMl+wdsEf+/03hneJFp7o+E7Ugey9uo2HRrP7rCRR0BbBPB
Hk02rHRKzjbc9fyPa/jzyxDHg51KQtOH3n0leaPAHkTCMtvfijbyXK//XgF7wQZ2o5Urv5dyTn8F
c3PXI3R5TbONIrJ/tHbNDIdSOVrk9ekgZOso6yxjRNDLLd0OAlscesDO851LNsykYRi35LI5zlXa
zu/4Ev9258RdPG+/GaDx8HzI+q3B3Q5eySDmNn0lBOAAHxltHHlhEhArID65EDefiKGoR3RVGONZ
EtawtgzqkY3aNgKij5Hk54wdGJNuvN4aKdnlx1d6fZKwsSyHe3Qa2s4hOPGzUTPlfYSP2idETKXk
irHJOImGoZP/id8RvlMhgqBQjEOrozhn1NkmkO3+Z2mzeI3UQZFGTUhd7U+U7llUJosKR4fXw7Jr
ML6AEd7HtrCFKQlCqjV/bl4XFQ2n1egcrVM6fUc2+0X0Sfv4gWHB2o6+/FkWc9CjaZW/+78Gnxjl
1tzx0WHWumC4E3T5Hzw21X+mZHtRmg5nIA6fMbMib6s9n4WAItybRKgC2XhFEf3saVGz590ybR27
xV51jEqMtrawyxLmsdI7OOVmToywyPQp1aM8jpWP3z+RLtUHfZegZ0OVUCeHI1I0Oy5kGVu8phBi
i9LCI5UMvGCr4qywJBiL2+o1wYbUy+tchA0zq/T+wAae61wvgobyMT/reNRQO7Gkzqb/ye8+MCl0
izUn4HMCrsk9cALTCGOE/51wuSNJhWlMVTH+RLQcypfxZo2OrYf7J83XGIdu4rpZ0vfzuVUiHfUQ
wDJJOHb9P2YCtqDHpE/0o9Qe0lJYcDUi01Qz7FHtbVkjLJnRDLazr+zJ52cf3qed6TWJe+VGFlGh
tZuRxjEgiKg0wCTYCIRfpCK7oJy56rMbx+EIfXM/7I6l5e+EmWLh9NaRpKg3N23jBP1CTz9TthfB
E0LawLi6tEMN7h+KzrEI747gKwwshoFn06v4B8H1KKpAYkajXlqV2/5S44pLEPn0pfwhZVGYeP+q
MfpAvtNP68qWJFEy817O4rmvOdUXnuzTwolngJqHoe+x75dW8FH/73BksYgUT5cHtLjPEtnruvpp
0iUDBjMbQoV4QZArE6lB3D0+nsMdH8Q++kA+lK+OKLHthfXTTeOBiqjtLI552CANCbReadQ5lqFN
MlKCU6OP9DMfostxy4yRGQfm+5KG/GD4ku7oLEPeWRep0W473Xoqie1EefCiD2HGQNxKbXkpKo09
ZrTtQV6IBifoKTxmMUugK3goYGp88teqVZP34Y2ZNbdpembAU5sF58FqVRLtaWqpB985Ys3jyzy0
5qiPxtxl7IbiZPhgxIJMVhG2f3rqMAhzBz6UZisHbTmzbcevaRZ69BnlsVomeBNAeoAZrs0Q9pRM
G8FU4kapbcupZLCuz2Na8YxW3hzizZPuLyZ4qEbw41d6n6QEuyE6p0/Mgoydih1jQP/tRUeHKuM0
qbr2NXH+9RIZMyI7/ISAd89mJ34zpX2sfd0euiDj9N7H4ZLutp5tSCBPuKXLu8c9ByTzSYYW8D9S
e8TIlLI6PvFn5mfUko4DG8EzCw0CGiz5jIqZfijg61Pxr5UoHv6cpgisdqlKl47MJC/FkGi6JSBg
+wGvSPNLFRmej+hsBr/FgsYvirnuH6D/Wc07NNyfUg1qPKdTtQqhzSBviBS0tWi+tABaz9n2BnV0
HDpJdiAb3PF9qI49tgWNjle9aQWVxC1hzIM5fDIqyNC2n+IJfoxuQlkAHA/ggt3+4EuXsWt06FZ/
7urTlfX6hLqbnbWymPH5aeHnQQrUPvffAEMbdGsU2VMot2DgxMCNamRZmaLF7D18VXUEo8LX4YDh
DGX7g27EyzZFWyeLfNZ6ehVB7ZzUQyfrwVPfTpFTRvpdznARjujP6ojJEqh8N2VfEMfvlxheUBQ1
lCsOaE2vsgwmnLlZTND9UxpjIbMUPRVcwvwv+Oup0XZxo77NlUOEDvqc6bOURmMhC2XN049xCkxe
j3mzRVvClvSw0fyqkBoZAabsaTiKQ2HfqrBFLTDItyGAYValDVgRlVn3zE94U0eoW1yuILYINq2m
mN1eH7Qr3TyIyNZ49GZ62ZQcWwnkJmG9BKMZ6RRuC+Vxr71i0Kl3hmQxFq8p+eLJMNaUEfpDWk7C
kBvO8DSuNtZc5iLvbuiArMTZq1N2ZmEE9B4yq+XXKU2n0vTEYIRw3OfbYAQshZMstU6hVSGIcKSe
On2qWtW0C8mp7IyvR6KS687eock0tczKQeCcuSNHJ5oixCPAlGz06pluRNvFOBHhr0TTlsAvaLSN
lCXixduAW8WPO66mqm8/s6PgVnKQFv4T681IPONRIub1o0vjt017lxY2eFHqP4pyt8xJjGywdnZZ
VfWIC/nmS7ULxoXf0fLcDQmWdv+CS6V1wCpZ4U2TawJ66uaMtVj+3auy7m4OvxAytWM/9GWF3mPT
NYXl8TnQHamWJbCRmJG0VhiIrnQmb5+Kg/NSd0JyRnTWXmZJvjpdlELLpXzrqxccC7TwDGWBsspW
gzNKOYPg1c13vB8LrSXZizPHzANSd/WOittiwpf2DFt3BXd2lvaDZwcCMQ/IzE0f0tYTYfogiXQl
YJXYmxaOLzX0H9u0I8AuuOdEKRzPSzhuuV6WhBJAT37jAs+nRiuxf2zM/aoeKV+NCxRnbb+iuD/g
/CnP6LYCSVSUyzBBHKFZervDBJVgYQd8Rk49jbpdhVZZeApJuDou9YqdQZ+mnAEbs3woDJ/REgPy
7YPiG2p+9eK70yvLy0Um8UzQs4IFra0uI+ZFpeCpOAffEwvIa6kUJgFnDsLrQDM4ftRMXC+fx1GV
6vf2dSzh8ACRLUmPx//4D/EImbX5WgreHpOWGuSkciUmeiAgbnHs2TuCRJ3jOyqqF/JBngo41fo7
yZb2u3NZDYQ3MywOzsQae1zy1WwxDXShM0XRo2xixYWtVXev/9kNCG4B4ndusUFK/wUXpi1yPy8C
xBYFZrJfLu3j6Rt8cOJUDK5+rA0Qq1aMFMfLuJFIYhXcGr9DecAzYQ2SSivM5nPY9iC0h1sGktIl
XI0/Us/1ENN811+2Hain01LudAP2Xl2pRK9iYqdudgGGUPoNidtRS4ZebuDNXpHDfvo92KoJHNzg
NEbeghdk4yaA/VR6/0r0kD+ZVUTRpnMv0KcJ3NGsOa/ZP3Sp2GWZqC2/h1WFq3+SCD1gCqNTw/0g
k0vBeKqB/puBkQN9U9WFxcTr8EwkGqPeiim+AeM/WnQP92dwSq1BhVOzRq277dTy9fQXn82G3fDk
LZMaDrHVm7AkPqJLpWYEuzdScxHq+gKD9MRLIaeNIl2r7Rwfyp/ZPIK8I6dzfxH89lMgbAEua4vN
8OUup7Ah4Gk1FZ0hLro45STV1k1/XncxBbHwHMuyZw9S4aNirXbrtSkADecOiqDE0TB33yf4aD2J
x4uwE7LpiUBl/X5E9z6ECnURX/ZXuK4e/zlzMWjLwHSH0nU8xqsB3GlwhzRzHy2GaNA1es65U2kk
KQr0hGhLia3TqQzqDk1FrOFXy904ccilazzyRdplmELu66auDY3fBBKLCp/gNau3kZsVaDGMctOB
Sx1QSNMq00d8n6KT0DdYY2TENKxn9kPoJIpEoLPik8gfiMXDeyAZK559YvZmPrHmqtBSjTL/0jM8
Qw3Y3H97fH7f7/TDsxYWic/xmf3TXCHPC02Bdna8pOb8Zfsd3gnVQpHu8BxopELBvd3Q7uutUAWL
HDqpzO1zOupZTxTJ5JOqUha9BQ8LQtciMa3MRPXkpWEmNfijBUDzvbXDJJwW41d/5M47F+PD8hgd
uUdDGxKLrUarFl814ODN5wWVyM/r5xIjNwUE3S/SpvD7IGtIq/vSeg2jNUUTDTMQT75wgkN2fVxZ
AV/QDFgWncabBg95bkozBWkCK3ZRBkLwnY1FIEDX7FcN/0+Ro1A6oivcg6GdXwjQIVHWe8bBQUHT
Qmti5bWa00+8razVlesNVVSQmP7B6nqQhuEA0D2dofNj9OahEZDfg+JpwVbisuyM1jk+PRFMl3hS
0+uBysqmVOA9SUkpDn1zRFr8T7bUBhOBUisFwijId6ayRngRfnXl7pNY0SJF/BWPTazYAvPMffLT
m/nLApXRVK27x+LYK79JynQ93weVhmLJIkK+WgZRct21QgAB11S3Ai0VhNlUZlhKtSYY0XyOEB+3
I6fNOljBi8NwFVUnIvkgbeRFhIJB3XKUw1Osb9+KoU4SM7ccq2d6MU144bquu3HY6wgzVsTm15xy
/IERyo4KpkhWSRcDcy5iiJMfCQponUpfSqHVhshwaFZvNaBJkvkdAZzMVsDg7r5GzDq7Az0EnVaH
n3eSPMU1xyID3Pak2z0VrQ0nLhNsXELcrRy4ISMdSv8xWPsWiJUr6jprV+x95GMLU9t/KEGjE9pX
KMZuVkuz1IL1bhaXCwzLjzuwcQ6guLl4KdbCl6d/PiuuXQtT0ngIh7yFIXUBTSybGj0U8CqzYWjw
mJUu6UgFnII+C0iTqFyrFx+LGgBk/Qu4fLDuuimzsWzoQYH/kxzr3fAxyUE2Q9ld2OPoycxaQBT+
76pkNhXWbXOla5Rh+rwohyrZveujR0NF3yS5wcQ/atofV1tpIIZFq7vazIGypTu/NQpMlh8OUnzB
1ZTgkthus+ySH6Yhp0sXCy2cwCKRXxQePz5Dp23WsgGCAdmtyORu+ZqIhkk+jggOZDTSLumalXrD
NwD6wTpQTcMbIP5QvSS3wsDuE7R3Jd6mGIueeP9tWz5hcwkdIcDw3kNw5zH+pxua2rVmLZVkRAc9
+62sz7I8xlpjqc2hVFAxIlMSa5hbk0fwb7CZWxER6nq/ydHDuZk+NcQm2iHDNdZWGu0UTVEMp+eV
uX1ZfLs+g1fm1TY/B0YRdS/m5itzI4mOgVM/WImhauqlRymilVmwu6YS6hMDp6HhI3fh7d2t15K8
PVBXQRqEroKlxJ1QbjpG0ugCUirHWmeJt1dijaa0nzJth19HgqF7FTONPBSrwt0XqOvgCo3XGPTE
OM5j0ZKohIltuK+GoI5BIN9Ag3ejHN9PDNEqVI2HJ0d92dptY1DeV07MOm6h6wrkslNrS+5WIgrd
shkdGI5OKCi0xl/BTQjLQKmasiF/bVFAA6Gtv3OXETsEaubwBwYF92RGrW6lA4eEX47/Ja3FnF1T
PccOuyXiSGkL0hhYO195Ff3gejlF80Dhx84X2FyD+V8c6txIXiS7NinYA8osE2gMvpFHQvrnT++3
3F97aiKKVO3EGnKPoh3faXlhRnNfk4bVDobg2g/VeLgjqkOOIkc/nvZ56LG1yPVxcAARp1e6W17L
6SQq3UgADE8XQJx+AkXHB4169F0lSv7EaYPIzimbXCb/BW/VPR42UcVSsdG8kfBL6SVmKr2ZIgFm
TqwSKhboraNUNbdfJrpAnmDt2NMpsk87xa/+8K5s2JA2UpRjbf8pTF78mlvcZcwzHKzfqHsZWNyo
PomcM0/lCnfakrL8a+fXZhJpPRd0eq9lH/SyyqOZi29DPPQvM46hodfM6FVzRCKxkUnpc48HKZM9
ksRVS7qg9odamINWRluT296zHBbL+GNfWaqeK7kxYyBPIUkzGo6TGXdhE+Jcz00J3Et8J5iVtms9
PAb6g/HJ91cTJTgnOvBQyA+z5amTx4FsEJ/+Jyp9+LqLhOYkdbnuH7ueoSaqxHJ2QLN1O/TP5kTo
hThOeWBvj4beRyl0E6HdjThpg4bM8dg9FV9vxv5pdIQId1cG+URH3g8ds8EGpSrgkdsLSxm0sYpK
etqFA0ukeSApR/QoxyO8TCGB+gGEAAX+Ud+jQ0XiX0FWWqsoh5M92Lx0GBOc7K8JgLIX1imrWpuY
zt4n4rqP8zKslRnVV685ZNBlf9K10kH6fPGQR8jo+FVdGVdP90SiTxszPTdF+it7ZDzIXRia0Co5
92Cw8wp1XSh111F2ax/TCS+bVrKLxEQnzZCP81u1x+30t3u8zW9Irv2nTDlE1tk/Gj1kOQaY/sPu
ebKnUeQrpG5iAet6Sj5KZ3Svb2NnqcEV4+EJ3aBunDCPe672cAUCidvtjx6w5CrHnFDCwSwPG9BY
A3+5Muk9c+ICCRi10dYRIq2f+TyG9vUm0mgSduN1DWqKTKSINOYoer+wno08DBvz+VWmQw7n366T
5myn13gMRVB8HoLoByHtnC7SPnlp23xTJxWIwoQcV/MicstwIbmQ1JTdvwdsx/MKJ77Q/YaDsVtu
bRTJcx1dCqTjlXljx3avrTvj33khi7bzPt/aZcMI6KM1DRzffgaVwvKqau0//7OsiNawGIHcq//W
bupnVT6QidUnZtRnjOrFLArs1lZ4BlVxT4B/evcxxIKLnfCDDite1AKQjD9Eh7qL2+8D+Bysnw6z
fBhqXac2eAqrdTH0LBysnMD6MmTj9ZfEoSiBAjr5whUsRhy1gn7NDqI2N0BItwN5fG0uNNP9+Elp
5jLG5rD0SOelq8F2RMoi07/03j5ijZb/T2aZjrwRkvD2nJudXAw8jy513Hy7XtGTbG+QGgFu/imD
WQjuWKSODF66Cw4IbSTinWMbK1iFiTNomIiF2BfANEnhWG9MX1Ba6RuG6U11iFiQckD91l+MW1R2
HLMWB/VOutp9XLJU3ZYRwSl7degQeZQnQlCGST1zV0jzeKcpMx0WICHI9bdQwUgmqLDM5TrWu8Ds
90U3hF0k9yzUXxNowBwuyZ+1NceiIdYrPUYVOJJp6jZW4bkCVTwWdof9FhPvXzZHjINdTtfrHvft
7TaImzPqwKBBFDLFwsxXQIlz4TlFU9zuFwkimcTW/GBcF8676bO5UnasTCYxygOj8YIS3TOZErTs
EtTGdqAJCk0cYlG4rjChaynuRIpC60zM7KDJVSKZawpI5WJsRKQ7caoQJZHZ1JP4Do1ZNFLUHcCJ
7B2einQHmUtOmvVbsE2o9YZqYrQvaj/D0BuZli5XneFWlzHtqS076cQ1aLhaEjsfk3xg8QglfmzM
9fXzrU/bQpO8rSLZxL8ts0oh2JkhcjB7LktVhGxpWfklWU4fsv1LcMCL1XMr+zXJJAdZhKJOktXF
CrlQRDnQfrC/ceIYuvQuLnw/6GSif5HENUfzwIWEo72W1RU68VP+MDJ32AdtQNYk/sf0K8napQCd
jVNUdMGmxVvsPzHWCqoP1Xqj0v6smG5gNmVjNdCEnNtUZMsUzpoUQT/r9qCA/+mUIeG/GpVWgPbH
lIvbezCIm3/ac4olqKc4viAZTeo0zrMiW6n/k7eB++zo6VgD0NRGWwDIgk/U301P7DzJPLeHrnGF
lUEoxj6BKiHJkkDMRE8jetgiiMz7RP1F6AEwkIkWBIHlZNBMUBTHrCLYgiRmi0Luk3hMXZlp8TRY
hH32e3Gc+VkH5UGFxJdkWtHM669Vgw8bOLYyslknsC0zzkA4YXz88zhIElgbuy9YF8ucu68c9eMU
PlwHvty9LcpdaLPOW7MW3zMHYZ7rKg780lbsmwWQoSmZ+23wq29Qp/0Fq5Lr5C9lBhae8Ip3G9/6
tUqy4P0KuyyV79WxzEVKNGSPEbZIixwuhb4z1YIlZYMmu7vLLoC4LFNsWNExvjvpPCIdmebd3xm0
P0+wLL5RC91L8vBr1PYsF3/JKdmZIsw3Xp6mrXsE4VYOitQxF69CwRRq8Md6MwEmC8VohLoTgTCk
2zsqaQmfEfXvCM7rfu3dfrtgZ1DqpvBGxqjWgABT4PReKQO/rk/Wn7PWW1BjoL5T6n/Yb0jrXfUM
b7zstRp9hDlLOMoKaQ9ylEngXfSvD88Ft2ntM1r8PTtrciROsnFTYQBW7WKRAxoXOOtxjClO8oer
Odrs2j2r6PEnZGh17OwXOIxQDntNbj0rEtJ5S4HJna0DZGILyLFKGPQpe7Gmr9Mjv88n6TMcjcch
Y+1CpfP1G4BTVjzasIo0G7kb76UlhtdnF/CI3I3Ipr6nhpEYCq0jusQE/rZn3XPXiaORI4kuKsXV
FaWDmskq6h0NsFyjsG2Y8NqiTyVdDYvDhg2owrI43r0K9jHKa3FJmlX7EXFmHBeJmMgUj/8k4pv7
3Td3dY+cIyWfhbLGQv5rJMMww+XfLMTfE9faf2gXq9Tg4pg5cdT5+pLSY+SCCIg5yxnQhfmEvX1X
jdfst7DGUvtcUacESkdRb5lOvY9QHWNYDpgzYmjcrC+4pednNEgBhAfYydnqsQYEracUkL8J3mpz
FXcAzzHhPLliIfXGuF+x6bCzCaXYR6v4ji5ZP1cenAJyuE5/jJqNMO64DTwHDVnmJ4oBSwYv6j6O
+XhFFz6K3q71Ly9fV0dGGB+t+sVb8pv/Gtn3hO4meX2+DK11vY+icCX1GOqeytKpXUeD3VDYz3wN
QQMVGWSmLlUR/y3kv4Nr1WZ9GMAGZsJ0izzw1Ff63SKGbTqWniEuIAtkmVG6CK/YnN/KPaxA/0eT
9yCnnCf+M/J4kkAVjPcbN8/lEj+nNz4vC4UFBldBreZNfy6uVyaSfDxEZK3AjBC9zhTYTbYigvK7
r6NFHcBWySIrY2DJ6uehwl9ciiuWhGtD4sLSiqPIV+t+ANrHgpppQ69j+zb4D1IJey+VzlfwFswc
hth8clqJsSdH0f4Fyz2dPsXzuvxLN51UH0r1JdvuV7gmAWcUj+B/ft46mmVs1MjW5Xl1b06Vqj84
CLFBuBUCg5JyQgZ7FEVMMLs1AsH4SdIJI1z4aduz8XB4P3T6qGYuDQqdgrBSgGWgvf5yBbLSRroq
vebCex6sCg0OzNI0cr/Tha2rNIsuc92ZdXFzpv3q7t/B4l7zlS2oALMmPl+IzMboovkWR5zlg3+b
tPwiQ9DXckyJXok+Q+DW79rrp+GAywZZmDJ4hPG18ZYmprO58gDG8Kha6YXbY8pmzmauCRAcJiPr
ROWWbgpa2dV7tFuS2OHgXMt1lLc1Yzh44uUBdlMPJUjF5GNJiw1pcL1LOx5yVLBIi5HJ5rqGp5eT
G5P12Exb69y16A+kyLo1OZuuwsvp23WYV8t65JJb7XEG9U9orpOVjMfu9LqmRQ4YSJkGMTXn8jYS
oPK8Eqwj9BXBvEr1lOWOh3ehWmgioiUj08VPf1ddxYe4GEajGtzZbOApQ6NzLQA5AgTlYotE3Tub
vQkH4K6wcJRZlTIQnJ+jwrKR/p374urnjaiKOo3MLQr/pExKVXUG/y0eJH1Vi02RkZQgWBJYPB0y
ByMSkHi3W3HmCl5gAUMmCMwTam170CDFVcz7xWqcNyD22pfh83IEp3ogZfL06vMdq6OcHdsOshHT
JGV9LzfcaeDfq+bLiT3hBtV3rdtesGiMp+GYeClcblOUVzNe5NPCzb4wBz7xj93M6+Qn0QIkGeZ6
NKB9qecItVXOC0ACxM/QLzVkQ4J/591ykINMvl7yAJLAJMp3MUt4xJ1h1LA+aNc4YbfRhUntRLbI
BxcXK6E2wxB48Q1Tso/ofURajKGdoIahEj0Dzk1VgXodNimCE5NBQsOOymvJUDLNP+3kI+JcC9PJ
r0VHrx/QlFnXLmdULbjggNhPLYU3uCa0GRgnEWObm0FbmhhyWml9AseaxZiNof6iRjB854dZszVi
xJr1MscK3VBQMfXIW6KJPIetRQKnax37cQYJXsbAnvzSqjKERwavaEJ0zgzU0PnAXAIJ3Nw/GE6h
owVEawb1MQCXnhMAzptKh0go34frbAFGTZGp4XRN9uCbSEPjWIKWrUZloNS2RNkFc3AP/XDL3zMr
hlO9ALbFOgl/d5QbHSSbNYpGI/bNnyN5EZqnppIbiKGn52mrmuh3SBe9oQiZEaA421MjIrCR95L2
rfWNjV9IIZ8spal37IJMdWVkdiMfnaRkY/55OtuBqMltg1/9EiBSHfY4pkTHqmp47lmz3jEvPNNH
R7BE6wHLCIucE72QousrXubQGhXbmoKZRP1WVyZ/ArhPsRIURdejEgRfoLk8NxUn8kFbeXGOjC7F
dsaDOKzE6JmasCW50J15Ncp58SQU2jfFUtUV4XGmLI46opyt9AHsZ5FoLKRMKyxO6hRzUliUCm2D
A3khll784QbygPww3zRVpqCT2CUA6xRr5ekdrlC9ivlNDjOeymeDVYAxq6utcU7L/U1DKb4+3guw
lpDSOED06tSLnieiwqc2u4160gfalLyUQxtv36DHnUmMzd0ve1wRB5FvL/E6hQl3gGA7JxlHcKWJ
O788z1ZIX/vMa+AUwMku8xqORtFmmXpT+tyZBKWcTb8csDA1XRtYfYwS++tSwmP3WpJpWhffz+EP
ff2YBio/PbnPMI6xJLSoGo3x3PC0+rH2Ywy1v4RKQgf9UcEtral/n20Xw4U3dAaOAqgJBNKX/CaX
iGKAfKEPXSdiFt/jifHVWCzgb/sgpMWv+376/SSbpLB6n5yghQpBe2zFSSwaAi8tA23PqCz4DPWl
fmbpXr4z9dU5zziJSgSl2c3L01r6JhVU1RhuapWh9KMgWehRd2S4+QnVudQU55r/fmgONbvuhpq9
Gj7qKJb2XGFUERrOP79R0z6nERObYE0RM1JPSwwgZmpCKBSvsLsakExP3InG9c1wJTvzM5A7sdZt
WqytjGDzKAlb9JX6aa1fbBZXtMUPN5HHqhaUhkpKxz/YMkoFayFFVsalU/dzU1uBbiQ5uKbrLOuN
RBxiocle1Wy28zQ+3rB1sisdzc9K5DAk9vN/1aXmoCSp90ucV4wQrirbeudwSWg7bclQJtGofVUk
NFZfakbSlLZiC9GpZC1NuNe6FSqSme2JBCUIeRUXO9jJwsUAk0+lG4JGr+GCROuH7Vd6xUw/iait
DrjkPVXN1hGE0nIhagaOQPxATpm7gVT/Qk687SRf9haGPIGUYnqMHTo7omj5wPFXrcNeKIO71aFQ
G2oP78++wm6IID+aidhy/dSJ4zwEH7t0dHxzFoUwGgbgbAsuLg4m2eZHQ9+PNS/Hx0/Q1fWQBXMQ
jb43IwVv1r9/qWyADs2SdpejpHqyTk08M18U0UhHgbcvWzNsDoa/fEx/2VIgwABumRmujKhKMj59
BwTHx6PLHJSEmya3nEpfkBKd2oOflLUdVhWOJkVSylSzhDlwtI0LRVKJynsplBc0rAn0luHMYGAn
y2xankwXWmcuTKeXQ4yj//p2ZdHTGAFilNDGOF1BQ2wcu6BYb2x8fskKmM9Khay+pNKECS6PhlmY
oPtKdwGdWVl/7sJxH/GOcyFPzMDkXFHKS9Nsea4r/T2Cv6yzm+zwZ+YX2xpthlRy6pMyUz4aAnvb
Op6I8UQqzGlpsHhi5mSBAdxHND0S9ctwBw9zQKh6gq8NKqGTECsXKBJ2yjY7j1IB2sh4V0zKIaaX
qo7UnVqprLYjAa2BCUWv9sZDJNwmbsv6ktItUCWpGAQIeCeZdg/9YlGbqE0iSOgdtT5TNFQEppK9
i33jFkKZIFHnuSEgChKlUVmwUsSH4ihJwaRrMPaQjSb9ZUMyYSsrIzoeNTizMCO3W7YVwrp0IWW5
+ySXZC7p0+hyjYiz4U4gI6Jvu2ycALuU5E1IqTkFQ1wXbtdE24rnGXytFpGGRT8NBG6D+hXrRh6M
4cblgv7lEZNB6aDRevjAXcOhY1v4OewV5DFFyV3cnMIwqYyodQFs0lnFigSd1qt2jFejRNj+Rewp
Kk5bbpHLbtr4yBMKL85ofN5p+7IK/b8B0LgVMrmXvp0SFnxWUqrtUdN/9IzoaaYUShxFPODAHYKK
ifiRh5cxbpJ4Vh4YouLo5ZXDwF/WCu3w81GlN7JE8hoxHGArcttiZIwSYkrw/FOTeYsKwXNGeWmg
Y3BPQ1XNiKao8QcXTybQ5q18MnUZvJkM3qdGtiGteelXsdLo6A4SqgUhk8Iqsq4OTG7haf15Ao7S
zCMWGcBaOv++3AZPV0Z2LKf9efKeViM4h3mUG0W+IbqKFjN/0nMPdoSOrFfsQbAdoJ3nm5ftc33u
UZZoF2wKKTO0k3mjqMxR2X2f0xWRlZu5oOd9N09OrKm7TkMXgxmQ855OPafsZL5zJjD2MPJW/9NX
XgfeDJA+OUoR9TgRoJlU/6/YDs713txcBTQ2HM8vwymny2+Hhx1U8usqZWfYH9WbHykEzIeowKvp
j1hthyUKlodI+2DyOv9k9HOgAaVy2D6MmlsdQzpu5RVyGuMrHJT6auvb7amHQLTidAUrlsSekJaG
y9415HV4GEFqPxAiNubdAmZFb2anDN/07yY479+7T7LhvNApWHIEjsELAFV7dmxt+fwo6HVsVtI8
HzOa0Lt4rMiwTsz0zYioh0LI0gIMFitpGcLb8gJyFsIbz3YUJ+D8LfqYjv0xqmPFo/TrIzAzK7lA
KM2t4haE4fRfjv5qPGvvec+ijU9Pl13XhaFGcRSWkf7BKNqOXTO8T+oknFrdGfPvHqOkwhhur8Yq
T4pFwaWmta1XFvmG5pA+1DMxEy5MMifE1VuV5P4EW9utICOx8ZSWTa0BaN8iMJ35Ti2hwJHCBCOo
FytpRdBYygEan7gmoH3ERYEJ2G4YLLFrixAc0mwrHJtdEWXFxztiwkfwOrB4BcDtzsL1Gd/+NgkN
ecxV4kmabPM7QTl7fBetk5IJO3roMigXp8tKLcACjbau7h03S+nMeeRLNT22OgHSxBQMiyZ4lqux
2B3jTTH+lCZgyTqENRcFpTPpDxjYTyVzo8V4UN47Tpy9QUbQsp9eKgguaMZ7+txYCW+HPk34d/T4
QVNs0727uw6WzEz6v5wf1Nw6uj4Bj5gJTYG2+tWWX3/j+n2dv1qubu8IALt3yYQR+keCpDOzCom6
klyVikn5VOCKj5FT2rSz+wwb+dgE6HuQlmlbNtrwg4cKV/xTAYsSMCgtarQKZcwxgex+xode1sv4
XcmGkv2sKXBE4IcESIs166QzVHSZZqnMML5ZFM6xcAhOkmxoauneG4a26WlnrQjASsfwc6xaJ/Lu
5G22Kpgl7Caa39DVfFdULX51VC+0gtWHRzhxBzDexRuww8ADp7DeQBgH4G0RQ/DTZAwqz2za6f1g
vj6O8B32DD/uF9q7IoljZxmY8adSmy6aFsiOLMRONyRiX+VxwTlOUUd1va4orRe6mLgV9AHxESYC
yHWu/jSpkYvwjuyW0A5xwhfldf4OUx7HkbWThxeZg2iezyj/cJmkEb/pIWGJBKI0FqS7dXp/n/4O
M1UhiwWSYtcenW/kVwm9SNhpLVDKdQ6MpMQV4AW8bXGwiEDkXPE/p85rM/sfDsN6+/FGy3p8uR2R
hXngQhDiDrsfhIswiHI5Ymvl29/k1QxCgwcz/ky69eyUgUXThFNjJ0ILBF3+q+GWciK14DXNTC6f
h/D2mieEG98T2EQKnzuIF9gWf+xuxrMhwsy7AKjBz9HdnXylxLGz20XT0kg/w419aSSG0ndnIpUZ
oY69mydT+iJfHXy3QIa0y+79D/Ony/m9NEdHdhPQQvsml5Lxw3aEhrwxVTeWfXBHPVCCG/iZhoK5
S2fTAFpRZAk0BkXqylTi/Wk7P97lYtkrtE3DejETb8Hkk2/rrlUxmMiGp1VuAEBCI5aT3tvAXYNU
bWxijbYCHA1ysfB8yDPC/ABKFeVUcKkUNHs6Jazs7MBaA9smnCyS3Km77DJqMhNiEYU/EO3qfjrj
IRxKwHd4PUL1YL6Yzo9p0Dyj+JScTcRMdQny1FNVHvxk+IZxJR+isFhLpp2iP3WSZh097ryBLuPw
FmLrUc5Xc2i9X/sbDcU0ybO530Pdmg5jbEof89hbVrwVIJlIbSgYcVN3Z4tpELAHS8hb2VBvKzMt
LKRsvtWFDmEjabZAEAVVMgqM/z9r+hAVA13+GvSsuXFxSSdpQ99S/LdRFMtpUi7WZVbEID1RIRmL
nB+epXczfBlBmcEZhEaj+BR2DNfzf/+lwnXT22Imsy3MMnMxnqDufdTxpIv14ddPZt4b0frHmWGR
IunjZv+w16WRn3kUV8FI+kug2hjf2P6KLM9eRFmc4xr4lzeoIgMapaBRI1P6eiEwj9oD5vlmsPtq
5wtutUOKrweisekvrC1J5Y1JW2aQGgY71U+f+5Lq7yT7pzV03IwdLrH/+J6XKOLe66ikNL52KwOg
ojG2Drpt2GcInJvgE/SXGK/DOY4oSJgGMXknFodrVqk8GRzXkzq/gj/4Y2P/wnt8ZhFP58RQRc8N
wZhiX8eXXRLOL0p37g9nb1WbMAp7GWdHvhJkreHO9FaeIrSmq3p4+dEaSoERGcDxssw2vXm+BjEf
ZZrmSOiQ16Pyfe6+9Oe5twvOq9Ex9N3Nx/J44muxf8aFQsa0K8qsZe44W+fOO7jlAnRLLrAsi8U6
v24pdYemk3L9J06RYJxmDwH+KG8gHjYIlokjCXX2hViYcOzij2FTl0i+PSRS5hFNNP7Bj5SozLNj
4AWRfVbj+zCnwTEcZuiKCWJ0Zov4DUdxmVo7/mqxvkjNwjop5BP0t02NJIdq6UvTAHzdMOqqyZiB
dfb4IF2kIlLyuqIp1fn/BGePHAlozh65bnPFJk90j/sNv7/VW6pwoecbhZgpltT6IvmErGVsOco4
8d6U+qYfNWjVnhk8G43+7FDAXdRkSiUiI6w4fWAMua2K3hw+2Ncq9qShg5E60eBxhX9rBQw1ZCQY
OR8ztavfE+Q85nfZI9VqVki8YuEffjs0sVMBvp9pWR9+m3LS7fLETxIKLAaGVK6wXhBSjMWYNS0v
XHsyBInRP5UZDz6lf6eTxndlcLOmDJ4alX2EBUYkWwwnRjVWw7RqURI0JTHm3M4/id+FUnHUQV+/
OlKKTtNAyJz56+8o2otUi8pDMPtkCBBlmhbieNqRpGJO3vW5s13OHkksqIjC6l4FAZqCCPgF9DyE
8kjtM4aBA2o9fwiMuABND6PHprwR/3P0ioxSFI2o6JuocyrVpXR3voCuTJjiKswyJjkDMEopNZzO
LRuybx1pgZhkA68Vz4nRoD+VTRfpUdX1g2O+7kOeryuoYUa9BHKqESyH6C/wnhlbInqVh4COenVd
Qq2c+plm3MI1gc7TAeU0BMxxAjI8f63Yx5Oi/AvwAIPXyHWDs5RGoFYBP0Dd2Mnxavi/zo0AUUdI
TCDuMlmi4TP1/wEJRH1drHrMNBiSh8m+9a3SvldvuaqWzl+66tYhBUPiHRFhANwzWV5gT2AqJPCK
55eTROE1tzYvbyyJd4WPLev4QErVJOdBwbh+3AXk5Q+t+IeYKMmZBAlqYYbAF4h/+3xBNY959FZ3
yi4v1KRnaqedKTUaum+Pev1oG350ZmmjZ24/Q5NT5YyJxKzBzDLJ3Rn1JuJNwc9IGH4D4yTfl23I
aAPFWyKjgphNJR7j9YmeuQXz9LN5rQDBK4xwyHl903OoyORLyG2E9QxtrAg8JSn+p3mXaT6ktOOF
hWZchFxdffJ0ZSJk0KIneXxdP+BUEtC578c6WL1LNWfzZ+Pub2sNcUdo8yQR2GMR9R2zDqSxqMvn
KE+rUQJseBxIfuEfsvlRy2JcfJ37NrFaJOFyHe/JSIlnY/kt4jXVTVO72riLnxFfopkq5KfGt8vQ
0CGpmbejwBd9r5lF8WjgEXr4/jVmzn27U+lQzRo9ChHaW6KXmu8HQ51g9NdpgBLv2lsQHxUEnKND
sHqmRU4cKpLU2h81yTPTbg06lg6U+OwnU/6rBW5ap3kMlLoDBOxzV8WYmaYb6/HNEFWNxXopGqOo
EFFCt8ptB5FXaCaMQauSn/pZmNxjgVIcjF7RpCLux7drbluwcfHgJwRxykKMysIo52JdrfE8B2vw
TjuYbWuAcV6NnaaGLnjy4WIUa68+455TnpxCVtB/+hoaI5sdo5w71cAUDA/YXq060kPPGzu8/mp3
LL3XhEUzZfTbDEXl3Nm6h93paWccWmBK9y79qsAUms6OZu6B2XyaTiDLgMsgtGD4/yjPTJkLI1E1
/Bi6gwFHnJlYCUEVEOwgyQz4WY0Q+H+eufSp5reb/v3xmgR0naotPb9CwxP/PNC8j99NBen8DT71
KUkO3bvlcE6Q1ogQZVZTScV8vX5v58eURFWgRtmcWvCg94AwN6nfK7yN95K6yGfxiVWUyHWdI8Vv
Khs79zO3+RiO6tqdSvEoaWU1pYAHg3DBgPzQtVooYJLUM89A2K5piLiDK120hCyl1HsPV2eDo3pV
i3/4DNawb2FmlFkciexKBGokis7MaXjVpHvwEqjkuoN2+tXrlWEt2zETdoNtnudmb0MhqMHUiQ0W
wWIsePNhNJFIsto8ppnKuctd+u8n5UaYnGMAFiC7FW7A9OTFPIKLvhsGzobDiD3NJBMlvjM0vGtX
0FHBCQOU3S/uXCkxuOEgs4poTWQB2AHLJwxPPvGz3IYcM2DFKNGAFyjBkpOcplYtuf7bCkCiH/gB
g64ONSbMYEvmO70ahB0WjiLUvAyXRfldMe5voEiQJHIEP89Lvr46xyW3Wu+HfhCCTNhjKZ3pe9tK
iisFHN2E1NABeHAaJyAktjDV669GdlCUnXcFersilzhcUws+9Se2qsJKo2C5oqSuwzDdD8f+vEWl
8F5jnE36ow2xcEolO8l+zx+rCoTsO6F3X/8knuM2jTSKYA7RXjj/ukIStQ0ZW6/lbXNp3dK+XJ62
T3/PfzF8y3YDHvpG9BMjIkc4FayjszQZiN3523OzcxHf4XS2zkgTJ9GXSrqlng3OEhZspLQO9eXj
8kx09VEMOlffX6WfEAqid5OwraDi7Vx46qfUpo6xJGBfCf3ABjaeXMbUDQXLSXNODtOj/NnFhntg
G028+NdmIiFH68JK9D++tP7pkQRwzbpGVVGUxHXgyIbGUpuk+zYE+Xz4uOLf0pOdQl6dUjX8lYYL
NeVM2YzbpI40O9fgKJNfNyP2PrQmiS/b3rz456NFvJcNI9PSFaDsJbIVJCQisXmPj+KdzOXiVwk2
Y9VescgZMlQYvXa3MMfMw1Wa+BbwyHJvC73AgDPVuecZdrMZ7g/cPsCh9skMsi2FRscSr46UIbom
/DXNZcLPe5+lU9zt/dQUzhTIjUSt8mkCQrqOI8RhlQvCxvFhr8gy3ovcx2B7MwvlkHE2Y1Hkw3vZ
dus4norwoIw/6VgPQD7grlQcYr4Uk5tiv5Noe7rAw2LUGSYPf+evPCae8OtovEBv2k9HQQ6oCNdY
4iZWRtW2+FKGfY50TKF6uaRLVVjaqLLLEsNV1+AuGEAU4sxEKtqTbgr2USRtw8cynolke9tFMapN
kZK9lV2VvjhmqSRzmXVrLqPdPwrsdyDhPAT3SZ+5drYWVQ4kmbcqCeM1EqRNwCQz4yAvDKOICG6a
+mZKPymNsOdYGr1NZiGBw1p+Uhz1En0PPAhV++k7fqIa94yCFUA/uU/T8DpHZX0ITaQS9o+cyzR9
czXKMQCYJKlHXS9GuA2rLB+7g17TOF4SiMTTfQLz0os4mL+/llMQ/jvJPyfnQIJi7g3fP/TOQ0xs
RLYe5bRFC4dBVSmhKRAEPuC6kynvsxaXBfqUa8gCwJA3cev+2uyPor88lRj0rJHqxpbZPSIeMOGe
CvwgNT8ck7ZkQ6DfMjjIWF9TOKCYQb8TEWg3WXAF3WJV3jxW4RxHLb7QOKlb9dv1amx+CvgIjtw2
IoAgSxyTPvpLSwj4fCyC/zAGxFYdavII5do95CsHVDX5fVEETmBA/+zMhxPROWGb88/lmRqawOOt
RouRboL1XBzDGwlRlsbcfkjCh4HvtfI8+bmWT6IZlsrjUPQvPBfAdXRXXAAXiy2FxEnGFAN2NUXI
q4hYPVdHbgbQysc+Qta19sYD5sltjxGWlrGztIIk0HLW5RDeskSFNJUxh1ZbVwlWw2CJ8Py35S5L
0QNElIa4bbT0DHQedDD2o5oe2mK+1Qody3AO0gTmGQToBKjfCWkwBq/VaYOlKleMI8RUI2st+Qs1
Vf+Ri0EnSZRl4WcWC0FY2hvVUhgGFVFK47gHPQ8R88z+4L0KZcDZM4SJrGz80pe14mNrGOABkw23
9Gq5HxRgJEk2TPsQQwwpAjfIiwwGWeke6qBnhXhGWT8jmgkBpbE4+1187fIvNU2d10+DV6I5C9qm
e2KPqiRRM7rDJMqz030ptxuIW1bRi0dJJvTIOpAcwdtPosd8dp1fW3bR86UHADcrQF6RUkT9Zauc
c8/nPxtCkOVhSq1+Sl77mC+iCKrgdZasD0ZpyKtd4lzxvX7HA9o8SZCstiuf0yqNFpo6Msl8RySN
cmnG30CFn6jngP0g70Yx47yMX3jHIrA/7uBNDd64cGY/uQM5EMqOK5FOtAQSluILFlqxiDJ2mtZy
pf0BUS0lOxiGC+24gK8RAixEloj/mBsHUdx6/jPUkMzFcQot9+NntDDEQaw1gFTFblnfyL/Zv/ki
61iiFZKHO5SKVrO6Q3S2bMFnDwdEYeUMm4PDdH8SgBPgJLwVmr2HysxvyrKGYHPbUpOddzWwrgvX
BL7+fTEV4gWaocly337xNJjbWtqiHAr0rK/qg6xs+ZiuNcWyNiJVVlRde67S48jlSiW+sVGfU1Zo
F5kxfxmugv/b8hJbDfICwk1DG7wgaO4KtreWAujq+EsQKQg1g3R320+BS5CPEFIXRZSh7odKMqky
vb3r4cr7IpDAuBaFgX8pPi2m8rrDNGqw/kss2KnwB+BMcRXDhfjBfQbag7T+w5CfYz7FzAIl65VX
g1umBzSbuwnN+d+e22fdGhJDh1b3DWPpqqvuu3PKp4wQmwd87JN7mjdjlpfzc7yqHKd1/W7XhsQs
1cwmyptimG5rtCAuvKd4QMqRH/YdjiD3LnNROcaV0Lm7mh4MhgLut0+DyDkC8qJOIo2TWkOlCxMx
QRfaW9zQEwds2FaKR1gKj9wbkZoLwv+9Tp8G66aFCGzk5vAQG5wVJ8yb/ev+PTRyuUQClgkPdVjo
9OMQD3q2CytNnqdiaHUOkQiJBqjBv0dhVz7jvs/WMQwXO+noR1ZlKXws8LPNYvty8Pfb66NhnbJX
kg9a8r0wjn0V3BU6wefa8yjEfDPcFSs80AIwepEBjVp7vKXPr8IGY2vNiZ30zZ+ueIrcgO78iSyl
md32ESmNY8qTt9b1mxbRW/4Axle3+1ndT6Ke+gD/dBzHSxrTxDdXBF+P+s2nMnR0GXTxKCqo+/QM
wuRWclvjgQHu2Z3Io/jrNLo9nu/TrxXeZjTYI3h5oOqYE3aFtRDW0RBDRNVkUQ/aqoPCxq87GfHZ
MLT1WMafTSi1m7z1DZxn0ElCC6t+yUaO6E5ZttEi10OcoBTMuLoGGpeTDYR28r9TlHsTIGDJw+3T
ArPQ6/8b8dxi54uEnQev/6zpk8Iwg/etpNuBPoPgRQNmj/8Ka2/zjJFP//lQZnqFvUUpTLaRav04
US4m8T6VSRcllGHnmvWyS3OcCMvfKuI9cmICeU7vJWL5qX6UbzSFvbGdC7DOGARlYCSSQX5CX+XP
LkKpj48Yw9lcCw/smFA6a2ETAqG9/d3g3es3Lo++2vCjOAAb+2IABuX1/iMAVmeKDGFegvxubzfE
WhYU6q5dRDXyr68yknS9wW5JX0EBul2cqFKPfOv8gN6poylYDxDRlL/0uKWUdf1ALpD55+v3XveZ
9TdIhSVU9m/xoLtXvgNRsZZH2oX2nDzBQEH+IAW6x+UkZbPTNQ85EWDhzro4hJcq0ZYX+lAJqIIG
C0wYgz4kc7RbdHIatdNSoHqxaWcIACxTbgEQegBMkJ+VyfJyrkicOd5/vDiu7Pe5T/TSZ34JC55M
pJlCAO4mhWvE1zBfbkUP1+wVwdCVS3z//bCFoFqi+7Veq1LlKv+cOdIAF1DBcfs+wkf9Exmwz/en
JYih+DfRQE6A55pJyiOYGIUF6aEs/bA+GfzHwBUafIxshYaHEfZXEHhEZUo8+SH1v6PfQooV1gd8
l8Nj4o25cZgeMpuFwXWkPJcB8H6Kl0asKBq49xD6uNHLPoycXYoTRCoczXpTKT8LiLc4pY7rpVRL
KOJ/ck84w65/U+lQ1iq97GI9RrLER7iQYKKYQ8f0OJeYne08JYrlFiP23xmtUFxexbvQLNanDeQ0
15OXE2XRcF9v2v5Ys4yb/A6joSSCUkSPvzPOoNmemkFmznMG9+dSRyb3Pwv3ZjJXj7gepKXoKbcj
Jw2e56hUS+iExHkPjI8XWNVNafAVyW30dcZLk8TqdulsMJOURF0ALY1m9TzvltIEcCFnzv+pSkTV
ePb2CA36mwtoKksrTVYHMOFex6GxJINQgZJ9Rdo3s6M4O2j0lqoj4H7xlqkT2pNIOLnHWtNRf6dm
xob010I3F4DEVG0QHCNVbYN7tab0+4BT1NGiy8B9imskgqacqWw1FN2+TcTRUA2O1AGmW+NEaW3P
2Rwflgcbf9tdNcNUtTOFCSqDks9iLp0BNEcFQ5cGrxPfqpm4wX19Wq+DqvM9gFn5vFK4DtpKlDSW
x7xTDjpM1GIHxo69nB1jhz4O0MJ5xo/kTHW8QxIpNkSkPvN4ala3jbo1aCenqf4+Wgf+T7RVBf9z
7dFK3HISiRX2QUDbZKMixy4y6E2uaHfrmEapQdIy18Rs9/BFTaSFembw0RH7nEzp08/Zx+0VauyA
6funWIUhiXUFsQHoVjxIjHY2LroeBGv4NnFWyxmAhzkEDLQP5mCfFkh3+2CxzaSssWWj3oPn26PR
pLAD5wiG5lB7xrw/sZup9HUTX58tSMTIIoJDb3zHKMh3M8q8nJQ5UncrN71XQLO0yiOIy9J7RjZ4
NHCnDC4PAdayEve2pIE8vS79PW7F2SHiZG6kndtocav2J5Ck3t7C7PvKHFwwcOoj8KstOSTZH8g+
W+9tHKfe1/2H/fUa4hAH8V2IczGExokpD7wgCVSAd6vjp569GFmwAB8C++Fj4eJGD6icfLKgxIu3
3Xc+UrhAlqND9dkVyEK/+wpESILCQwK70r70Sbk6jXT+tsDZMOjqr8nbjQFmLhPXaZArYXm8NJ/U
OlK9pOWwlPivxf4zdnAtGS8w93Z6MG5blMUW56pZ4Q8VSJhQN89Hd2Wk1H1cbxtcuqRpQcHwrDuM
t3ZVCIQHX0FZgNqwSk7OCe9cLQ1fsWEBo1Hv6541vCyDkmFS+dvFvKyAIMfAQ5kuJ/o4czsuP4T0
ErALs2bJPQw779FYRmhL2zwLAkpDrsh93l2B8buoYPRt7L/6cJlIpm8ALGG7IDd8w4ZjBqKppfsr
uG35zwZFRaSnISz+ooXQU03x2UEMPl4sL88bflqkriLV0VcF1m33mUM3nod8t4Zw7vl+gbnhHPUO
FdVzGIEt1IWLUd6ciFD9JDzSGq2zFonkOHWHzeILRzpMYRC2KBywDceiRka2RbiruTxMbxoyLc/B
YYYCkcX/l+px5cWmYX0QypKYBZeYO3928ddCkL0Xbhk0hqu5KpCVuKR5sjxcser7mlHxMA4Vy6q6
xHCEQQ18asYcQIrd6tv+CdotDxh3Qjn+xjfHMHFrOHYOetGT3oW9DCqaP0qx1jfP1DV1ad7LWpoV
I9k6HkQ0BkCzFMeQG+K8rqkm1bqYL66kL2cDYZZKkfjh636CQqUyUUcnUKtYFBsCjc/4snxG+/+L
sYDtz52o0zyG1HMfjDWHGYlRwgSr4fM+f7NpEK0rGa+ZrpbjO6SYO4wxcg7Y9WmFbor/d6dtiNa4
ywiRuLjvVAGGLFxn87/loghmOFfyU1Orz6nyunFc9MxpfNOyBGt132uOdW3i+LSSfHoTqBRfOyrG
8LV1jslivLNad6GDrV4t1ueY5ZVXUdXBjgQBSv25bmjKSBesqX5LAhIOreJqVggmRg3yCodcuFMb
8n+r6U3VtOZRexWWkhNqKfIWgoyj0/0slJKm+hgieo6aPFsk3vsltn5/gVfrxHWPLNGMrG5WmWpS
jey5QaC50SJ9gc9GPiy3SfVsvP5SbIXFvxEWBVZDTyDmNvvotzScfNLLGK7smGcrg5rysO2Ehlj9
igja91BNi8HXWhbD42DeYYH/IqUByaqHx0ckxCuebHhE8m8kWYd4GEOTy0Vq16DBKJQ4pGqXtKfC
33A0oLCaX5TiZgzdbKjXlujvu41RvUfqas903jsyx7Ec/YGtNKMpfC7gnmuThiFoUpm1FCCxPHya
xgYQQI0nogUTwjtF4uq/iN2U09TVbARDoU9KXLo+CQSgAntF2khvD68SxBP01XTw1LN3Kw/SikTd
VDV3Ar0MycSjW4f7sA6tPkZ8uYx7Pz6NlEWKLLBJsea8rW82F3FNtjp4vmBRpjjuGKW4v6OT4hS2
uJSGFtHUc0TX6zg/bJauG91rV5i71k/oCknCfynL9FrCaTAENh6Qig0T0BH8A3G9I6xK2I3RGrgL
bWhJ6ePV0NjWr8Pq+6SMGEKO83MIHi5saaJG3Ba0PgX+ceZuwnyKo0DSa8xmPvhyeZqJgsATb6UD
01+jyLv23YxcFKNzT3t9Vzb8Tt6qAine+gLmkomQVIci8J+wwdiRUYBZ8WFsXgQH7I5e7wmUJN5j
X6BQ+SdDnxE0u8JB85IL0qCk+Q7oifcqQqWTAMlgq1LsxaY+JKBwdZI9SqZfUxwOhGW813STpLUk
Ps/2DGlvfRwNogECVl8KTjZ8wW1qnYLyEe+yVJHkydJnTDMd9BtWrsGg08Pyw9LpTJIyjCm3uKhq
iG1LvKZkKbpky/M8hNtaYgDRQe7sLfYrhFyL9o9OP/DIeTFjRTDlyEv9Htu+sE4Dl8mRmvI2LGZo
9ZtXwxzvZqL600EYXbLiaTb7kSyJ3oRDCUk5LHLE3dJAAzHwgK1DdGwgSNgjew0d9RXc4UzP5llW
1lS5bARTEkmJbeByYgFo5gI1YELCKbPCUATR+QEXa9Ah5jvun1SNEzTKtC7efNzRmHAPCU/tWO5l
Yr3dbSRmRZFKnmuvhYWrEYU8+a5eqhBYB4ppMoj9z6FhaJUa75UTZ5fB4hNvfZOWlHRbQYpt1fud
GOk3zVqGGVoVv7Enkw/tBkn9PDcchlixAIgtCevLP2EDn1edzgRPDX2IU2c4BX7jfSI+2IXQslon
hMnaFCEo6T8p9pfG/lW9Kn1bYLbeMgrW16yNX48w2DIcY/hNhD2wWhsZs0afdml2FJgR6TufVXlD
8H3ncAG3ouaIUm4qbIyUrhrkXQFBguSYW5KS/zuO5UFltKLoYS0IegWleNmrptZRMe64G+uucjIu
ybqs+4SlloLjYrQZLsWlstn5tTRGj+0JfkO2YCxnc6n8BjjqM3FO6QSHQvJSV0jGPbtuYPio/QGq
7hMpAa1e5fsXV6oNXkeMaSXy5+vJqRyxP61LXMgyS7H5qAwRs/W746qxB4vsXPBO95yPU6o+Sv0u
JGOzAEGpAxSuaSGXfnC4/DMC4PZHaOeqf2Fo2xKo599eC9fR5OTSnmbJVsqDoh9VTjvEah9bEWAU
4ELoIblWjoNUrYcbdUumTSxvhce7Nrqoxidg0YyVjBE1/6zIRwrcyn4onQZ9gQ19MFUR1dNVrojK
SeWBum7fRyD7FX8qW44wNZKgpNULNlykE2aGdKFe9SZM2WCk+rWZ2feFRumfJ2E5nc/Nx7UX1gfv
t+2eXwA4IUraMHX/X2LusPV8R9oZ3kteu9tXl4PVORKYpp23S6cbM7ew9rM3w6umM2Qt+ng+Kjeg
GetC+AapYRDdPg5nySJYNuKWE7Z2lRN+d91DknNXcmQhuZbKyuFS2gsz3I9k1tyrgRtQ+6TzerQ+
KFzrnjBnMNcQkLC2LQAwW1X+lMkOYZNk01UBGF+lrw+VijRqcc66rZlp++0goLOd0imCD21uBhkF
FBDM/3s4BUhRCa4l+9B/nMO1keOhZ66AxGzvWYRPgiL4S1hPa7wKmhGs3yeMUolxEX45c/LxBa7K
LKm0zIdiNHCEYzzE/dW99sisEi2ZCFgx7a94tpvDQKmtmANp2CsbSiJA31w2M0GJfh9xkKKAK4Ju
5vPwhGtutW6DavW6sHOHaaQ3zUB8l+reikl5ugFMK+IdKaIxSDQGG5Uy2IH1u06YDqRw8oCG1LWx
DQwI8GUFjREasRJDr986bu4MUk/j6+91ZuuUDCcBgTiElU8gYaS/X8LWFovHlV5znLlKzz1/MBxW
0laMSdgsEP8tljQ4ODdnLrVIRZ7jc2XV6VQoCQAM+umIqbmcR68LzY90EYKm5xq2OxCP9il3rAsS
+ah69Q4JmmQEpbm2xr8wnrqjt8Nm/gZP7spTiqiCSyqviHLmuLAlsLOY8w+8hG3Qwsa6ZNVcjrOS
+r5JlOOfNO3LdHwG6HzHcXmsdtQTd8HT0lR9y8N0aOlMKxHAy1ZAPGB6FZAzM+hRaZMGm0J/z5pP
d7NByhg8RbwfIIY84uJ/6SKBgY/Sut4wKZ+c3EBapELNHbyAJqapfSFkpz5gS9qqDIrpurh+1x33
16kytZPMTF7LEX9WalKyFEbFajyu8Zqx/uJsfM/K6JuGbd5ssIQd2Ndq7ZcTeqncOsGjXn0drRgy
SFfqq6DcIMyqXw3mKuDXBC6P2yqEfwO07bvE6K974+r74T7+TWpTRoBuBzmEATqViamqduywndFN
8XsXbJ4vhGYdGugsjuG38njCiQvBOI6QKjZVwcNVySEpqyVRSpRkAsMndt3bTBEsVYQ6Ya57ptGW
LgYDZnopjk1FUImNUWIhfcNnfJQzQvh4/vsPJMjUwYfoHd5WgQhxVeg4Mu3rpSZOOcikzlIREnXt
zxUsGhHubIIl6PK81exSRQC2TrPk3TIjPuLiH4DNVeZnDHQwOq1dpq4bm4EiD8fzx0cucvUcpdT1
NldQYhqKBi5ZCPdacnYnTAPynL+42cMf9nsF/dxm4phQOGI4VqjS2NpMoFxyyMBhk+uyXfoPjUF3
aoPczuzL7lzxs1GvJaeevPHdKe8ZJSlVGY1bGY54hO2+nvJEEeUbPLyNjnnm3OG/CjGS3qweIyW6
Jlf7CAdNFcWnV9TYAt3UjH0idPBh4PHBM/4lT4bUJ1XbfeshYC4e7Xx+OavLSGsiMNE2avePppkq
X3X1jOsbaAvBvg/cfCiG37xy0ITPi9kIZaQIfXfCHnxAH/e2EtS+F7MDuFBDNlSr1P4xriWGyfMm
EJUyDIF1Ztyrhudw2rFDdjDulRvk+emHELzRNRp4xhFzxzW2kHlLWO5OkvXFs2zL4XDC1dMQnod3
TOpc2g3J6HDhFLITJfCo43ea8c6uhtMpfc0k7OOh8esTVAjT6JcbzHbzl6MB+22sY3ToVOqUQsWH
d2KgOl6NOnOgddSlkHpJmhGyf0covePRbatczW8aaRMchx33ggDx+QCXNDL2DIkOldZaofbSHf1a
82P5qcxSnlzjNXjBLRID8zcM3rYZzdrBQXtMLh7uGroeTCeWd0eQtWnMTgOQZCG2VEcjIJ6cTxsY
d8V1XgkmTBUTY6G7DWbNOVJ3NH9czOeKDYfnhYF1Qqz4OYCVaKm3rLiFqdGVGocMTN3HzsJPKczv
93cDg3LadtbqDdeEVqhI1UmY2ozCjVSkhTorl0KGGdxG1BcJb6OZm2DNWbTjQavoYKbShqMlSVlW
U64L39phQVNHwdJek5lyp8hhAt2ateRC7+v+SHKSWdiNoFe2CR/aco2PBjrwumY1f9ArRrkwk+jQ
ItVEgN9VEvdNkx1iGeRgMY6dVxfVBpjcSruV/KNZd3iUedFFIWR3k9DsmBa9AlYnUBjjbga3T77t
zpHxFRQ6nqyUa7YtHvcKOxazDC30Y9XIqwcMVSj5sd5MHtj1Mvi00GFMf2KVB4s5kp2snR5eDvqI
eoAuFfgqB3KfR+Cq8mGwC0zXa8wy5HgOeMR5aKMkYcwVnLx+rYhAzjNahDqHpxsmImiIE+9hyitU
xdx+fMpl8GEbOH7JhC9i7Ggih6vJl7ekwXXBoKkr9Lu9ZZzW0CmW+S7O139CDCnZ6XujULoiK9oa
AIFq4j844nX5nI8G4Yy8l+Hxunr1bo3GVFmCTPI4GyfFVV7LEKh36SjwfDrcT+wa+Yn5RU1mDg67
abMz2CqMvrF1YDfRu9mq0wrMpcoDLbYARy0HdoQOYMwvmtyutCpt73I5YbaxtnJBN+JTOUApUmkc
SE6Gv0w/B6G45hjGLhGCwP5ns81IbC5cA2H65YUTyBwwB6gv7Ks2ZNe3tLn8E8kP5dITt+BmLbbg
CRCi6v0RmXdmBOioeuNkYEbn/JKSaZrkWk7jKpstD/E1H+0Y1c68fRbdVAfP8J7PhuGhK8nnejmb
dLG6njcLq1YTD2a0mxshXiIUQXO13pRHXz9F+Oi280LIRnfA0GVzmZgz0oz/8GjgcHN4S4L8dK39
hjczw7qeTbGc7AK7S+ZnKkiwTcSVSueCyq9tc5fYnZ/us+shkLxbTfGFA6vRqmky1Ws0B42ZPKR1
MlclFJAAvi9L9Wnfpko9kge9h7xX7NcqBx39Mj1lX3FMStErwmeWC5+di0nsXBhg/zwXGcPifJxa
7ovQgW7DvGYTHdw2z4Uo3vuOl4ilFD5c0z2ZzZL15WvziPOsOsbeELDyZSSPHfkMhMts1bzjl06k
nfM7v3DCYLuthLVGG7V1/rOvLa9iKbz+tRpYooSf/eohpsh6BvNWo9ctE/eEAFmPkNGWIZt62nlS
mhGrL6HG3Xb1OmY+Rnbjjx2pFWnof6cm5EpqOKyLWGcGO3rMLbR30PIlJO+rEdKIuvx7FLQiBfAt
ajyk7ifP/9FocBKnvm4llrbo5RlT+GpcaxKwtB6EGN8Bi9+q0uSQB3bHbJ7tQ91Y07T/3FgcxC3t
nioHzfu3mhlCWEaCjgE11bYaRSJMOP2pl7jC2oIvc4kK5NP5clkkrZ+fvyjYQFRQXgILw0yNOzPv
Bovhwd6WYI7mJSaBfoulEn+4OESU4sDfDMWz2QU4tMsFwa7nFc0Wned/HobYbMeQa4WDU9HUXBli
zLakN6N4ipFyzJY/yAYQfIG45oku8psGrfQuC6JFytBmXUzTLZWFmPXUIcYF87vt5xE6d/5a9u1X
P4YZG4+dENrCkfifiNbkiXYctu0sSIE1ue2uKjFp3iGVlVWWRrwI5AwiFOThWEyiIWT/T/jEGJvC
jX40QZ+WyNXGq8dk+EbaAr32JB7XDfiGlZG+2/szz+RrrQHfOQKYUQl27RbOQvgozrpXIjGkCxSj
b9SSmXkfJPOEtzdLG6q9YI3LITVUJdvSVE6UwAuWcfiSbX/tyTeRefIhla4KSPJ5YORBGLplfY5K
Na6Kg5+NgMuPpnNyswK93bKi2ffljOUvraP3bJZr7jec6clOlqm5Eb1CaT7GlURGQdGGat2S7txZ
0b7OGA7afXyVAzZzGvU87FwHO+jCn7aSANzLIRPOBXjSGPLcHhk+Tn4OS9etv7rQB+gSljMwTCeh
KtqNEn7yamIgtSfiIU04hBLN3OpLkmSrMvBMdQ4MOS4/X/8RKkaxe18fN9Ro1alk3w309mijtSp4
MAVH9eSp7u+/d8QC3OoAsRe+wO2tGJp8v0iTAbnmsYDkf7TkOHu7th94MjFWQWbY6pTHqpmfXlZm
06tUn4GUOtEXRa5JK2m2IKfOVo9MUGSiMuuhpPxik3MJ1dhyl9OulvOdboyhtjxA6asFvSzcgaPq
X3mCV4N/dLqKmWsYUAHeKK/Aa6Kotb8p963YH1zwgibOJLcde4VFioqgm1pOxNu5XthoJx2p80ZO
BDBWZ47UOYakCIfTUU7cP+0MPTMTYj7LqxQ5YOWiZx0reb5xE5nHuYbY3bpzhBvHrvQ6AwDCmrVT
0YlpiR83Bz/ljAryf603rsWaPE9TsUrwWZNTiKo3/gkLPylnCLHTta31TjseqdGHTz/b5e3h9bOI
GyOQn3HcBrXA8uVkS9fJH1zG0kOSSq6C4JzbTitnpmv4uN73ZKxS/osKE/I7zDFZnIiUOBUSqUvY
8ouNREGqFBYG4zQ4G9Y69gIULWfOipyW8ukT7nLWVFfXNF9OkKKIRinQYj01Y+OBzDBGmO6X1Vfs
Hltr5YOk7bciKFpj0Xba4Rt0LojRCvGEoJpkfX34ZRHcQNr3juC6ijm+iGVoKQvpSeY7PRpFrYU1
Ulq9CyBhDkRUSSnCZ/RwJ5Nw+CANQqASHeBd9qxwlQkgjcS6dWBmMm7+arbK5JYtyby40atPKzTN
UMSBhj6i4R9eMUAtcSefo8qrfoO8AC6WU99PdRRMxql/Y0M2j4xfSTTdTrDAb40AwubQwy4ZkbLb
4z12Psm4UiAA9WgedB8ij5gLCRffG9Pb34bLPJ79T0mt2Yfz7MPY440mEw7iUiGRKlOrrDXtxGot
TZbar4IbP9wPZ9YnCdkUCghuse7ahCHnT5wLsvc5Wcm/YjFLWFcMovE9oJxteP1NJUe0ctn1B6kl
ynLkBxqwKEQzXxK20PFWd4vs2OyMduOV+fgrJLWLkDj56AM6LBsOF/P3LL6Lw2TXinbwwSabLcV7
Kgx3vLd2AWQDCGmmNBPybbLWkwFP4MM1gSL9yjQbVMZhGSaLcz7iKpHSmhfJye4haFPzlZr8IUdP
SweZdh6aMaeycZRm/N3A80L0uAdO/jkH3m6sZ1fz+TuR4EpxPiDpIHNhoxlf9xIZaJoaTRA3SpqG
P8H++CQesBfk6cEzJnGzifurwZme3JfxRTB/eienpb5M3HGIKWPNz/cZR9rexGh5V7fIhWtj28o2
GLhfNi5o4kKjnMkz/ZIIrMZJ+hwHkHRrSxkhMI36iBmSr1fw0u1NLQGrqEE+ZOJzgJaPMWfAy8M1
1woEO9+DMLwuaoVAVDuj0fKiir6sUdZs94qMEeP8f9ZVQPpEUmWeyI4DZxm0uKSgL8hCpucAFIRt
vLialg2q2Zve+ThzGm6DknaOjmYB2SKJVV+37muIXikIg8NChoR2MFFnWGav8PMzrRbbkGPJK+/+
cSw6KevDPhL0KppJdgKhn1sCuz+18/1Dp0THef8nFREfl0p2Nj2purTkH3L7JKvUGtxj1l9XLxI7
6yv5EMy/0h6KpQ2kQ6hHsw94e7SPMjxtEaf9a4v+/orsUmGW82Ch8ql832b297feKBPzeZ2CjV49
oWHRy3FbY3T3c3AspbRjGrYnAzsHe22P3q0K+bp3AQnIjH2xh+A/tL//+6omAPIQiefaSRWGGzqd
lQyWeHEcZ2NcDcz17ZGPVKAJW6c9t2ksYHW2honLw8BYAuJuU/pZ+YPYj7NdaEgmr235pkzTv7q8
RfvYL1151MBbml0fOz6T/JMrDe8JE/AgCOP89T3S7aba/05tZLGUYsXd28kNKw22Ww4d5teZs0Xc
zxnHHxz1fH5YzuqD3hgskBUf4d8n0xOowUUy/NYqlLjDJBiVyxmEmQEBIwEKHb8AmKOvF7Lp7/DB
QIUtmgGQszPyUpS4U/tZJnAIh0gTVlVkJU7u6rRk/h+F1ztefZqr7z+ls9Pwd6fBBiGSdOXrNNho
Mw1rGQWAsfiv8yEppYKKSVFxjexZPeDPByvEAq6D+02ALy7e2OCP2+/X6O20lOj0sS8z5f5Uu3pu
XjKvHTxaVxTstpJL5tuynxZZ6rbWwZLGgqtWdRsZFgez7ixS8u4mr+rZpplvbe/S676g3kQRYjSD
DHaIqhTbrBgQizxz+1bd+wviP3VqCz+IxPCUnrqp2mtUyLSdMYZ1g3/ePd791UNGCocrxa/dtVg9
rpn75UxBxQj9xf++yZEth3UlqB3BkPv1HhaJXIxOyaFRTarWclUsEyXDndHx/67/6NdA+knk+MlR
8mhfyjTx/vAI3JTCDNuk4ybIFo8Fy6qh4UAm6M9BQ9rfPVQgD4JpehnaOSEl8+vVhqDT8neYOEH1
Ukj7DUAqYDJ+IEKN8mi18fV2YLAHBXnSm3I63w1Pp+SlGmQcKlEnmF+LZxvSjZUMMhsVNjv5FUk2
AJKli5ZjFYhZY4Zd0UTbqmy/0gsQXnKfIrCexYZirYhZpMu4JnNZDdURWn+gc1+0DZqH9+gGhzgt
Zo2inBvhPeuJhQt83EsbHjxpLDMbrhuJgRbXesoOiIJ/1u5J1Ix8RoLt9iion8LVgD0LLoL/IZd8
IBE9vK44AbjHk/Qn/h5zByKhLeZCYPYw9PbRWN19hR3QHcNOxjYXyMwLZa+L4HAnSCzgh934XS/W
xlKq9Ol/5aR6n0yUGv7I2NlldqWTs6adltvbgBS172+SLuXjOu71/GpQO9IrqAVsridIXgJ8Oa72
N4gIR3Unjtwke/r1DN2IEqnVxZcu6ot3Qd7FaLxWd3N0w3ArSsyGlgXl6QaC0Z5QAn3e3EqG1TPG
VKpjJo0iMunlX4HD96zufdUyJDRdxJdv0gTQzdhBkrpdp/DM1DBaNNmJxNb+5q28WCKY98V5mZBh
HCJ7bVSVGI1Skn5e+DSb38SSfWet5ULPYbJcTwaoK9a3uhmv0gnk4RqBc2hTI6UEYWXeTGwQ+hke
2Dj5DhHeBD6ha8Mb0aOho7lmgsNZktMO2AFN83Yr4BfxMAjm7bjBYrmbDu2qgC8kMk3DoiSWmIdE
1VuCA3Mh4H/KfDGogx0wOSylRe5pej/Qay2R7Vvx3o/r0wI/1Si9w78TnZBVpbXpoJgaA7rptJgu
rwgHLaiJbFiVt+9MA7x5QatMJdkgUuic4qo4SMpxhtMVDgXqtYP0hah+YhtCt3gRMFD1is7As/5q
WCRk2ogVqvt34JRlZ2RMOrHP48+CAPc2GR1x03fsnTW5+Swo8tbcJfJq8nHAR0FCp0h28Nc8p4iW
0KN5VbrCY7AQMptgRC9JGc7+81dc4q0YP3dlXyltr6nEa9NkvVAuEK94xYhuKiRLpTsRAYzPU3W+
zhcwO3qiTGSbZIiauBUSY4HDHqmQIW2wceaq/GO1edYhD0cSESW+6f8BOX9gjywRuK2SHNhs+ILB
A5kF159+ysIlsJ66b8rGbZFtyUybQ+d4yQF53NG9Bjp62hRjmzUpTQ58oganrMtp7yVl8hPgJxg0
RPPTHRhLWD3I/Y32FDqAeeof1RTCCexK8mplSZHk3UNGf5k0lysAEVUNGwV3mEAP1BwYPkhDtSZN
Bo5zbbATLJoa79AzG0pETKKD62uWOn/+CfQUalgBpdrYdRkwes04u6u8XXWsjhjoObSoCKI7ffJu
lXe93vfKpv+ED/0gGhappaOdUjFKhcpFn+1qZH8SdcmCVYoOWa9BJcqyWTC//AjSQ3gjeUEuHkyZ
6Fvzgh4x/upyWaquvyD2tlQHGd4in0EEpUaAZdX+3c1Yxpqy+DU/fpvZLldw9FlyQbpOHGWHCwkQ
uysfA8AtJQXTz9ZtjTZqbN+/TwgviAKMYKxGYF4qDPcfNHGs/DtRUi0CR8D4PUBfe68fMPMkHkrC
EOxsT0JiDZ3UXMsXEk14cRoqT0DkRTLdpQM6s9zwakYbx9cLDe1NPuLzhjjPCOe/8aCk3RbsWy9I
EiDrMFyoQRb5JeS4GKYG/qLe1ceJpeHhah8d5qEO3XDKPOjsow7RxxXvuXzO5zz/ae9TEuICiqtN
6oitB83+sJr5lCQPHgWw1syYr3e20otigDPS7/CHwu5HwUqOODK0MLwpohfoPxdv2zSMAOBykQ4I
XNyxS0LZtTXaAya2BpsMGqjie4FT4JJ2xJqci4tpCfQvmGySzvTWIHNZNWB9s5n+fv+cX22SbWGR
dSWg9FhPXu8Un4EF4ujk7H6fqFUezObTfymSvZuS02//eKx+OnV4kf7NLnHX5juRn9zvXSOEzhxX
dl9VEjQr7ERqn0sG0k6lZ+MGNrImf2PSYK6Mf6x+qJrcSEKTinKuNOhVkFJLtjsJCzjFz1jLuQIZ
56khJLOg+S6enWRuG8OCHCR1d0WCq7I4oTmdOLBg83sulUzSsLGnpkzGcTjFuV5xtEpCTolERQJH
7EnMBALHqKzgTSfXIKKV1HA90osfw9g64lftHXJorLkidIqzWjIq+56k6IWgtqaIx4FqHRV9/kbV
uT5E06ciUVEDUkQCCDnK8rnHdaiudmajYdKA975uS9o+vjTmLN/QCHj4vvkL5ux4G9J0ba/Oy3Bq
FTYykVPMglIhudyoPTxWjGFQZE7Fgb8mz+ubCHuXQBUxUGihlJketUcVykGHnXhV48zo7eeIMzVD
dRiiphOASzvDdVZsm1nePU+4mITAAWzkzwq+g1NIAsktX2nN/MD6yESzsWLVVScgKe6I9yTT2GW5
Z+Pk5v7EUEBWMWaGlYx+MPEYUCCxrb6DPcAmEVPW7k/nZZOHYLpl2SKjocVkK5akKuvtFkkP//o+
sJvCNPsp/zH+8JlS70C3dFYrko21XuFScTV4qnhuLAKAfb0/IlE9EoE0vn0UCidaPbE5o/e25pxY
9O7dKnT7oNegPJEzEWXRflLLPvUmcE8grJVZ+lt5R4I2oS1GRZFyCBFAjYQl0OGifNcYKZBEIt7M
b499LO5td6Zva5KznhX6d75l0ZAg5/PFyWiATW0oL8LT6wUkmOwa9noLHSyfZFjRHdQyxeohBH8m
nqKnaPH65rIA2QUboiuOJcnXz3zRaOBKqB51qBnfDUi5CC16whTyWcZXweII0CP1JL7xuUt4JtVy
GFpvN7j8TWai9qif8J+nF3uvMLvUds5lgw+YQaeAUSa8UaSNWXDbYKkrL2B1X6lxzXa+A+FfpnXs
ZesHfxrZhYFcrsRGhHrlUVF/i6cZE5yAdkCifmNMG2vNT3fLwLz/ge3fwXfwkMEBu9PDaZQGlr3G
DA7xg85WIzFRp+SOrXgfp/jI/b+4IIc8MIUpmEX9s7aeq3tbG+kiFEBVyWbCJtBLGkLvK5nhX8K6
BTjGoYYuxV88lWZrKsQ/SwmAUZDPDPmWTg6WURuBUvvzkGIXHJgj3C//eiTV933bL87LuwDPoNtg
VJcMDUYUcs0sTPpwVLoMsuOszbPJNcqmViTCN9hpaNTBfLkyVg3MpoDXw/49kJkeuTte2YPqHOxY
iMZswD8RK8c2JPqpRJ8QAApM4+3kL1z5nfX8PUZgiWrnk9gxw+klUENg4XPvfEZzFLGpyQXMYOz8
jLn3EP4WgyNO+KyW957U8JnmqoyavwKr4c1rwIJEqqFciE/oMWa6WVzsIP+doMbwolLgglyP/LAt
cN5Dyzjwz0R5yqCt8BkwcpHQKv8LnL384TiTGWp0Bv0LZ/nqOYMLdB86y1vvn4svnCAVBIqNku4f
KkDO2MLDhsxkzvA/6jt8WtpmLP53+zfpao7L+6iBgP1iAVN+IXE32e9EsvwqjmMcJQoLwEUyT7ZO
wP/Wy4TQOXEGUrEXBZyZ03N5EmVlZUUg4eeAHHfONTAdDW0uuiq/mqrNBLodcqwk65lCQ4tBktG2
RR1SYMlC27+twO0ffmEx8N9rU/+pUAhmwn4HT3MZQoqKmU97nFe/SO5Tnyu2IBeKHLZPwT5UcgEK
oAinTaOSy/n8/nVm0VcjWBmC9mFmUIoFC7Uhk8zDXmWbwUmnmCiM2BblgSedsH9K9CK53VDqDl42
0t2/pNiq5xaj4y7hVF3PDDqVMoZv8Rm4e2HllB3awpDDVQ+Mua209PsOmODxC+G+VfPVDT4O6clJ
SyD/Q0tmiiZDY4afAC5R/z03ZhPYt9A4WRsPwj1UPxv//md1Lo+yaREj8Dp42v0JkR8wmu6MCgdo
ploI3jPBmiVD+c5c32s5/2LjmQx0xfD8qXaZR8IFrxgY2S43hy1FpGMOOxalMT3DxJ4N6jP5M1Hh
lxcEfN2Vwgm1XBFd6Euu69xLq3a/D0TS9R02BCJaPvC0acpTyYjFxIiDtIFDtu7vPsdqtOVxbtLD
B6WbKt5hGANbmNJzcfyEaQqPdQUCAvabfk0ZOqKuT5Gjb114ldDg2O+h+kndVf8ZoZ14ksJSdq/6
YiB5xka+BpdI8cyd1I6PndBkXzuHywNnHC9lqwu0IwMaBZ7oHyEzLEk9VIlWr/DsZ6dG3vFKC5fe
gKTv1P/AvHBg3Jk8HJtfRT75bevdKTZqx2j1zcYHEAriIo3y1VVNs78tzt4FWfqyJLsHlDJb5WQ8
rv7hB+gbmKyO7HvnhYk4MiToN2FON47yO7iMI35F7A3fQ7eTYcveE9uiMIMul9SOwJ9nbDczVmtN
q4t4esq8cXuzjJU2fJmdapNjAtvwlThU34WWhmyz9DqmowxLXpxSdI3VtFyd5LocCp2lIvpi5b3y
PZubV6qIwGRvaCq2YlIUyyclL1bPB8j0OGvegcRNnUFK7zvH553ydtOzGvEH2GmXGzQz8dlPXYtT
nJNqCRO+r5EptCyndUfAqFtjn97sX4A2ISh/8CS6BNlbHG44u3+FzxoThhFyBfsq15vvMTinzMGC
n/KtPFkyGCzZinKcmNnCuHoGl8OjGCkn8C9R11kb3ndU8kSrOJySxL6woRe4SuhZhS/cyPgf8L9P
EABoWV3ui39ZfDLeLW6mYjA/OuGyq8y0RtIj67AlMtdUz/N6NoHXP7H//n4q3LYrFMEZYC8mwb4w
bAChH6x63kiPBZZxcPDpyCEWjAKcanHC9HrfO2ZThqGEtUnYk1M/lCnlEOB85x6yuvgxWb11XCyb
354BZYfwatxs7cnDHACl24leAZ5ZwhQ+0ZeiR5JqenxUFy7z1rwP0bhLKbUiZ5U4+0gL4+Y8IGxh
XXow6cQWL5e9W5cArWz9+z+EnC2iyzA8GOM64L516SMVOq/IAgKETUXvx+5+ofWfjuCrVuC2DQgH
5lS1TSixPd+WKrSaN661TDpneODAkOsOo1G2o05LCFylP/iAIH1ULvZB7k4zHieFUr0caeuO4aor
eVa+BdmrqDHZJQyMCxzZ3GC2uZOchItu6PTqFdwJp8waZNxV33Z1R/fNqIuw+8zq3yvvYoYyH1zh
N/bjQM7bOWvtL+DULs+jE9VrgS/Jg38Cl0vJBak5SdqfGBWLITeVlG6KEnoYjPkMJfb8naxDhqRb
orN/BsGNBdH2RkUSPGcFY+x3++/ZM7S8ZKKbtYE7a4Q5GPWapHJsxplXAuoNZ2TtmwHViAxLkVRL
3iYxJx5LabihSbZ6tFyoZdzOfqqJLZnxJ82mQbcyYcZvqwlIwkTjzJBnH+uvmaiKvoGst5dgsJ/K
ezMcm1J5dABZvVsvwlPvi3u9nqGng/gHprCGqg+iFnjVlnbxg3mF1+f2InAlbKVl8uaqAWL1aeAX
OLNr5c+k3n0+asWJv1tMkJEuTTF+YdKhjsMcSVgFmSN4mSU/871Jozxk32OznAWfgGlFYXL913Xo
hcBLAN95vlComoXwspP9uFWbHxsyWUai80rP8t7scCOFPnwpFOkms7W+yG3WsRbEhZ9qzVhutztE
91eaglAYpO4sAjau66yRwEo0+Hh4q0AhRAmfvlOCzAkqbv62mJ2LA8/Zlql9jzD7qt7zoxEH8pJM
694lJ5VzrWObzEDQ+LVXXcUAvNQlfq9NpSuS5qS17oaieHQZ+EsGsX5KEoxB6coVPBUd0eQ3hc5p
06seitKGm6Vy13CShpwTMkKmHzGyGpXRxFC3W7SoXBg7R46g957e1OUqR6H8bQy6IzS4x8AwRnwi
FfyZggXLmHDKiKred/KO1WNzM2CnnYvtONdAJ787zQDJA+dCg1sjfEdou3e4OyazV8/xPYSrbu1Y
YRd0jgiYdEFyPeRs/M+VGDXuBNPMV+25wTvlFp18qeN27zkMMVn/zPCuqX46ABfO7n5vBH/WGq59
5rPpqK+gKUVDlqWGdO1+qhhX/XUesF13bisHGkL/BOheClE3ax4EIDSuBFAPFcIRxBkm7jdjjRS9
1z874SMupCJ+fybgctSj4LZU+6p6PLE7uzZ+dzbePIGo+v2AUk8Efyl4XtP2VqP/OlIEl+aUijFV
xDaVoJ2+jWF8A58ivvn5+Z8xu0Ks+7M/8POF9oo1tKXAtiQaf1fPscxmR/1lc5UdqPRj66hDJ0vT
BJEq/ebK7TQxUMHeCQcu3PbH2JRsLt9pYUGw8KJmx+xsV9EFd9MY9L45ceU0JLMvBiKvVFXLYvYZ
vAfu81KzBQATN9hzbVWa2yemSFASuPUsIAtKYswNt81ye2Y/5YmUmD1c+z94K7QPK3b/hfqEU10z
q3yO3hkG4YBhznvWa9FzPNZZDui5zp9QdMNGl375B2IJSSztZPcHIiu0s80lrHWuoiObkoXGW7Ei
wO4mblhiDsinqjQQ0uqylyyGXVSVhfT7krA9g7coKu3xpt/T8A1S8rPSl2Ecu3k1bEXmPH2lC1L4
axYSrmzOLu3b9xG3WGmLLIC555Celt2+Dj67wDuKxxSl3kiH4Wxq6XWSnndmDZ7Rrr2eDv1w3T0u
BkEWTLCTFq7Bd0ImfJGVKl2qSbvVa10Ea8vxkBF/xsD4kVwoH/5HAldXrUf3E4ldg++4zn5clpCF
+NxAgNKsqCZjJrXPAgFB97oC6tNZ/qPJxxNjdAQOrPKX+AQrw08/YZ5gP6qMtkLCS9mjxfb5fs/H
mzNEuOAKSop5nBpmWa+LKrDJG4HDi21c0lnDk4Tg3U2LXZd82dSjCBI+bWzaLwYX/xU8UN5Nc8BT
YDl6w+7qQwI8rMBMNdvsLbR+5lq0wRwN4wpPNjcMw7EAR7K6+VQp5XVrfdDEAFTxVZBYXLbzv3wk
TLHCz8hwugnAi59MbD4mffyLl2tpDql6/N9bhxFUCEKogi6VKuxwrKtzlsA630pW+tXHxX2IMqD1
l3Bf2soFoygCyNYZuiOAICqACTu+JlG52A/xzMB+wXtlkEOPkSrWJP4d1sEBlYq3DZ8mtcGLPrbd
BcYXaJ41yYY+2ogbayUbGW7LHsi4tpqXoPGIhWsZoGGDHn+XhoGVk+RxReEyLKoYcEQMNfEt+ZJV
7nkbOQBbjw2ByT0UF18uFwi9R5iU4ylLXafYpBBXJnYvE6SB5QjI/oe8h5uYn7c2khXqhSWuJAUR
asgW/IqElpivjgRdvfBAy3HbjYFs5PemonuX+xNqi44abQNlQMBGxqOBkXBcg1cWkoxaSkMq84ue
IYOp6i24FEdeeU1sfzO0IeQ2wh2gwea7b4HqC6QVlDyyw+lTsxUumMPlVC9vMUmqKHt5Rw4twTpn
KO+we0G8p9EKMWdgMwptmX+E9xjAAQvMcC+J8f5QMiouU96Vbn3RDuGv6I+FSTJb+eK3JsrUBim4
RehgsvEC8VcEDuBwlV9erRGgag0Myjtp5S8RNURpYkf2OZGfvIl9lYBabDHLgqu/MXlqtH9ZahvG
a9yNO3qt449UG6L3SCc3zjTZOjXZMOw6oYtA8kY0t63mQt5fj0AnuNAwjz4UJ7jTHGZns9Xjm1vG
YOUUO6wqRtXmsIYqjp3iaBEU9HRQZ1lZGGVZ+4SaM+lWwGEvvm4LX9MGqcTAKyZu58PDl2QDE+tV
QydEVSBlV3Jf6nTifBSYE7f9hQPnZkwhIxAicSPu3ImS+iJqMcZru3ARz5007rkAEB7Ff38KVvMY
aoyrkMXhegMpR9zMxURC4vksefhLkCwoIxPbLAW/b/GqngikKTb5rDHNoT1s4xMM6YmXYxPd+C71
4+w3gIyaUGy1tLOjSzJq/F1M36jpFVSDGb0phl81dPqZtmxoSnB6rS4RNYaZPnEaqtg/SIAJdSxU
uFLypBL86H1T/chgtT8x0gglYrzPBlNPTDyBIzHWKjvW1YhOsl5YxDyPh9KlU/2N181lBPJO+FXq
FUTNy6SO/Ey8qZmi9+LhDYB6LQPO1Pv4OyA4Vj2o2BX6lW+tIOToYHHweU5oVz9mKzrixRkZ10Ag
7ROvXi5g7pmA3zNwEBXo6rNfPApa+GazsA1OFMylZqJ7QE1th6eXbaWTdskiE0y3QQTu4aWiwHB1
S89fJxpZXHYVUUlw/YOtGzm9qZ8Z360jYfNgVFSzlw7GI9umS52pVDFW2mtkOt5OsUMZr9qhUBNP
oTci2U2ID90FLUhDF2kdC9GfBSeJDp6TfSiTLodhELBBNl42eugLLtV/7P4mB7PWZG2zZgFUqSut
8X308TQUm0f/xvYJKmSQYYIiDCNofnK6vYw/oxYk+fBkYYg6wnJDo5+hAXdL9E2mTVepLcvSqgSd
TqczAs3myerP4R42NFgk67uNZiOAndaQTbPgCstPIN9ThmmQYqSNXeblmaMLFrtKHZ4ReY+EujEp
Bat4SOu8akkuafKuTrqw8EcnfXKLrjruD5VNWHG1aRnu8cOxNmV+25mbNep6/BbY06p6XGPYY99s
CzKxicoUOkHsjD113byVDmUBzsC45mbQAopM9/xEkGO3x7DNBxh33QAAK2UgVT4G4vP+JV9PSzJ2
Ygg/4hF44JHvUhJk6u+AYapkIE1OArFM2xSCUiit01Y2jv0j/z3Fe9N8mBvpTClx9YBxKp21RnAp
tzwLieM/8zfQTAgqBZox0bSXeqgJu4mnr2II1PIUaV6wb5p1kNScGKHkH+f+Hf7GW5yOB+XN6v/C
fndmje9ryPzhX/9qQL/P4HB8B7QL067/66Jy8xdXaJMAlIMX0btW8b4QnQg4W67J8owgO695Ow8b
3Lx+HjlUsg0KKH8Y/BClKbkTupWuHRT9/aoI5LjPiB5x+czG5CO+rUhruFDX6kmLnHl56FuPM/Mo
yvQ6dCkQx9Tnf3XF/h7iY0mCcCIFgBcOSMQpFRavOeskFEHZ4fYIHC3FiFN410YxkAXWUx7yx2Iq
Ckh0FusEnNYXdOzkgdPh4tlc8CDNLa11iXuhd5yFGdNct4H8odbF2kmTzlzehXubt25KKQwpldc4
B/yfEPDywET85cZxqKMAfgRjuQCUDFXw/t7WJt6v6tepOJ+pojfCeemnmQvR9eualiQWUYqoxUxC
fgzgTmNp5NIu4JUwVjcuy69/Gy0bxnIb/nGeM13q+7hnQn8F5xmC4InHKUs5EsBzM4Ca3qLztIgH
sCJYCSd/tXH4fK9sAhfz88mwVBDY6ft4tCAL6r94VuEHtHG2MIpOQpg9WKLkxjavj0sLKYeyYoya
IASAIftXKum81/eiDZQ5Gju9dsXiaKt4dhgg4m/MNTbZg3rSNIPe7VPRZ/OTNGeH+R62lc2HmFzl
shUjXdzq+a7tP73YwFSI+gYPu/s7jmC9t97mc40hkUAl8tilkXrfNPyqozwkerA6j39JnIHehHi/
2zf2wJkd98tVnlFKgimSC/22pWKJqMG0RqmkZ432qY5/ACSUfBuRVISJtRbjbAO5qZcpxgLqL2lb
4SkfTKVajOR+rKxxRvHvRj1Nm+JwI+Is4qJkNUr2INew7J4nnPf0xHltkNv4JTcUwH96hJceXTjI
URT4JU0O9AEN481lTzYAELsNVIPxFkq7+YVJiacw5qBDdIQpNGsR3trXqW/MW+jnl7WtffP7mVVS
PpLFKVssWhcVPm3jjAhF6sGoS6pDQCGek99ZG4x1pUejwybg4rei1EfawfE6JHffI4F7K7nNBTT8
s6ZwwWIGIAB7jaYYr+b8GFGofcN5zXtHdzDFNUhzkxxluMTKB7/HCkRmWTfED378J7sUJ7R7nxzF
TuYsB5aDHy2yIDqAtDcqwgIRoeD0wBr644zUFCQ1JKBNxnGS5yiGEF+4vVAFetQuSU6hMrkIGXlO
cFEn+LOV59PzoFInJXeYYh1EtbPY4lZg23BVmVq4pYKz1W9D8r/dUuBIG+SNo4mwSKLgHBZDHSlA
5leLKyq0mKvdc44ML6OwOSZcrW87Nj9muRxAZi/0XhO/jmlPSN9TDhTbFkKSj4VR3KSne2j/B7lv
VJRmVjc8aE8Dsbjg4ppYIyg4Hc7Rb4t/Obbms1way+r5lCLpJUQOZM9+xhSVpEI5L3V8VbgvCHSg
JGlfYQxeMYOHsvg8mYjiKpe9K3Y+6RHiZIMnxNM4jgb4HtIGtctcqK4M1jtxq4vsXRlqmMmldzr6
4AoZct/xpuG3rXLkslUjjBzLQ/W0HZbq/Z7bxqCpCL54Ge5JENLzxySlM1bl7eKRKR61gqI0Xwre
jw1Gf/Qa3XajXsHpWyd93asdnX8huedYIK6mOiRjP3EdFEuHcb/NS9ok1VGmJsEUYZbNP9S7Wh6J
LaDdclqHxB7c0nQKOWy5JfsMs5XMBxACyQf+WGwUIJw2+iSHRFZPfTj8m7s1q6z3IU3zjkhDxpNL
VrJudC0bdWclqbVRS7ZAFs3qunyysFCUhL5Dr2oY31g/CZtt1/TIdH8ygekha7J0yV3lkLRTyeP5
JvjUiZSbbnBbIiV8V+iMvLvYGMupF9ORAWFqu86MAS+RMY9XF6rcvK/n9BD5uUoVjzeLozcMo1ai
prfipe1pdy8WM2NeouXklSfEK5qOOGuJc1CirqwKBcI6uHDdD6Rq04FnrpanzKkSPCeMUhIINLj7
DpNjYrLdmfdTaEdpIvOjMZVwdMbeQ8KzCfkPB4ZI3m3YhXrlyzvt/25dedZbJuktzF1kaj1HGwPd
Mwwl+HXTQsxn3nr37HxMWNfqreVcnEUzo7jZlgqmUtrKxyCOZoW7RBbQ/MfE+e3Hjcm2kkpDWHvy
cA0i0fDXQb3I4CPPj8bIWHb9c8/MfxjIQENCgTp0qlVzuu3mViO0q2NPiv9jncMFtVxptNJq1/pA
qwGIFKroG4JzAJcVbBH7tuMy837VRjTvozityeOO2QhwL/kJUvB4L1bQzhhclKiXNa/0MSPz+myZ
ueddPJxXy3TX6XT3wchE/jnO71QT7OyG7OoC8tLzaIVN1PLit5QJmBrN+oaugXGhYLOepuGipRcn
puJx2qW+OYp5UN8hL/NVU/29Ow4V98+RfG2GQxJgIdxl26CbScWWgq7sH52kGWjNFq+mBLoYncqF
OW/roHsLtx3oX716rvUQirzVgvnxfId9lboOQLegLR0TKz5ZhwxxfYhYufQvf4A4BbsvjwW11riy
Id0GyuJByXNlQtpjP7ArEYh6FS79kQg96lCQJpaxYFz6ZZBRk8YDsei3Np632gT5K4auBdxnfKKe
6SCtnzK4tnDngo51PXEtOFZ//zoHToLyyW6PhIKt+Pf/mnkx4hRgkbaWZ77+6LjRFF647fb/uDmD
hmEexABNAFhcfG3/Vxvg/GCmk6v7RJj9h2tgjsWfIAL37UabUFJsBPrAf8nZ+s07ZeUmKk5wK8QH
lj9Q0I+9xPZq0WUmOg92qOtWSxszTAghJAf1Se5CuyFDGFOw/+Lu7Xk9PxhBoBEA9EkMi05l2HJh
+aw5cIexbrsDmZCBWuj7kqOVcE4QczN19k7lpmB3ZUSRVUAQPbSvVgvaV9NnnVlslXUGbuhkq3qw
qsSThAQSztw2FWCWID4Lo6JumtXPXUFdVvn+cLCmjjaDAamxshBi4C5TCbG/9/PZcrc0FkXbMC1j
puh9pgZ58ZuVyVWbTEoAO8KIB0qGKyDeIF0Sj78xyD9Nm2cmNMSxDi54wCiMKvIQO/l70I1y9D63
g9NASBVn7Y0pCI4Viqx7vm0YTHOlaQifDyMZx4kxfVS95iO/VJHs/RzhSe18jaJzmWZSFoWNOwpp
BbB6tvHKEh6N2Df4YNH6KKZ5jd/5mn8P9Yg3W6PMUtD7b7/R1nv9qDNtyIWASNSxQg9i1pIVSETZ
tt+uC0bnqD7n4Ploj26TERVpZ29Gc4a0vlpBMbhVoR+/3+Ju9+ehaIjOWgk1kben87X6G+3cjoMW
k/KST0wqhLkfnJRiM8v7WELkeUq0dip1IYz/wAn7Ui/Z46HxZbrDj9o54mRDxNy40HuQUGrYmMTw
xKS0YGLWrj+B+WcJFDhrEowLIfjqi69VGxSHmTiTWU58KLMH0EyfyfjZKJ93hElH3b9YIxd5UjJ4
yrp6jK/0qh4bLigEfcUqWN7S0js2CihKMpRjUjYTGwnf+LS2tWss6xDMkVfRanpFaVAysKi5p22k
B9LeOWHjZaIO/0MMvOulZ6ZVESl7v7LVIGKzf5iE0BQKkPZ9GmGiEAGviecflCeOzTgcsIYb9TnL
ZDFaJur1WKstK/u6ggDhMK+R2MNsdYrMvCC8l5/oMSDqVjeyQZQi4Iv/UQwDn+rqFQRC5uHb8R9N
jNY+RGCXUEmp9IisWDR5I2nZVHl+6jNGU19AzCU5MHHXKwRka6l4Ttn8v5TsnsRNe2pxCHq5DnEK
1b3VxCfPQW8qpA4zeD3cp/RoHioMzoav6Zv61r454oJzfQFCjNSEHuC82COCTqxaoSnndobJRm5Y
ipwPAiQTMuft15ShoW5Vari9YnqxWGWKI7UJXNTSTVtkQ7KarKqmTPeRX5OnOYNuqBND/ZWWh4N/
NB7I5oVTJbcfJ4lnEl6r23GWYG8PyMWv6HI22ARqN6jORcgS1vLT+m0QaTfFx2dBH7ie2UDTbZYr
mgovmCGJ5976U+QhJYiTJPwpLixPgeGpRq2TkTR3ucEF4cGB7a+q6hph9Z5YpQYtVIqcQNntUdil
bJXFuYR+jRlwenBD0o66ULra5cO7teshOrCSFetBrqUAA99m/QGtWfsxWoZytE6Ady0FV4eltbLx
JSP52QWpcjkuWdycdVmSbC2V6YNLmvPQPS7AFhLMzEuM1CGl9yuWjFZK0ITzX2iOHJF/VTrEtnvX
s0v7gLgT8nrhHodKJJwxUq0XPzrIbwUf9jkUtyckuDlCLVutgNf2hPD7W315vXQKPU9LpQyrpkpd
wxjtr+Voi+mH3joq4sQr8Uxd/l1fuCP6PdipxnS+mPFsrfsvU67S0OlDATT44KkLdDekDW07crbp
WeJvRU7bzAJcO+ThpulbqxltI8Qd4QzkeLQljrXKQM6cay3is0jNaikZOt3Of7YOtlh3Eq4J0BWr
c1lUinGazgxHpS8+CmYXJm1k86szeEQEvp042ILEAvucSbhFtj2gvtBdqdSHI3JzQg16tl5eA/Kt
ZqzUpvgVqf4WcY6RJ2Sp+sVAqsD1qy737ktLXLPKBz4bIM8AIXPf30VVQnbkNWAEclc/C2yka4Cf
n9o+qeTCXvUDwTkFBewjbvn29w2Pb4sYNpV5DI8Ku6zPyKyT96cg3fcCtgRSlZcEHg5HIWoTzweH
hRrVjlW0jcVnb8JBj14AUDPmchBtB4y8jmDvIcdyH9tz8fx1OZoIQBJ4OZa6vi7YE0IqNXOZ59ga
zoUYnoQRYMFhtDber/gjPMpba/CGkjWo/cRRzLgg6XMlVsP7K7Rzt77Gf3lxoTOPpEOzcjVfcuEA
AxHi+hankxtqxiKAkgeuOvETtIpmvLhRP4IYJx9jyDNZkVuvvgRKTNI+VA0Izn0UBo72wtTeiHlh
PSduUNZBrHLk7G0/tmPu9UjYqdQlGwe9mvBBQwfqoaanSG4E6D13Xr/5zxrHKPztQ2GwZRNHvp9Z
+uXt24LMkeCYMfKjyZilKImq4Gxu3ahCMRmljb/WuYldTnXgrhvhb13LSfa3aLDGwRdkDGh9U6Ph
ktEPj8YCGNWMm8ZHwYXxJuGm0oIPskKJNMTpTcbbVENpUrrMgn1FBA+r+yDWtA4JC7JnDcKziRl6
HrpWF4y+E7H7sZibulR7GwFTJtT/hyeHf1GBcQ4V8MgSJ3+Rjw4UJ2eCsljKOYoTp7C852hdBmY3
W0j+xAumkNEcPhV7NVhiYvP+QoZCQDWGjq/lIRdPx7YEhuBGsLlPwvyIt4jmZLcBJsgYU0oQlfvO
9p2AXcuBrJ19Bohfkd6ozqBCRVnzxcmUEr+uTQgBLlFVT/QWDTeC86ykJ2PxWlP2MbaluNTtJS0F
JAH5tnn2DYVZCPEBfaoNb5uofKmcuOJi9l+EV02iMKSLr0MVQBbVa4+0pEZ5eIXjeIIldXf3OiSd
G7F+pYqNnr6+XH0AV9P6O2sQkq05IPn6Fcl6Hh15xh2BETDHSuotdm6STtXoFWvDBnXq+pRmlBsy
lFSYtqKvEnDDEP2Nz/FBruUUILQ1yQV0WnWdS6TkvDc/VdMinliX4E/8jSglSVUvFeS0+IXh6eGr
yd/nO/OO8xnXqrZXQntmFZzWjvrq7UzF1AlW7Ura/r+SwH79DaPTqdqUiRjlgwvmzLJDWw/Aj2ea
8GM0hAL7lHHfgun1IddfuChICNZZgAGBcmF00QmOmMZO/NuOiHlOnynftW44k8Bk6H79YxEoQfEu
I9DPPxTMiojcf65IthqpMQpJzD8qRiHIxt8Zt+BVJz051mU0vdjKnYnNaXRoSbPMKYc9pWZyP4aA
RyGEppgFbbQj4V6OndkzeqZ42YBjwLG+8+8xnU2b/T1oXEW6JqWDSroi4pEwLZN1lfOezAsAuaum
lDZ4M5cgsn3YKKabfCIvFvIF6S89ST5ZrsMxnTKxxbG004AiA/jRa0zgMxR8ao2nm0sgUgqJEscc
c7hP4ZkLTroa/96tzkV2I+LUCqWQ6dK/aolmKh7cWBIGqee/u2QESB6yiIWDHyRWrfyGnEyP1Hv5
RSVTguo/IJLJjuKWLhlrUFJBu/C4Qmd5oAegIHVd/hWkVJqYaeFrytDvlRX5mOaT0+CFlScPwamX
5hN5KRvm9J28uLRXypNIZo8SlQRiXXhjMS8rEb4Z7AvNwdsW4K9QCSTW7zlgto0Kgtziw7npu5R7
Ctta1TS4nNSyMOXopV2AvgPw22g462zsL1PqwloTVOrr/VZKoXS894yRnksuBeSCrW5j+zpivnjh
1KGwexbX2AREpZYb9y47x90q+IQCBNVatG6DG6HI2QuWg76Td1GQD4EEwKgJYqMcHOA6ZYCAO7iw
GXYETifr4Ii6ITzJIJvbiXmiv7VF5o/A7emd0LbQRtoKHf3ekjW3DUuMFyhd10lrdbIBhDg/a8Co
bLOG1c5n+Lfco2GOtMeIcgthqydGbTmpEhHbMy0uFsbGR7rYeT2czzcY/LnR4bwK89yzUBHwwMc7
JWodFuJkoY0DBjCPuzuOsh1U4T18vJ24KTq8OsJiPw0IpIu7c4E6jsWIYz6n2ebkWpn9tnC+G7sH
axGxwEqaAUdu1BKSveBXxUzKvPgkUSjDER22yjKYUcWJxp+omLBNg2hVpkRUBfiZT3A/pNuwtGvE
7SzGoKczlwK1X134LeeCuC0M2fJV3sKxAzrozQktCg95YF3iNwP2hVcgLna8s4PdNQFKM8g+QADJ
1RN4VQ1T9JLCRJqX3/G9DoIwy3RYX7sHHv1AwE5xRPvqh7JYrpOUKhaOuBX5zx3LfYGrBhnDobXA
f6Uqcvys0Bpyhif+5LBfYHRrK3jahBZyIH8+x8X0Th/M/3GdLSfoqHeRVCsU7arV/6TQTN4EOj+c
qYKOvNuh2RP30LZ4TmoNF6G0mwwZa69XVLGXbWyRrccg1wq5ui/vZsNYTXyO+Nx8B8P4O37jVXFA
Gy595zRRO+cK7rgFjb2vMIA0M7qunzFd2vX3jiKec5Stlu5QySKeL/rbIZYr6ywftWynJBufLaBW
0JYe/lejNmUUWdWfhqv+tEo8Sl/lfnMEr1I1GIKUoqhJEnBA9WU/PJB/8fmgqjEP3MzQctGl6yeL
u1/1ByTbV2726ZP5d9ybIwKH2zus0ZPXMClgJXWiXBe670grxz8D66rXwVPcD71pIZ3qlTxQFtlw
fX2WsCLCvgtxzr7SeJssWW1wXw3v3Z6h/vb0hyeh2hQKDGWvrrCGPHZkA6lFDdUS/KrCxYoJXyF+
4c7xfit3pa3yDYuqy4pInBMOuCl3L8Hwe0pdAX8P+Y1aa/0zcS8qIP7BYiXakb57h4wHtd9eyFx8
Q/XtYNSDvubyErT2txi+SfgL9wiDDtabgkT9inoS4RILnFhm14QFjbmDMdbWkNN4Ytpk09hgN0T9
+OcdtuFsqr8NXU2ovC8yRO3OF780wgJuYxxSwJpkmiEaSMD1j2k4e7sEnIEIZmowvFdOhl8cZ/QD
ZSf5s2/hIzc1nPDBKWAqlyUFx5mfKQT+4V5sGOFo0hX43JH7Z5ySIS1CG7m/CNSYS2wbYKFE8EzS
z9WZ6I1MOgXDBBmg4vxShxc3A7NwkARgvoCHmsBdwpr+5b9rvoSOylCMTpWMiv7ssD7ghlpWlIHz
NTQ6BPRoa4GIarFW/PKYLBJlKMQsS7L67HrFYnidpEvtFt2uMakexrgIsshEPQCSwpeniIV0MtYQ
VQ843PXiXbFyC1vxUN81LI/Sd6JhxP3gWWO5DeuQ/s2hPUet1EdT+/BqoZk1NzDx0+89sUYMBin3
OTaexWAVUVeDnlZNaep6+iiU2buG1p+1i72kkKTuztKRFC5fcQglPxeJo8HP8C/UMa/1BOuB3Zyp
qvForMtZQ2U+pz3l7XnrgZNp5L4Z4LlPbKv3NMwm4tiSrvR5SMwM4Lv+xtnp9mj1YimaT1+TNYSB
4iQWcfage8Aj1yOMJAZA6PBaQf9A5maci/vo/VbHqEDH7z9fk106SZkj4e5Zl8/9+3P4vccmdLus
bWFoomk8YYG8IlirZBCAxmsFL13mpg1A2ZSQi0LFHZTrqOVRoTEmtWlrMa+h3qS83WNkmK5C0W2M
pfAzHr8qZmGFbf/NhtiL8KMeRY/fZbTg7liRgRRI3TGUK3I+8/Et0aIbwwfjqLy6TG1Flkq8TCfC
1NQAFwiga7b0ygm/e2qnmUYcz0k9cWio9/g/2M445zO0sO8BHVj+x8ZE57xUf3OP6NQEExg/RWEg
rNXuX5sALgNfq26O1CnKYaj4LlOr5MYUdYMM5Oe1G1N0eQhwCAmmEcs1SifeU+Rap6WzICZzmhKz
1f8dSOY3aibOUSS5sp/O9qzMfd+DJ7KR70WInxUA2wsMZh74+fvpPnOT+mBhpShrLhbxMPTrDyds
3ko5aLZig1kykSQXg36+byL2x69vixuPy4GzkQibBDuADDFejPmMDRNO4bZzeSKwFDn36SWCnNRN
FuS0HAH0e48307XKy94mQBaTt0suM0XuVvodu7Ez/JZcu3VY8+rNLSyy1H69zXS7vuefwERPhTQl
CE9EdYhZI5yYPHAYCm1alHN1iGGO6tCp6MLda4EumFQwrCWcAEXx9HEATZSQ9otF2N90TMKxNjaR
L0TYxlMG7Au6SfYYUWwUK3Gj7M8CzqKE7ARRry95iCe0XrNhYXLSXT+wie8jxuHRg2gKsX7KFiUv
IYVX98ZveBseizG6M8V48fo8Xzz8+dmmWm/KqnmcqEssVR0S63n8RWJyvsP71GJG0K2m2LUHy9LI
JSUaZzvJmr68O4ohfH15ufq5NFRMHVeoOn+4XIsfRUmUcwJYcE2X3hZM/kUoS1c/0PM2R8GNYkqH
bByJGfw2zqaPxwdPsjaaoepjWJPduYr0bHNHt4TDxC4y2PduHceMRNI8zocLi/4/DGvHue0C7sbS
nzXstdV1utfpzo1cYaN84dLMIFPgNF9yqN0Y89Xl6YHbkQzbs7x6HpXEr+tycSD2Ek3yOpnGmMmH
LQX4X4TZS4ZRaOEW2bq2JIDJQycJaQaHPzvVKvGjdl69sku7XMArAmS5goYI8PiskNLvFWdotVqu
UbzK3Jq3NDUId8XWPZj4uMPbhkvuOpXdk0m3Ikw5Y/+PJ9tsVQpzz8U0GPDcC5ChhLvIcPDPlP4q
RSZi8Pvs+SW6FkaX1mVbAZXYYUnh95Tsk8oRezBMozRmO0aCfrbQ8qqnEo8vGgvgHoMJO62I3/Pz
gwNoXykh6heMWuL1AgWYsrPldwda+CGwlc0Sj1R1Thk6ObRt4vON1cOVZQIsaN+66rHOI5oxEx2I
mqjdVVpT2yPsWzopNdRr+mPXO0qYT03YjJTm/Sg/gxGNVlW4nXAZAUTpZsdU2pge4dXfWwo4P29a
qUJEl/lfxUrw25srKBTUmjjfQhVot1uWB8S9Ov0zSsSY/no4wVoyvdex43kj8hLBSOIQF6dJCaA8
ha/0hT1zSBrrKoSs7KYjP2pjZs/h2NTf8g0vLn/mI+CcwFe0YbL/1diGb2kdYTIxb9twEDzSuQn2
O5ft87ViOt6pDDSedA2FQ0YlbW73Ai2T6ml50DeuK2+ujY8lzkToEjQxWtSi6UtWdmCVVZjRbIXz
gTUkoP0oIM2HGFeccMTrrvauTp4RUWwL8RBxSANFtalo2OyjmjuDuWH3idPC8rAgQay0UMeGh8fp
xSBvt82dp/dbOsdGDtS0/h5+R01y4bMN+VGXGbHo0zpz3tnPE8/o15o5a2uhoHLByy0wM7w+JquF
G90LlOS8QXEUYBcIyHoFZq08v2vC3InWJnNS2XcKw1hjytMA3Pvs7HWIAWGsDTWlhL2wB1NrbHq4
XUneZzgGr0e/DHKMKYNu/VdrMpq/54TFCUWF/if9a8tASoDwhh6cdBXLzXTts/wFNBsrwGtML0F1
d6xEb5YY+rXvzGgf5caspSvUWz5O9vTSW/+VGVAviR7o5y7gzSMSyFUpUmnE7zkwxVkX+qkM+DC+
gDRzyVbxUVU4gUzQu2+r25xoVaA3QET+ffO12MdoUfPw0IuqkHcZ8fCZeY22Kp7l1Q+nQ7PWE/uF
66BwiG1h5xbLA5Jrw6jN3/rgRawCa9W/q/XOs+zoWmWv0GH7DcnM4v0vbNR5OW4e/yAaH+fDLdoe
Yj+F3J1nWbXGk8ksDpf77ry4Zyk8yO8T71WtmaV+f2H61m77WkGWj+5Jb7DjtygO0ykaH39ia80g
aSmwoczeISYM6zNg5SZNT4E8NrNmiulCwJYLU/JIkBnFDBSYCk1pmUPwjqmphQG2U/SL36PrqGRd
wlp80AnKj90RMv9Vqnt17hge+5o0/ZfzmzYnDX8gtU9abrm3g2aqOJDvpHkvr6b+c5TRbc2xGxTt
F1VG845YS+WwyCCzoM0lOv7TLyLBuZTFNmuQTnKBH/RxCCl1w+hodIBvYgq1G8m1o0qRSg5hrBXj
HlYL0fQ/ga7I8iixFucv1nJyx4RhFa+yBZU7hnffSmbikGZBYSTw6twVf7Q27YoDhVEQQKzVgOUb
4Bdja3xJjk7AV7mvI/mLlR1srMEySHAt3ss9cNYd5BL0PZU+2qIYJKkPpgqJIVci1Dy6Diad5cUU
m0Wn7WVERiGRnteTAiKFeRckfPsPSe+V56lwZk+S3UeZDm1WfiPkbJOZeU4nI72MpDugsRlFfbOM
Pn2w8ZdHff11eYHl4NJLWBod7tVhXaV1ekjyTM9dhCEvuverGqJJC9Oz0QArwcrXYdSv8ucb5+S2
gzX8XtShJxzd2deROZPfv55oam5Csyo3cHWHMkhxoH9bQuiUeTgjfqWhta86LicasZHQCJ56Ip/b
KeBRpWLdU43J5LUjmImNt4JWD1doRJUb+oV1ibPxGpjlkLAUirsMjBnn4Ec/95I5W0UoXECtj/vG
GYvAbTjmKbrXFoLxwrL5sQNb4174ptpbJaewEq6EUg8f2nzl04izffLdGM9lxGLJcG89mms2Gr4d
GxDoh6+cyRKa3sgj7eQ1UDDfR28CwKLcm591pSEPb7Zt7V8ZGSDDWlWGeEIngFrYi6JJJzgIfJvE
fVv7fATUtm7YkwcSrrl3VW2PDgQlkQf8tn3YhgddJ8mupdX8jO1LCzqRuI8hEYQXSJHjTMKltcMx
Gk2oqW6aIK0FExEfz/6uFj3qdNyojjHHwK2Gs0c3F0zFvKEmcq6i1xzR2S63FwRb+J5jXNUSUxWa
N/Fdl0tzxx1ODQj8CR7EghhOWN0/u0uiXcbr7yvPNCJoR9gkVLUjVoUjN7bUSlYEbU+JI+UlfPVY
iTAyr3Ac9LyJv2YwB+zwo1YJdjiRsBCFcztgnj54Uvs1H3mf+pew2/EW1TMmVDcLfpTdUWF4fljV
0xM0fMwRUzz1cAWe/VOdsDa7iU/t8fSApa13Ohcs3sH0mi19Ttm2m5b+A6qlg+UQURRwLJJrL2+J
OJi+KIyE0Jf6MEmns5SXvU0jOhMelkRn2zMnKbP+Fy/woSVFLYQe9/lmGvZFcuNmgHVNeTM4/4Ra
HAiK6C8S2FBmg4sWo9LmNwxgKJ2q9A2opG2UBlZdY4LKy8yV15j9IstmJ4QQ/7owGTbC6JL0WSvM
TcX7XrE1pb5I6b4rSgVQiv3T21XnQs5g0AxKYVtDiEOnkAn9UT9oW1eVuaLA2MTeeeb4QsAIuGVD
gzc51SzLJtmVco10l5hsVPlX6ejCMe/V1aycZ8TDbJfsNzn09EDoXjWgz83rT9nGpHJIXDqatL2D
zhnYEMTVABjA7pTlDjdCrCQxSKwOmjatASoqgiI6YfE/Qw4/SHX/Z2dR/9aQECu3Y/NKvU1cDQ8E
IdFMeOwIGkrIeOisc/QXDgejVpEFlHUftW9R9k3CZK8q47hDKYLudaZ39AOhONDlV75gXglCpy1J
DkniyqSnD+cGvYxokA4x7OPDOsc1xe1H6rp/kESibTUeE3l7y8eSBYztXShHiSc0zvZP3+TVkEWP
+nzFz6jhiTGaCUodT5du+Fk+l5tfkTzzFErkyjqId90Hi0M5w+54yYUam6RmO+x8EBlzXZJfq/wH
SimZ8+AHOQ8+27R77CpCSf+C5T7iIgyPzsIA1SnBA7V79hYDqw4NCitKsFVYnCEYj46Sl98GR7EU
khpT1p5+smnZM9BI/4m1CmLF+e8CiqE5cQw6qGytwJqJ2njaG0jnRCMkGcqCppRFKnPNqmlqbMcA
RhLVr3321++tUe6bfY0wpoYKnX+7fRsBIVDAl2jSmTiMGdhf5NZr4T/EON2c1axn9dASKjXVGiG8
k8knHH5171yiD10HxdyxlUYgxzdnejuAY9x1mbi4nslwqVOM+Ji6aMkxrqranyv/61tC+5HllRsb
uUvypy/cEfuVXNWYrHaQl7wVCpN+seT6ZgC+ir5DK+BZregDNztEW8PLyskuy5R3zAEo9TN166b4
qulpg91415YtD5/qJCGO616vEv0lrOgwuKdn3KQrHr3mB0kjf457xGzJ06g1Cil+FWtRm6TZM6n7
ZC2iTtESFlaYb2uzizQ8yaEMUPEWJEJo2TPp0kcn3GTiAK0azPAyZCw5uE+VJeEGWr3z3BdS9G9s
IdbyaqxWjJST3LNqW0INJS6JplobSpQmJr41ctVz28G9vOae5IWouGFCkAHGb8g2t11/OI8+RUfU
7AKZxbjE8xqfsUsJs5lr2UHPiGxwSpx0fHQe1VE1fgwSsBMdNNcXx+VT35qTnMbne8O2OcEhWtUM
bBGVYJjygkTedqWRkdW5wYHh84gV9W6bLHrbwpV6auKijGIiY4uLkMtZUl4k3nDHbNoS8RT9oaaA
khI8IYJtrT5oTJoBl0cwgeRNePInM1t5cWgHlF2jGVumBU6G/68GXZwIWM+c2i9tfpajgOMiYusr
+V/gOZvsYdToYJIaFWCHIxH8HLOuZMFIkjPghWgTFgjpOLP3lHnERNwLP2zrjGO8iljTdDza6AA0
bRLVInYc9beAU+2+NTP1BZsYN70wDuOQzqvH47YL9wXRX0Uz7xA1o8oMP+Xc31mnnasw9hXSKl9j
qqN3VSIGViEQ17cJttHMCuduA81d06Cu1N8Ho0pXpEt2Df9u/8xw3UTlo2oZlto9/wHCat5HrrU1
3Gdz4sm+FyrLwVjX4shdIQLqxzzP+h9aM0Dw/WXzwiYo2Cl5hUs8mQ5gg7appPbqBZheUMJXT5G8
RWs5bg9BHbU1HLI+tmXIfKWzIGLfZX/EPgn4Vi77j3H1BZhZIc1B7I+STbv5J04wxAsBLHCSwKXf
CQY+MABNbPmOTZ8MDrROPc/5eO1u38Vk6tsCSKgshQc68Tj3cHVNyEnOGuVJ6rHHd+XcnTYj5sBH
m59FdSaJElqHsDe+T9iGmNzDRMXxlyYR5zOQKcr4cx3BrGgUONX78RwqueJ4A28oM7iMlDJa4ydD
Ya2osiC70tD+YmK0XIVla9OOzKMllp5m/UCbTKFTTDyOI2aM6u75Fxs2Wl35su7dzoUSYHPputpX
TbW33nnyR/rIjJ0Xuvliv3/hlSFZIt4KPJN6ROabzFDbCxzHSO5k5c/mFSYWbYHuUD41/5EIrlvn
N6bwiZQZiVT/CfGgCSYQH9Ae2H2+UftgCmVwFci8V5HFWlM/8Ja61Oic9NmPixI8HrfmA+r5R/MV
NqEHrEihO+9iKqEIBb1PlOen2Ck4I08GJfESlB5bz3M8nXX53PIt6QYB6Lzgj+uUPlD+ve7RwGl9
Kt9uI2WFaoX0TByFoLzfjpl685lugAt44EPO7FXS/BIpQSQAbZhe1iDB51d2wrIB4Ddvo+jS0w+5
d1t2E3B21vhK4pQnZN1tqAFIjm6pKIWs4Jhb4QtRngXWEPBrXfNxmTWCD/ZJKrDoADWLQpUn5aqs
je+o/oc+l7IKQqdy8kLR6Mwha+SMG0N0uNGwwJA4UACBBNiL18U/wrudw0uk8Kh16l2czDTj7zsX
sK6xSn2264CTH1EyPEFYpf5BTNZa9IC7cQ5Z29VaRwwfeGVb9AlpEJKH/11Dxk6/WatjBn5h2t5Q
Z2LAMFlkEBfoYwfkftM6xdKALCWEadBNC/mFH7XwszluetVHo1lq+jTRtbpYmLT8mK97moNFoJCV
Am1fSfPz0Jam+GBZcjG7Ais7Im4bF/H8SBFUkqTOP9O3HgcEBm3sg140HqUGEZ8jSnLDi8R7rndt
3ReystxSSEq/OIyLqYYWZCmS5Jc+A2F9swJfgWDZt+x/rKMiAHYsdHr/CgW05Rl/Scdl7hlFDQ8a
5W4EyWX9Sf/gsdUZoVMEUh+oVvqdbc1nFbp4ptB+j+y+eqXe1UbbNed3lrLqiSmeFzQ06vh9+jCN
BMId3E6xioNlTkPy1Iu/VkLQ4hjgV48LCAbUFazL5GW90bcAxc+WTwLjleI+oRpJYnExLLo6+lOV
xi27TGNYQFunfQ9Vrak114SSErd9ssLOJ6BzIVMTi2Z6aAvuWamrSvZJpNqSkazHpZZZq60Iyx6o
eCYPVx5sKqPXcUgPD30060Uc2kuB6NATq6FBCYEukO1LNr8XpXpVtpqrm/TgCnSIBuryzpNA0FRv
SCl9tEDE9uY+BryoohVGs+aiUekKOa7MW6PKN26Usb9XQ34/7YrDE8SA5aTlpi2IrIpSzpNoNAZV
uQFBzhM0HaHB3kiE6jc/xLeIPDlKgdKUXS1Lz9alZikL54U75lVASMTFHTytHnNB+YXyWNs3o+E5
6wMYC1ji4a6elHr/V7hKW+bnIi4BoyUx6LaTDtqmbqo6qPmoZNMaKQpFLu8NeqE6nuJH8yCybzc0
kY9TlmxyjmjCBvaijELLQkshDupPjgWfy8DcmSLIbS76i3j4EQYo6WOotZNuYILBsEGkReT6tS4m
1PSN0dI4Kf9s/zIeSbDL6ZMzTu/gwI5RkF/CWPT2xTVH/b3cbB/uV5e5WCBMFrIHnCXlgSo5mhEB
+KirZfYgxeqpUK/bnVdMRRMU2YvHsw5z94ka5HTpku0pwIKPuBlFrOJM9W30daaO7k4zE/amI77e
2oRs5q+vNATJ8FMtasDhV1oTLknRoY4lXINQLtJXcipRfZZDmSLgrUq97raDw4gkOqLGlkmq++Oh
UePH8uj8c6RMSqtp4lVngMWYvDSOP75HycKQCHhUco8EN494U8rRjvfOrSr6/ITmkov9eNtLJjyv
TL+UIyGAPFKz4oC4HNAW7+1TBlS1tZADIFDS33lUCR4hsnPYv/X2BZjnbHFGmLIVR3D9pmkoSwO4
LIEnF6me7+Wi5pDcJ6HyefKzbqqpUVcy74a2QaNjLUgeCf/2CQ3CL7MWI+vu80b7V6VApHBtSX+Y
ABBCgibs2+XzNdUHQDPM4p3gkIJKtxpidl/5AEJ5WCRXIgQjnJ/iFJ9h6qA+XO5yN8JNI+VHsGDb
XDyLK4o4KKS0PO1f2HH2YEUp6yZ9keybB5nSfJ7AL+edF8VhslU2SnVrYBMGdw5HDkJeBgVukZSc
GJvpiiwllsFU/ofCRa15Y4VDo0XNCDXlJV5uKq31heLNsx3Tssed8ICoQwumXBRQR61/rRc4yUhq
q97qcGnmGaB2gHU3jhkeUTpLfjChaGMI9ejs2kcW6Ksdx2NxC9f2Os9J/PZjabdJnM5RD70QyfEx
nMJeEPaGnu9FHNqTeAgTFRN03bAVllUIPr++2EtZ48Rfx2bIw8c2LJ87vXJXrqINclFfIRlA4LDE
5+i1znyaEozzTk7DvwbmQJe8BMgP/gfY3Do3cL6KWvJzayCTfYOHlQKoR8uAvYQvItonrViFgkzr
U54iQsQrBdNjbnSUiD66xim6N2tEWvHuwkyt2bchBXgrmDH8DFUIJ1lwpEgv0t1dlPFOklBIWW7F
01hVFMmrbZDsSmcFey8kKyKocH5nqDYGy7EmDlWAivtViwxRZq9Rx7n6NFPXfY0vKDrYgoj/P+oV
OXEa0j5hIZKuk1iCZzh8zWDHx34+/oGUCfEZUteQR43i8xn5OygFJBBCPz43ylfRetN1e+diTFns
gIxl14Y0T/Yk009Qtpe+IP7asI7F69OU98RD0Ky/Goi/CO6y7xcjc5Gpr84M1teDKsR9hI/4nn9p
vM/7ZvswEGEhuVM3F31LLQJByL5wbgW5WULZ+mekLZxrnYB/4zuCQ9yZh+ChBdu0sqJcZT7O80cn
ULHgcHgeI7DalHNg23pF+qqjc9qj5g1rdRFKfdoktzTvtbd94vggFDfWqKMo2l3/TuBTED0MC4pc
t2T2pC5+Mwg/IcIXScpO/zoMq9U5gZUsb8SyatKX5scnu7NG55M/1DpcT5fTjnvD18Sa75nJGKJ9
+3k+JvXOcyuPAlD0mHh6UWwvUJebgEE6M0OKKT1qw6xe0fitTU/GLvp0jF1wbmDPlGf2TxWiCRAX
9fqif9xXHOqVsJAy2DI0XDGAotY+k8S4mCwXwm1SPUyTVTCNCS6fikdQmG5mVQ70nPftvnujra9R
z9Dcg0RqonNTjQpGSBBXs8seILUtXHVETK1xhumnHOKQSNOIA0CXSA1dVmPg9gu8Qm7ggocFKYRz
qyy9mzhOBEYo9l3xinNREU8aAKcgX2kaYq2LDjuJSNMH4IoJ4+Sn00KJin+swh0/7t1ZuHLo33Ik
3AZDuCrzVd2vXw+J/syHnLdH8diozex8oRYGK3nrthcavmTnygVNJVt4VlnbscC2rWUpBo2IqZ+2
2t2Cxq86EDPBBNRv1Gy30uWOTfE0SOWi1fbaEzgEtHao9PzlSAn02vZYAE4K+MJabz93IPhkCH8e
DdV/ZtVMfQbyABgOk884uKzeQhaNAWf+BmIIfrNJFJu8ys91li5l5WmCseydUv31wk7sZbwpaWBu
arhKmmCqy55w2YyxPG3K2IVXPssSgA6RvAM21ertCYVOASymyGZUrIuhrEt6+l8lvVOy9nlZSwpG
xDq0sMahzJZdwaEabK2zO9Ty+7bnDMHHVHBCR5Xd+S8o37hqOMJ5Prsz1JBXn/8c1VK80qDApRBN
6/52NNoL/HsRaJVxahGb9cULZon0d+xhdE+rYyg9PRgm5+d2HRCX8xY+VCV94DZN2l/flHpa8qtt
nIjjp/ozoxP+m7cVC+IwkWmS3xhcz81PSNsh30gujUrjOco/eqtxB26fgQHqcKL16fuzCCqyAzS4
kD5hC7Lv7Lfbg0BxcR+Ni6go92LpxaAcGkRVaBD46zILgY6CMdPTQnSgiIFnpjTARk7sa2yoPsZy
lXWEjkNMzSB0Dj9yFCb9BVoY1tUGOX13VWrJv/0/Gg/8tiU+RQUoL3oWZ+/II0RPCmRG4sdlYJIB
Jb49eYuXl/IRPiXTAyC4AJ93BUtWc3r2qjqC0R52M0xvxyuRB0B8QpyvL+FPwT850O5W+Q3jQ10m
VX713X+PjtZrHhG56xyFxazr7eCPdVhTN27esmngc86L5FkBe4cC37PX6gbloPA2DgvlY+JjKlDX
uh/1OQEvSuPiR52TMlzgELxABMQFmeeju3v0Wr2Z7NX7WhjUig+zmbT3oN4RE2eZroa4XKQfZDAc
jXCU6IdeeN9FoLRxSd1dp1vREi/MrEIZKKvk4/KtTT1aR5HyuRdqufK96WYC9TCoTDo4NY8lnOTW
8uJSkYkRdgHVwIzG7Pdoim2iVmTo4GvEtzRwpw/Yb35stVgFmvERCY6cikFN6Evb0GRla8yWo5LY
vYgFl3Ub2CqbS6xdXoFSwfj5HL4Nv2IUtw98dgzg+07sdfxKSNkcmQHEcQKMWtpXXBBJwlpSDRIQ
56KRali4U6HenH3c73+wRVZYpi8mUMaB7iKpwAGQAjR7cDursyOOwGpHHkhWk1G5f8VojPn2p2cl
wV//jqvry4dKcu4XcklKdXhIM5erPv2JGJ4HCdPTk3yvDvZizyloK0fOGd2UxbmPTJfAdtLPbvx3
n1iNiFLeyunMgIxtnfS/oHqX6AuAJthSfBF1XSgtN3gNL0SqHODugzOxfWu5FLujN1YoVxVIplId
gtsmqaxama0M7iT7YQuS7xOAd0OKR6B71TWQhp87BJG/Zj8/bEICxPu0UYaghkudOkPFSf1sk/F9
kkv5WGWuy0GXCe893ECsn5bQcvIZYiCXOBwZJYlgcdj3BW3Rb5WPGaQXFJh9JcfpBeaE27NqMSxI
pDVClU69kRVp7EnS5XROw4lml8FG8C/GJ+2Mqq+e12qB0tOPDfU/ksF82VXdz/uC7VbeK8CkQKJZ
d8RD4Ach5yxc8SyTtj6r6RQZkOkm2VA0wY39AynyV7psfQLXu1Esqsl6cbVKaRvIg1XB5u4/uf0w
6baQtYsn4zOI/ecBbNg32eX1FWojvSZ5PCmFt3r8cc8GyylBq/Noe8bfDGva8y3Rkb8DiPHoR4q9
OVJocCaJsyMbsWmQI18Qd0DiE1XNMAhJRmyDW1+jTmLl2Kk5YmPv7mbJ5qQhCBlH8pALEcuveW8n
Uvv4hAPJJ5+sOTqCUbsx6aIci4fos6DzHYV8pO5+GdKWbuD3/Etf0LohJUBUk1Hd/hqFGYYIeU0G
D36eWVpVA710AGqHZ7+Z8mVWuSjEiaVvhy701lWuEl6gbJMMs3CUVTCPUydgfIIBtkpisqVuQWRS
beIy5V2vxtEi+IeyrQq+xNHTfaQHK712ZAUQOMwrdtMVEWgaY3fj3WOmfNOui7U2jEoL7Hh45YC+
+TqfPhLZ5kfBXyozfQmh7WG2Pf6wLTmJPaRpSOqEabXfoeibFw9huaRKhQbgWN9DxnDoo5Xnzwui
Nckwxkx8ymysFULhdQ8BHWNhZMigWxei6C9mdA9TdSFstBMlJq2MzVdCooTItM3CTXwAzcnMzQZ0
cN2gYFslC3YQsG6C5GzrykZKUoLWgnv9HU67tUfzOsG8zvVobgG3f4t9BITB971MaOJO6j4EWZpO
Azuz5QrFNK4XjqQIgyQr7a1q6I1MUuI/harwpuWiGn0D1leT0Mn+6VqdNveX4aQG+i/me7bhbYE+
kIjKfcqOQxmL94ezuSlBfvm+YdMguuf5oaAeRNBwUJi4AI1dysS9iVqrljwyrcpSg4iLV46nMOnE
wy/7pWz4hzDdtuRaun1uMk1iMNvUd7r4402NG8O0Zcbt7SJ7JKE13JDdIDqeh9gxybSPMT8ySPGm
FZkAKPk2mZK0ivdicYBtG59opkp6xfxv7iASkV+3cQT9HoNpTIDYjnejrrdxLzL46OYCHggoA9cO
cNI2jCWwg1FCiL4EMM3ckgKpOyr4IrwMU2C01ygxr5fdk98nPBlIpn0Aw1FLOUtMnKsR76EcJP57
DUAmqUKHcBvTORUQAqxvM4uK6UldZVon5blEyz4EB5mH46p6pERO5I2E8spQx5leKJJAHeCJJm5v
unbTuknWM+yz8jFjcniIFNgvxvu0qIzioZYBDpbr6Nf+Q89cYEIrRZhkFq7b2ZNPfsvx+pZIHrqC
G82nIqn5KydGFOisi0SEPrp0wNd/VBJVJjZSKKINj9XHdKTbO2YDNP1svLHaDfnplhhPPX+okA7b
CXRza4EWYN0B58GgiHjGur6TVRFAgDVG5pPb7N5qUqAqVQpEpFR992YXqjH5yyIQ9s38wNe4AbKZ
2EEPTM18imVI4KT2kuPmUbotjVhXBdiD3DabcNcXnq8l9bLaaHyLturnOBp1+gYlgL90MHY1rH5r
16TPCMosvxEO4HuhgYVUa2OlQBSNFXo0E0XdtluRGdAkQY0AZco0pctc3yOvwyUC9cVXBmgniBLQ
kARCWpgD0k1EZzeXw1WsBjKPK2NnN7y8ioAWSniRN15r5qDnuvtC2DjH1b2heC9JG03InYNmHkpq
0REgc7SC0PZA8HMb9uwUVbpAGkC+BrnMCUJEXyipoM9ibZzi61h+j0jSo43hRwlDgXtNAU8mvOZa
KntjM3D+gyNdD+G0yS+92zRj/UPecCWXofUY1mF0Cyqh+t4ElKTVyEnnymbt14/+JX6a1nDDB4YK
fciyaP9im1JnCyB+Czr8z516eBG3q2wyVE5FUQnj0fzwWiSZ4zMvOWorv1nnsp2D9AtpyTqFUHIg
+9xkXrbVpYTvT6csI+Rf1QXneXDJQI5oo5g62j2vh5QnlvF440l9tEoTUebnh5nSSjdX3QfyOz5d
yX+viKxDHe4ZKGLQ9UldyBaY8I0zB8BAhj6JLcx2fCfoBRaNbA2Itt3eiId3fXYC1LeoI0oLnuA7
y3+0AdHf4nsX5e9QlgX9M1Wf+vwKj7M2TquzmHptBVTf2KOq0tD81B2IaGGcKaARxxuICOKeVngJ
SaOBuNOviXdwlXtK/YTDX3d1Mc3/Any+mXZVgUq6a3HUlS97Fl45X8aHvvZ88O8GkQyR6VL68grl
16V/wT0wevF57FZ9rDWtoxCYtxKFYXWUEI49ZAgqCberdlo55Tjqnw86WU6hoqdTSG0p9+xqRQLz
KrDPCItlK+5f/8fZDpjU8Voyn4evE29aNj/tnJ4pN0EbMBOA1U750+Mo26JrST0mivFFhJ6x2NY1
zQNcHFXKutRAk5Rpt7KEj2r/tYbbJaswUGxE5np5+kb3vYEEfdJZ5eh+5rvExNEJKb8Mu4J/aCmm
kcNEMhwsECL7WlUHP+AnZK5lL1k1a09UrojhNQ2QVbvd4zRSBFb7vKTTYpMSJsv4xtZsWAnbdtsh
niNVK5AQtDiyH3b5J0EwU77wW/Qv1b8E8w7BS+VXB6RJJZW3Tem/ObHB6OjKapTN8MaBjik34hk+
gQWs/eyZ7j/3avEt8sFV20Swx2zDhSgu487IHyBaZx+Gz0xm/i7sMIqye0xHuRx5k7fJQ+QWRBNx
GZ6N8CUxgA5yOGbHJTcnDJ84ONZxQboWfdHlYYhypGp/PfPRFOnvPAFMB3vax4dQmEo5nr3iMU6A
NmrjSjtSg9qc1+015DYkJoIWQ7OAmwbGg5wg+pjer+Wv6fCkagOyvJqkJgdwyeOVEd9tWniI9RVs
JiUJ6+J5DjhODEZDJh1mLsC9J4DwboxCiOLKZLNymtmfz8pJeIHhKDAMnSgrP547aw34QbKXtRnq
hPY8NHafdbQ8y5JoqQkQjhjDURO7qW0N+0fvaA/lVYZRPgJsPlAuLs9cjlJCufuHBwacjFzHzARS
N0buoE8BKuLd6Qn6HUZfOBnmjJRLouYbm8FStUPCfc3TAYyQhGGv1xkphnLt6Vz3/zKpupdkUGbe
wbWiuMdx4LyyolQoyy8KDz+7Wixuh51TizCF8y53ST7DraahNipbYUSvssmJeuPrtbuKdz0NpwhM
B5SJRbFOHggj/6je2VMaDdK+l1gCJRzjyqLr8p1h8TX2KM2ILdMZ40vtynQUsDtxXioUwdDZ6dc3
XVWwTRMgMxJNOZ6LijHTt5DSD3XeznW6Fxu4uVKRYAs78mWU3ZrXFiiqBb66kMdAgxfuIortHb/t
a+HMqt8iuNoVtns41SPLxXgwDD8m+BsUOMOByazwH6uJZD1KlEspxc9AwsksowEzk9wkNcj2+frO
BC7+I3A5mwyQzqRIGUfznYgFbuBQjb/QvsRAWBP3lyzt2srM0wb8ctc7Sugj+R/EhYMyaY5weaRt
3/5jV51V4Ks2vo80DngaxBQLF4CbJS2Yz+cQqRdiYAt+Ybiu7KIVHuH79+qRpQcQAFuvJZ2t5VJL
BaIL3XFZ+WkcJmk25uAZrgsk7+LTpINhN2/dJoF54a0mVlxpDyrMPbTkAHZgARc40MZmOgLsTrDB
bXp8karLUy/wr6MmhvANnGBXtGE4apkLzGlUj8XLfOJJzOt6OBC8P4fU94gcFX8HUIZLr8OKvSQ2
5gi/52/DOOOsDmQgpJKQyruDu73wiDxXc6vO/0DKukO0jeEyLAVaxIgdeNtQdomKz3izXJ59jPrJ
AC2SEKKbJPj5xlBCy4LMBfljJGW8j2rwa8+cMGKOHkKltB3OdCN1vU/uMbfv+napdu+oKdPYSFuf
JL7jjyLi3pDa8YHiBLZuwOTjHGg6b1qadHVHBaH0govfclj+Xqy7uqHVGnhePI9fI44f/wBP/kVm
4mRYxjBFXPk3pWB2017zTCG8XEKWXNiGt/pI7ozJ8Lb5ANQDapUrIWaPt5SJ8F/K7yt7cYOTURWW
Rij6cTBlHsr5ZyWshnpzO6fWaQ2jqae1VRj2tvW/SvGAm0VuQ/HGmQvb/CeyUSceLLJKA5g10r3w
MQaScz+IgRo4G6b65px2wWBoKC71faUimTyLlVbWm/xnmrOH0erEDkW2qdAIFabpgWRzF5DsXxUd
ALdBxvZZwZlrkOqMD8HCUdwDEb/nYTsKm8RM952557lfG/fvtb/VkfAlm9H8W2T4A/KcC9BEjA6p
UqpvGw3MZSUEHdiyUrthbk4n95adb84uUGtA8SQu2Luw9M8iLP+1wKxazZDu2wjuXZms2nc8x7PY
v4/ozElye9aMnQa8L9ctojYaWKaIDGWWZSDVe+Uka9YfPQuPZsqCpIEFZEUDttKp/989uSZ2gJew
Nam++qQvuqFHh1y3Ht6YpWuZh6Df6pgUiBqUMpmu3xBK4K+gemNNs3pit1PaXq7DPnx+EeYxVA0e
+06LoQhDJr+MvmJL5B//6qIiHnC4k5oP1KZ4X6h5gnCgZA29wKF2TfgKveStkM3cxT7lLGbR9gfZ
0dYakcVSgxyfsHapB2KyqjGtFLVXCuPjAWHy/xFDYL3gThi5x69Mbydx4FyPAd4hgMlAb4fSEAxT
BN7GORtYXtYfrnDCaNrvakA9ayziAZGo851K3Yif6QJt5VPyzlVXxTFWjOqGy6ZSbcfROxhf6ZET
i2PClzrt7AaicjICRNVVcDgKchSC0NJx+lg2ByGParPCh9dtN25TWBnqEXNGpuaTzfEAXlitkW19
kdWqT3gG8XZJxup3oGD+HMHOIp+X4jYfVUGSok0hfUEdWWzvq0NZN4mL+RLfwSBzGbV+kWUPADUL
YNIxjPtWyOd+8717mrdLzpoAcMdSbkqCsDPL6h5dBstKagdGSCRNzPee//XW5QHJMgmXyNopVAcc
gLPxx5vYyxQw7fjFEBT3wP0qNf01LMxuuYeB/Ga0iOeDaq0Jm8SnweQKJ4mGEQVlFKAiWN0xnaHK
/UTbOwTd9RKzEvHOIlvv54MTql36GvdIyqD80ItqBsX5D90L8TPfVFS9103NmD6ibHQJAuqBFGZe
iROYsWB2nWZ4IzrV8rheL+MRDu0Ozl32kuPpslSRDQwAZCTZpNaaH35DyI4zYRG7d+zsoReNcZ1v
md3kijD+eiRaBgT0UsmAJdhhu9msc/WNYYGc647N9KGMcFxSiHlP8bYRKnbg9lsS0O3njIjtSUT0
eJbuDo1UmEOmJYaAreF0FjH7RCNJ0Nh/wMzve84064SvUaP+lBwJso8bs2m+fy1Q3hplD+TwkLFT
Wpx+lmzEEUAcYp6BdhbgT+oBy3hbhs8v4oyUpe27ntYQNcV/i/WhSND663XZwUVKrnjSBr1GAcWO
MQ/vIVqPHDJLRMoRbUz+uvxUeUe+Fv4pOVvGBzvd7OlfRfyGV6X2hbeuBRlDmeMLZnICblXisP3+
XJqxEH5t8v+uT8m1lbksWOLm0/giwE9Mv7mcsIN4s583Mw1HwhU388s54JqkMT2KxKbo/DHGFMRx
h9M9PL8FUy5vNDYaMIsa+Cnt6C7kuzrY4r9hX9MgVpDn8mRqB0GC9T/1UrO+bTzN1pAsb4N9SQsB
4h2pabsSufYUBM7zSBR+qA+Jh0Wbb2l59Bs5vDD0+f9Bpczfu/HS4vzNKfu8bl8VnbRMzX4KwWh4
VBlfsqb0J1rEZBFfCaLpOOYD0jQv7TVpOopEqm1mnHlGnRtKCc+C9V12m2wdd0+X+mmiPmX9vjbU
gLa+3OQpFOFDrX7W3W5op/7NDQJLhmGlqg5janSznsACcD15k1ric2a1Vlxo0MzOfgwrdDZhpa5c
tMxDjLp4FgUx2vLvfqmZtwdBWoKZbYaKb3xLLLhsJhNTltD0/mBTNbUD2PKVkUfcgUJxJooBmMzx
CEGxGHf4SGND49AOKd5bFxgwzRHrpobn0nWJKANuE7KNZdpGNJwuwt2qygkw51hW16DRE8i0z93o
/Ay9L7r84fuuP1Qon0JSULKOGja73VixdkMyC7aPTafhsBFJ+VLWCnZ+5iph8w7KKUK8Ia9IEuTS
VY8ktLuYQ1ccdfB9k5pjtarV9uS+kav61X1651ZO4Uvlk3f6DcMkNvsL5VUmMK9MMMOWmPa/Mxr7
wGTBJpDmX6QWwz805X1ZYTtJAhuSM0jnUOoRPYYI7jVhAiH1nzEmGtgwUDnDYTzmyQpim0TrFtf1
GiL/GAZIieS3KhK74lxsCMAvDdwRIwTZMyM8jgwmSBA58OF0a3ER8xwaWhwfmnXkhzdoDPJNTexC
yEMWIRlpD/YpgAqBD/Ypdp7XhBof/FnJoy+kOseuJKqRjF1rosI7Sq3uWWZD3JVL3gJ5wA4SKeBV
3T10aePF37DvwIsFpM4I7WLs6HBUOeb8jICy5A46U2K3feL76LEvv5d079SLy2EuxBzSruTUazGM
wOb8PLeZIhKtPopO9Vg0C++Ep4GWuojneXJamSHzuWcxuG7dpizi0zVFR0YUdVeaGo646RiQD/Fm
B9AmQA6LUuB7x+PsGhrTLNhn+bfVPeFQgUbFD4NnSroD2fzOYU/L19CUFVXjVS8vonRLdg77eciO
+hc8VjoLzDglD4YZocNxvlunDHUPggERamsyRfvWJjCIftdofxZmRWUE5AvuI+Jr+/9uIwnHyKjk
x5fn7jWk08FtgMglOWlxO0X3hFr2u0ezaBFF2KGBhK6Cyvm22XvgQ97qxZUiOIbtBsNrHRQ+BY7z
WKYUF4APpwcIzriuPhzc/YvSIUnwmOkxKJY7p/YmU4e6HwnWfmzAAgwUf9ZBRkash86Kz0sPk18U
NlDbDpuB/M9Ep2rXsj5KB5GMeLPuuWXtsLwwBqmKiyct83l20tpx+tPA1b18iBwbgggjrfXxz+ft
LnuwAIBiIHCkpBT28yHByRSmPY3qpew+1uMlA3ApYjBe2pcvt+GizloxJzLWsH+n3KSnQ0Q4FzOk
dwwNV6+fdfq/dDCwPLPAQ++Dv+iQcMOVJse9YVVcaSOiDgwFMhuixvjqT0oKtxBe9oFRZZbq0xdj
6npz281zoQwaTjPf0jrwW8yzanA3Y81XLBQjwwCTNKyCxH/7FendpX9IbyyF6St/Bjcd3AUXwI7J
trAFqAqF9BAlFcZYL/zjnaxk6Bl62vy/bYlIfPXv86RV9vVCNDg0v7EtiHyQAiBBTtwpeJkCvVB4
vj5AiM7h2DzGlVDIRNhBVv7KKJRZ9m8H2FG2Oo4JaapPeYWOGGgbrbP+f4NYYk3gAwIKwIlFeAzB
B2f+PP2oOCIu7Uaadw45zEgFcwAuDvyj9a06SFrhnUAWo9fgcvu1mN7ANrBKnQx56J8VyX5QROwQ
P2JT1orn9mzPWVKbboBhDs7w+A5Pg9znfyG9xLqjcxhrieEJoxjjEefrn5JQqBygMprMAR8Vym92
IxnXDJTGYepehx+r3PX7708iSzPBDNzshLHiYQ8BY1PHM2fqyHwArUDwBIz7+1y5seBLdiHFmaI2
94EkeiE61I/8Yuzei6ucecHqT6GAajvYLc2v695x77T/MnvREWl48Yj3PSNhppjU9qYkoc9cIccA
3nvkmdacspQ+p84E7E8V3zZxh1ROheNCIoVIHOGm5PtiIZ0nopGrpdBx4GTK9wZbLnFuDjaLXL3u
gLbdcrdTRgoMMj7XIpuzJoK9CPD9Kt2rwV5O1CJGRvgWggChFpJS6Z/Bhy2VgSQp1q3Nbp5OuQIs
TCwBSpBKkWXel6k7eMBDaLSITY0zURpJV/cNwadEJMS6IJPsOfu3hrGoggBu6LOCwiEvw7xy0wWk
AqH2Exa99jP3GAZ607fGIxELJNQ2tXVjNkoODcAr4wl3qabv8i3f6vJJHXctDGB49wl/DtJE9/r3
h8s61FJpcROuY6WbdTHouCl2myjVWMYnrJW8TEhzU8QZ+ZDaNSw8tEJdrN9xWsJEX1dz8Qs9T82z
ICHJARD19afxEqcZCcJ9UavQL2OHgCQRufJPSU+/d3G66YQ7Ep5zgWeLGOcxHp3ILDJVtShW0vGV
b9O/WGyIjussgqAm7EvCh+4E5Cnwmkln7TfoTTVjv1hFCSoRoD+Jxr6tZS5sFrMgLz2fddWGU4qj
3vu9Ci8/DMb2lP9OIravzVNMV7rcYP0Y8/Dyg1zF+bIr8Ki10gG1oaXhUrelJhvjMsc1IOBrQGiT
g7mmGS8FHNMlqQS10cKmbhhhJnOqcPRBTuPJkb7IhuoRzehAwu86MkBaXesbaNd2bnVBCKW3Ztt9
X7H0vkkrM1Gi5atwufOry6/h4G6FgCXPHXqUzne1Y03NHaQypBbFS04GSDIQ92pGE8AJw9SV15et
7b3/7WiKFtcVNB+RVHFOWppg7XSqij15cRpbOIiQXyUwiW0ztmtx0KgScxVlweQllb7XdXqhYdzt
KCspIJMvl+9Sb8WlcoN9p1yKfp43WyvHWWgvKLOvMm5D72A6nBj+6KG4sIByNQKOUCzjXD6KHP30
zS8RJbIkXNxceaLTdRFa5fpoKLBVK3126L8BrLjz0nLrLWXUOtr3L6cNn4bRqizmotfYTfQ6t2Yl
enFMEMCyvqAo3rBTRLyQR1KkDfEoYNdYQaRDqzQ4bJw47I3okImEZNYKL/iJi5jg0I0mFj+8H62b
jVu5xS8ylmevWrw2f0yg1Zhj5Eq8w0Cq51ZhoUeLUX6Z940Tn8I2TgPgBEE5BT91CVt6CjXClg8G
p+yvVQUnTgFaYFpts3vZOQa8uAXfQs3PGOcYkbC4LtANrhqRtpbXog3b+l/R9deuTtPXkmBnX1Sr
QgH1adVzHASIMYHPy/QPkxStwVI3qZqdaU4JatpN+jN8zrPwHOOinPjCrLDWgjwQuE5i9Y7M6FwK
SFQOZGngA1KdTqQ0ZgdvzEyYA9lWHz4cvoUR7Dz7hJ+JIfSmah0JC3Eetdcz9L3IL8lxSLi/uj+2
QP7TrsHSHjBdJeCV8vrHJ8DtBBLjJVpgnn5SiMHf9ozrQbYA36uy88JeKRs4vbAwybcWHMj3IjGs
UQekLcwjqovuKwphkGdIehE4BMa/j96WygHacVCVk2HX253UoX6F/WBN7SYlpi2LtbmgBZqbBq8g
fEs33j8rgZNRB0YFBYbQYgQV5y+3OyfyIdUXTZGs6IijwaWTQRpchJ9GjnWkj/Ctub3aoJd6Ng92
ksOc7GIRrmA3iXLE/wYUKiz9mtvIXQJQXz50/es32io3u9zWkezSGfdGbau6PC41npjfUE3aCGpe
e/YXS5KXexf5Zz9cB2YUxDW0uy2kIf7CoSFjodYL7/4AbyRCoA8OXnTFaBQfcIMENvFKynrI1gRS
cVyM9xNRLT4hW9Zr/bN32rIbQrHQA537aZ8Xkw6giG8givhDy0FN1LSrUVZNunGNHBCe7ro45iwx
anQlLRHRhAHe8NQhlBc06zMRRo1xwOD+gEAenikoH+++wO+eoKYqfack7UcZHk4yHwAaAWULJ9xp
Om8hFme42fZs86XiNVcV3l51F+k7eqYu300m0zJwKOCQsfB2oxKT/7XqTAjGPJalZ4d2RKGaREdm
d5m2pI37u+iHE8l75RNpgKUSlW+vg1OYouqTqfQW1iLhSzej8oxw/pond1tMSW+FSreSzkaQ+cnZ
fWxMY8tB/t1oVhtOXepHXUTV9sLaJv2xo7dcIRWa842oPkbN3v79ZvlgEZc21S8kyS74qc1sZ1K6
nM/WCHk8Y7P20gR3evYDRvYAlOjIkbY4iuIUGtnpq2t9Bn0GQnGxfkbkVQkEg1Sr+Dr0bx4swrRp
yXRtSwXPItJXbcVJ+LQijVztK7Yee8U/9eNs5dxRoACTHYORRJNyYMGdRr0iOlu8kH4+o8iXlbfu
WVCxZeXUyJR0fJ5j2wOeen9O88W4ZHM4bbRLtts/D0G59vnU7uJhtb/aOQyRpAtRqGNsfUhmqiUR
CEh0fWgFLLXvI1jr3BmStfT4wm5OPQpqpZKGqFT8tIw3G9+vDqSJL8y2PDD2kjL34cCakwQOCbsS
qDB+t3QcFQ87usiLGYXoXJtnXGv4HzDI4+mwP4tpYOhr3cEsnRFMC4Yh1ZVq/PDuMNLIVSI8trWE
GZAjwyAn6buzN0/tzwMhiwmk9J3WzGDrFosWY/3JbUtk4ksZ4+hL91jqTXLMTpq756U9HUj6GRnz
Jz4Gr00BuOU0gxFi6t5LtS9bDt4Eque/YgKxfbOvMHxaE5xAt1O+pTWSRYPbaJkG4UFKJEG+FbJ+
BalCmWnv4TT9WWh8PVFBRzNeDEBAFXllQ+qhNDHycQcMK1yz1h4M25qPM/BZnV/ZJXwj5tLOKfoG
Bco9WldLf6GNe3Yi8zCY8bCdRsK8Yjg1A7ATsFdWA6rqClYKOMSWKIEd24WGToeuld6TDgZGdZfq
5EJFEsWPvP2LT+vmM5IzSzLA6spbZVjBmgkpDx7w+jt4eCTNXZoh+Zj5RJ2GBT0G8j1UMN4+Tx+o
lEjgy4jlUh8S7vNP0sCIm27e/JlcJzQjTiwz8y5r87LLhPjdda7J2EH8zoeL5A8xMZZb++Vd078F
e3QWrvOekUgN2qXwmy8vkEcuCcIvWOEnHiRqmE72tlFpkC6zpS3BIBJuS1chrkgSSDXYHan65acT
9b8D7XmyDjpHhRuOq/gzSoYXZDlMe0xwbrADVLzUVW6NqB43FX5poLWMeBKQK9MdFHlI0op8TNiq
FIgor2HACYmJQPpQJjDFv/iTasbUIKBEbPqrAUaap6J2Y6V58YkCj7dIpuicT7xA9kG9uCIazxIz
66gO+wOAcpSwF77Qe3F4rXU7EwOaCy0qTeIxCHuV+cedSqwMEK8uk6EvdKKaux769BUCAaoc94JU
5UJM7Wx1Yy6cjeyryOGybgurKJLqr0HmzrSU7mb9uroWR3UX6GPhyFX1Jrb6C9Sba3/6OymxVnSd
lOMdhENBc6ddUD9VtUPJPZxiMWNQbHkg1/QOFPwEwekcp8YJ7tM2B5Rqez7LrbKBRlexZnncdrCq
jaaQKIqT2Z/u7D7biveGWKLoZfzXgMs+TK4mPcl6RM9aUGJOxI12iU/7Uu4Wt/rAUN8DZiHTVzML
ff5g8gfiYEA5KfPPBUVNqF2AzXlP8DFT4Xn2c7L+i9w0hNr4yVcdc19nHmDKZ+lew9aqXoI+na9t
qQF1xY0bRNah6YvNGBj+gdEieoRCs5Y7xWprwIr257s+OtDG06tkmr8BrXe9Ka2B9OAdyQisL4SN
8DuLZYwVR/OAhQ9pV2dLsgB/Jv7ZIzIjz3cwhLBTUI9igIJDKS7uxtTG7tPBwoDYJU1Z6Xv8Fbtg
t4FBnY4S98FaQgOm3qyrdE8RHRT30XwKcNv1tIIqiA6fh8n9Als1/IqLmN1rRqk4QyciJmLsufSF
elHZzXc545N95vmdDBEoaZvfUZ3hi2oMtOxVS6vse7u8UW7aKwfKgTpQH+kAmDqA4U8nPHPIsEWC
PyaedXbPPWby4OAaKmOHIFz2lgx0wwTIcNhJn/rO8jslZ7IR8REk8X4VC8EDZmr3o5bZJH/XDYVY
XozKWVSVub82Z/wdua8DJwPssLCb5M3wF8BEAptAT84OeG3C6wKn7nO2cuxcl65kBRrN9P+q+LPj
M7DekZc3zJ2Gn6Bz9RunedYIz7R3h7SxVH0v+zhK9Myn1/vbIO/93mmiE1EONkMep0/ViLMoaBQc
1kvG/BeGL4pPFVmI6gINldoszf+mZz3pMLfrSbmJdTN0kldVI4vOyFJvTREnVD1w0Z1WHg+bnAQN
QwMlA9gZkfyA3enJwjF96hcyuWCRaYUU4OKORPtbX3va96+QDkLZPtFbfX7Z7wXyYmT9qU9Pvomq
HoX4p7h8BQEo8qkccFGGpMHDwLV0qrmhs5xSVWPadwRXZ6xNN7Vq03vT9j8pm2a/sznRB/3XqrHV
ScfNRa/xkw4mDFPGbp63lZ5WLcP981tWIAsdDNR1B/6pOQeSzzy+yaT9STMVHuqaQgiwQ7F1E6rx
sI5yxS3iC2/dPLaSFJdlbb6kgeD82E4T4B9B+DKy58v8Z/R6QBUJbOXg53oFHLdopUjyHEKEUCe9
K7sSXdYH5L4c4vYjS6MFVvfqsYBC6DMIhhr4yL54jVpwhsG/SSHoLs/RvUx0YCtT70w9LPjwJolg
8MF1UikcEOUpNKWgZaJQDDMwO4aYrK0Kg5gY7bQVjPrcHuQzzIX7ou0Z5rr3TmfHFcBl/a7KL6Tm
9EVCss+ogQ5rRW2iL385RDhbZ1eBpwBhq2yUMVR4Id+rkYMuZNoP+SZ/iaQFOay8j6NtSTlOmbsL
tUKzKVlaqYHk4CHa92fd9jKoAz04cJeaZVgro6aWB0U/QOisYmImWpPCUUBCGFGhYGlEtT/lr5Tt
Iz5KlVxOpCuWX0LLOkjmneoEjfO0rjpK1+fJ/dWDhHtCzCti09Brnw+x+I57yToSvGoaHB/pETLK
9TwIGOEosUXn3BpuaBalFHZmjhp/0+FosL6b6IJM41TJznFOV3k5harDy/A8A8220uTR7pB1YhDO
U/1leJ6NpAx2M2L7lG+qxAeQr/pbFAe3Ef03eL8dLrCZ0asXYIsrtuZP1zjs0HTv0pdJm1XTrV7D
SkDoZDkDychfsfsyDviLMustAu9TcdtdOype959nq3JRfprjmJlRYwlRwjLdttBq5/cjEWW1IO27
jAwrLah5xtghO1BGwaPPlAcYD9ZCwZdJYtkIxZhgCFlGtHbkMew/eLhFw5VgAPxaLHkWUYLQvKlx
BiuAdWcK3E5feWoqXLHLwzAb0wuB3k8vBcAH8jDxfd+AF+3mb3oxVdOjsMgOp49wfgV42DEFKvhr
wnbQBr8i+WcZepurMj4+uQr1P0oowuP0Fvld4evlyAp+ljKM/89B4dG/A3pH29Rpg1Vp+huca9Xz
01/ZdU2iokRLO7dQW76RKn7JbZumfrxMYsEu/qpRjcP5BUXwi8ndguI3q3UknivlhZTjtxE/8Nbs
A3KR2rDF7rdwYGslZjH676ZgqmDFU+Kb6yS4RWpnW+HSy+NC6XN239H2J7BT/V1Z7ddgqkaVZEzv
KOJ3yGjxo3XQMsTps7BkbjjyC7nQfa4PvpZyQObJ8+38OyCJeCa9y4Hg8OmbMuU5K0VXe+UXSTdY
J5pEWe3YshgZc9tdgMmp9vOOlo/g9daArgJEzkO3s5/gLgyBjCSS/JeRmIvL6dV2237KCdMZEtEP
LoRGPsCYdA9iB6N0xROE01NaY0NVvLZj/SZXCh9gpTqLeZ1v/D4lJvSVq7Em28RoiVp7cUA/BtRG
mxNRwMV4NOfA3rbsiZy6Z+1XRarJNlhg79B8pPEOwsl5sw3TCqKiMXbjeTyU3DNyYHWjVHPG3wXw
7x5mxClZA9FJyPjlCvzBKIBFQF1UvZIA7pQzzi8irjgCkepmJ9BofaFjqbJxlYvwKmP1eWsNSHCV
B3A09grb9pIH2ycYeBKnKT29wrIa5yrk2lDrK1iPVHLXPWg+YOeunSqGaWMuNV50MNDRTEXzvyRe
a2UXkn8LB/TfXFrcA2sQQbQ9beeBEBR8ygA3r6t6B85JuNSw+kZ13jPcouxhqx7t08xmtr2ye9py
XGlfBE52lAqyHDH+mY2qizrV8Qh0zQq72EBeE2mXKTON+1oimtzMNGwB31COBjoL2j3U4xBiZhzi
bnn5HAlGgQYfGy/f4RZpQB5tjVb2saPMj3CEJKPWTOq9QIBtmFQCdpj11+Lgai6BPjQtpMlnhu/r
stFFrOb4LK3KlBI5NOrP3F1DRyM3L5o/Jmp7hxcjrPGGgvV+cSHV9hLUlJ65j0XHLs5IQ4CwK4O/
brn+Pm8Hc9ZZZFYdgBM4MBOSpvVKa/9ZIl3Zpfm77SbJalNTAKsYTHCkbnyYBWsPeS6oIJ2wILOs
uHoslrbG6pxTqZIIwtfd0YH5wM2DpVNRFTztRvVv5ZkqTAS8aDNfDxyn8k9hyMxTzeA3AMepRTsg
qUqAuK+raH5q99B7vYWcB7R6TGpXSscW8LTK2xSSZ7TE2f8PFMxOqRwJsS4mMMx31imuCrsx76MR
XIl1dQ3H2T2izO9ZmNniyxHYWf4pKYvGzbViZLAuH94gQMYKTZMp4Vd43oBb+i6LeyuuY/s/5J91
Pueka6OSOb84hcPCE30V2Bfrp1k+Dx85NZCJYcTn63XtevwlTJ736qDwobiZv/KSM4OhK+RNzE4e
9McOaQ1taw1kupO6Sx+mQZmxVM9PlKJfcSJ3PLs8u1KfXpELgz7mV4+Boo1i/gO/kAI8FuXm7Xbu
wQMT4HE4mpghguI0szmpElRH0XZxNImsa1lkOveIrvA05Ys+t+ENLMpmophCXr6WCokrxw8GwUQV
DxDumU9Xt23nhkLpFEZheeVAp40Z9V7e+1i+rGZe4P2X6s5c+isHoLNIHjwLb4r/XSWHqefb/Q4K
h5FT6hzI27EQUogJ3EW1Vz9DivwH1AZKxl9pF8vSrvXqHl+3pi6jOKM8D0DLvruyI8XhQDp9G+N9
0bATJ67KpySOfvGf/FWASGytm9NzY8+30ak03YlSuFPmPynq/2I0EWB2Rvr0N3AMEcVVPXsz9TuQ
ZGjmI7mXxBh1IP1FZNXEkwpyrWes/Y7fHPbtby7ZMZAXsubKDZGK4sWvjdg8uq5pLuJyXIL66YPD
BfA1apJp8UyoY4pJQO8eWSVikYM8PqJrO+A6MUqptq+L3IBKD/Ko+8GkaLGy5d7NEyAZyr8/y6ks
yqnSzJa5JgAdmTSmERdm+B2MnkjDgXnVGqvg8HEeuWSVuPqx0/K/AZ3LevsOTkoMxOp0Hz066xzm
D8u1i0Ys534omTvYqZP8r+D7G1jGCPYXvH6PABf7EYvs4+89vTM/8oPc2+5mYqcqvvxnbGxYieOp
xcssNnY1flTKY2AvUFUGF+8fXsTooFWVpqZndQXGUqUZYIZa8ka2M7npu2+EJB1y5oYx6EwP8o3z
KBrLj+Pzv4D9TFOLad9Ajy3HKp5QbKt4WhYUHuDxcQPt2q5qcYNZ/uhbYDFjryL/VyklBYRJkETL
9WyFfWUFzLgUIopZaYGXxg8DD/xr7+5uuur15N7qR/BrfikI6EbiJeybewMssp+DcAj1ZMLCYCMX
VClbM/tPPe8P2l35MIFwyBHRsWRJPZds9IX8ZiJMbR9KWKyxVXiCCtLRRroet7IkxkztgP1dYRti
yHNEQ15ebfguyJaW6AIpl/XU28PGs4sP6FT14h0zzgpS2vc5ufIBInpKTm36vhfsuXtRY9RpyPZZ
ceIsIdAlt1+jTqrcAqycwwoAQygS8KyHXxumtWIMTkoPHgJj+iBtkTAJyJi9ZwsYvllhZPxtTDeJ
2nJH0V2stFufzhqTmRn0qW2nKp5gBU2tfcDfPLFIPkuzBaOHgVHHZn7MU91cHx6V0wmB/SdNbdhP
v4SlSGu7j+lKETzINHHdT3sV+zkwcZPBK5M8Qf/KN8l/lhdOkL8Zz0rT89CwWjUTkcDFqEQWpFv/
vE5HpTaIIHgiMAWIm5ThO1ox+tJPfgkhFvKTWnQjEDJt8jgFKrcGttC5Q1KpN4VaTaX1LU8lxaav
1OTcWNftejqD2YHyg6GcXM8uNmA8U+fLBN9J4Q/IUN131g4uxGgPGUcIZe8O6G8FkHycgkbZa2A9
Np/tW45cd3Nmb0yKqocHEI0BQOqGY/D5oZsItCTBW7+QUVoTfQWwexLGnLfH8OM6+hX0eMiJHs2Y
lnXm+bLjKM6rx4qv3AEgxh/by7kVYXC/fi496PS0FOKpBr+pHT/Vndhw7sUwN0arAJIsCZ5VO8ZA
XoIEfAFcQKuf9ImmBANqWGb5LMnMST0/pG5d71kL5ndv2QoN6rS1DDA+NLXtwPzEs05hOrM2W4Sq
9+iYDM7eSTjQ/Wr9iBsFSTcI4xC0JonAw6TXwObjp9Q/RGV7D/JjtFw1fuz1MLpZu0n1Zb7uxGBk
TymCYpLwcGHmS0woA/lqxrBK3v0J5hTablZ1VuM6fl+jtPA4NMLMw9QfF1rmqd08Jf9vr34EXPVU
pBVu//J1/xV2E2kHZfZEXYrQ2Quo5PdI1V0VEfQ+oas8gp+Lmc/xutZWuLEb/S8vedvySmXaZ5FR
nvBRxLb8YPN6p6kGFqkob7xppyI04sY8Q/uAI4oIaC6tKEoZJAPMhVXECaZ+ekgnGCOtq1gyeMdt
noKrBA5MXtZfCLSN0/aZJdXA/PE8GVtYxGWGEYQ69ALImIulUjWoejQERnyp4+TUPMnYPatfpFUY
BUrzdKDy1j7JaIJIBTdTMVvb8wPvCaV22rdKC99q2bOjZnedoRqqa+bXsUIU17KISZI7O6RR3akS
EWauIKAom84ffWOxt6b+5xPR+ejCUDmonFouc1OH65EHMX61OGj2GTwvSLT3Lw2w+JVf0IEyPhnR
PK7Zy3j4ac+AA/RoqNgxi7+jrZ2gH+80gEkAf4kTZyMYvL1ouS66fiBi8SnUn9V3zzRciWecaVuO
X8b19jM2rUlS8hlA5xLS7vOk5WGIcUBtdgIoPI+/koIrvgpkEU9fLXPmshNZbztmQbAS9L8h4kgK
1UWJuQrjSfldo4bNkeGiyr893nn87CErBWfcyKvsU/A/47c8S2Nw0LT2ikNqbOShCDMUKnFRqeP6
WUzsyMIPsqGICsV7vZE9rokwf4Af7k0i9B/rSOXKEcnaUE+1q5HfKgYQp4KGwd943yhJ9ogtA9aK
UHvqzL4TbfGsqEZGzZHAD+Bc4x0RjEkZ3zVU+0PnnrG7/0AtlmuJ27DtahCsqzZj6LdrUlMo8YDy
u8dI14vxoxMYeAhOep3NyuGBCjpBIlNKMiNGDZm8W2HKv3747VF22ImSmgq7pvioCXFhxY7vPzIJ
tJM/bpqYQJZqM/6YBOizsh3SUqF3q0XU70eqKLl6WtmZyMVSzATeE/le63I8tc1j1b+TZX+noQb4
zZTxK72kKL7oDjcMRdcZjcd4FJhn2utjRsBGm7rlfZAzxxVYasT3zUr3UTfcVYMpcCwHBD9SNzD6
N8W79thCZiEP7dhNRNAjjdggkjx9PAaOgkCP5KxP2Yj5mjesaWEvklwFX7E3puz15yUJrNdLVVdZ
iM5iVyL8zG8rrVNNhu1BHUgum0PyL8OS1FgWTy6woUu6AvgIRVQ50s6ubvfzq374FSaEb+LozOaL
z/amGuBH9iKf5laJ/NGsxWHnS3dRPEn1wnkbUjiqkOWBVF23NFnF7iOa2eMrG6hYNa7KgJ7RPYPa
V4ZF0ZyVz5O4uVtCoolV3K5XO6RNI2ARLLTS6qguvmFi2/A3uvzFCHUqWNALKUf0cz6QFLy1jH5o
h6iHTdzQ2ZtX0iLgNm0aboP4vWqMGiZoGda02w1dvUL/wG2X3QY9wUoUZyWDSZNj5W2s2E4tbWRU
xS7bvEnxuUc4Ll4NnaLbKC/yXrlFkTtWVHOu3rj2S06vnYznZNY1FL8XkuzEy2/lAXgCfCXRQaBL
gCCdMnsFaBriRi6TrxJL2o5ugefV7itGVIPc36HwXEQzLGFGWzrp5oC0roYY72xpTuOu6RWhIKDJ
dFvl6jUNUy//fNqYmRX7jOdP2wEop6GMCZBK/IUEF3UdyGg9bIWW8OO+ZVZ+7Z0kNpmTSJXdyn+q
sAf97BOfga9I84so93Jj/gBBQXCFvUwlY7kZ4J69KDNEdakJUa93okKsXgqAepyqnUxhdPxtKW1u
EQzf9a5JiMTtL8dGzey9wt+8nEZ0haI3Tn4GQw8tJycEfa7ir1PFsAnkev48/zYS7EMTWtYyuL/a
lZBXkZLv4mz2611EqRxvtJdEqBd2uKdNh2hWrcM62Ltr1mp5gYYtGFqLIc8iKcm3Y2RJxqEp4rv/
42KTdMiQxKlV2X6vwODpQspRoNdSBwD7gLmqn9ebuTQrEpUyWOnZGlJ/sn9DgRUFTjP3vlrIQI/y
s17zbCGBPmOnWL4E8G0HuUamErgX3bTqs8T+xzgmiLFf81gCKo8aQUxSJYoJoHLSPt9TDxku+O3o
SlP6rCu3q1fQTJm+avD8mNgpQ57ZlGOlSMrKLajMXAbt4u3YpAaJw4UK2PT76Pd/h44Mc5E4LO2m
1chL+kZNYjEIkhC7wXGar636uNzhkiOfu2WL3tVzS8u0ITkEt6eVffyfmVzjXHxo7wQsMolFYTw7
B8I7RGgo2cvShrqXr7c/yjxsugCF8yw94i3d7AEOZt30LhRBp4BhcJ8lwbSPgQNHtsKDd5y1Xp73
yl1BLIgNkmzwZwaDofapdMstkj8IHW1Tk+yARuevULDN2qUyg0FjZP2pikGLszSVjA0gm2qmO6Ns
GQZ4kGdksOmRnf9/yOMVp/tkzvGt9wumbJnbIg50RyfPKqH3sy7I1h1BVJtlRPawnGuXlSUVGX3K
41Niytk0v+lvZzgB+xBuvpFjOOvUMTdM7JclNAkrEBZ/s73s6fUbaMDy7auLJWbxp3z/vlXe2Lta
YEHuISs/mplK4yeGcz9botajEOCyd5e7cxOpwB3nBEPglj8SsbeAiG0DQM3KjMLogKoYn6hFckHY
mnW+kCww4y1qTHAnL2qxYGWkuTk3Obne9n/p34WMUvVd+Rrf6DZbD5AClDxUz/n4TWuNK+KOZ15q
HcgXpT43caP+Q7wkdjEVdT8eEKogqt2LpOuFY6oCTareavgzIU5hrDhGelKOBl1N4krWYzMM3+Sv
dX7WRPR5fcKurjJD2ZCMtlDDepci+CND8GoXYWJCROYs+WCnhk1WVUOUS1Ro52CKVMEsyW7jR5yZ
T5BlCh4COqxqSMbVkuuazAqkTZR3jzI+EWGJY+tvCnkrkqq6o5hJ8ShedLBl95ASOZU9rrALTEGF
aJKAF52AUyW+qpRwctMU5XPXJS7uiB5O5jPWeJhfbz9Z2+5zHpoPrtGYwo5dc+hLaZ4SvqKGNHmB
5j2zqNBjOlvTpql5Sl0BmuNl7wyJxlXGvlAVf3AxOKt+L2ZsKSIBPWWs+8u8rXLhK8KnblGdC7ua
Ej6p3AOYkdbmH5ez/IiM/8YyCBBO1dN74pkabxtVqAL9f+BmpR24ApltA8YWY/d4rPYkWP0/iVYz
kFDm+GDCXkVOArdj7NrK1haZtDxwMTVmEV+x5bNcpfVAzEVe3hQF4YlEAJJew0NZvJNDEM2K40Ig
61pmNRr+BKIu2vApTx51KRAeSaCqadlamaSJnz5PSjjLKvErEekKPOaMj7lA5muD6hlxxHWu64qz
B01aaDad42iNBM95Ad1wJBdmYyVV+e/6l5k0yIyFohj05iQTV6pJMU+wLR9YOYRF1vgzlNpSp8Xy
SG6u1U9p7/cpofz9+EYDpW1Ayjy5rm4tXdoWY2FsoD4h8TJBDJ57PwRZIGXdpb/QLK8qxaY9SNfa
W7Vx4S6FjnwYINbdy8b5OKOBLEq3XZcGZ0rLBj+n0ZVHROnDcEOqQH+OPig01j0cR1pnMniI6uFE
devCJIIv7KzM7t+dSsKNO7I1/NPb/6ffuBITga6VDNMsU8LAsW8idW1Jz2ZH/TiXn42zZg1LL+NI
ZPDxJIJpnhHl2I+h99diqf6lisehB5WAv65dWlfH9F3Z+ZZEpaNTh2vGb5U9rE34gdcyV6xmT8lX
hYNHwdsH1rEy6ZJv92FwlMKsl/oYsetOCUx2MM88JWBFFHwTBZhNkNd7VwUOtUlfVwwtCLNz6JRa
2nWAOUE28lU5Pj82YMK3qTnjZ5XYE8bm/vsOFkEFV0IKLK+fyd67O3W3K3REEiG3qYtuByqy6uZ/
j8jljqvvWox1x6GYa2soxeMUS8DFj9A5ySMQ5RCJ0Rs9xnIgmBRgTeSN5a3VZ/rps0Jmrw6xPYvy
l1QcEMy9dAADR8DlJJkSNvi6EqmMcbFKyIXQ3o1UFERGZJS+PtocuUwFVIEJ3Yp9wx3Fs6Yw0jah
cknZrMO9mF+fsdjSnorCYhCmOWcxH54gLChB3fVLToKagQTMVJCljfjefm0MIePbPoD+Kv+318OM
T6kKBnJOEqiiwEi4Gy9MdsQt2nwJmWyZE8UO1e4/wzfm1d+r/VqrMr2n1rt2wYXZIhFkBTKDzVLh
h4MPGIfpw7vqf4jcQ0GVoUW3r/+1FCI071+7JEUeTwE96iBjk9NFe+QPF3bLkacVCM1Ugu0TAwvh
xoMJGUiC4UYazTmXI3nhdHZD2ZeJpcg0ZLNx2enZdt5CJ55EsM5jeiJB/xPnwci8fWS+HL1SNRmD
llPQWSAOdIP9ASfGU/Euu2rv+qhKDLrEQKXo0w7+7KRbB/vEG6FPq1Dy2MSPsCzocRfvhDgftJIK
wcPiFrJSpQRNqveG1PPt67knhOywI+jPQrzjQTwW5Hz0vI808KvxO4eTiplTEsqx2tfELvWP/vI3
NYNa4EdAUYRvT5PbL/+RiChOHyMHcIqF9cl28xyWFKoWBxrGZCh9KcIs437Vuohk2PYby+SA7b4X
toJETo0JLEOwdiQS3sfLFiS5UXVW9Ilqp0kbH9xXqt43UPi4ArjT/IVYLd4z10ljdk5AadXDGzCE
KLpLvbx+XTdWZWRvuE1X5GWwLG6Q51VMQg8kg/an+pT8e10t9k+WQuE/d/hPIGLzSkeElzxJ4iKy
tet1dVJluEXMqrijofgYlGM7uN/KczIsmapCo+Joq7RC2ekgzlmBkt8mqruOPd7dqBt+mXNF+R1G
NlrzVBW2qw+tmA/PLNRMoMDnpN1T93JtpOrVDcgJayJzM+g7N6vkFjNELlgez3Z0H6pZiZZ7RCOl
7xm5HnzgDqWZhXXw8mer4U84CkXVmK27JQ59bX1zyKJP6RthbD6eVAhvu0mvzlOBklcrGqephQOl
UhCxOs5E8DR7F/JEj2rpxgmgWjPbGdCwLVCCESb5LBV7L0vX6OuQBLoC8nWvXnPUWF+FJpmvVAPj
u/wGRj8ZPf3HtkayYkaHBvJwm9bTsID7z0UwrA51bE15aHwwJVYOMK1O5f9QB4CSLmLSutXa5X5N
MbbVP28j1mzcf9i5wbsk8BFykWbcMDhzLeph6nqrbYmPvQQ11tHE+QTIekpWgho3fjaPe+mNjqMz
YN1faVDxZhUuSZxF1EICbP3CoFljJQkIV7DBLwATpeD0m/L3TekSNMhAwhRrhJwhzqL8YX8HAI3g
yvC1Zi7vZQW+jlcGminn/MjDO/2T/7ANy7dk6Nx8fn/c3tynPNi3wFUK92o9IF32kbmTy3CaptWw
vn7VCPhMNj3zPOPy1BMgy2SsRZtfS6Bsm4yJjL7zlPoR3iEPjfAy8ywnwDel6W1KL6R7KocK5koO
Vd4C6d9h+zaF2E7I5/Xry9op3kBnqMYlK+MrZfpYB4q9EaTq7ajj4gt62lsrTslXK4SY8hE9ziWd
WS27YY8pkoptPatIgA7+Zt49RrcAAnxoFYFpLb98y8nDjmtktwFa82Zcf5E22zNly9FugoRwhhYK
nX0xklW4dmUKwY+PcllBljSQvwPnpjsu1gH5pouFTFmUVXLXqm5EM0B3FHEX8IKJ/bDP9dRZOttm
ew3QsqkKi2N0qGB1glj+Uw3g8iVfWq+zNBcIOHP/TGpQvosrRfUNrm7uF/BBTC+8GOgsEfmxm2y6
9y+EdxrYrmSgMANktDRWS4lh6HLN7fyYStdndYykXNf/U8ci4FV9GgtVpsq50s7N+jmZkrZ43lTv
rhQoikk6xJE8JhSeG9DZQa763fS/xrdyZ+KXW93KroN1c4cj3otW7dMR+tZ/YqEwkbkM62whis8u
ui0nUH0QXKt4NhxOG4RDjSirAwwWOD3AWSG1Sign4ATKOij1rcAi8eXQTihracYAQ3Gej1KQ2oka
RZm1IT76S0ZJuP+TFBYBlfYGoWMn4Npw3vvaoEz+kzlEAguTQuXfbb6uKMyx4k26rGUcIfqkSTMS
bfa3R4ixV4CJf8BM4nnZM+8BWwaOaxOwT7XevIDG8fWL7YjT2h/61pfXrdGHJCvwdd7kdF5Eeldc
2EoMV1g1pfWLyTnGxnZtNjfgkQaTvvuOPQHe+m69zXhjxQSf1WvwibnQRNvwSYE+D85S06R6nMwG
UQPcCRGwF8z15RN8iBQpbxd//HY8BJqUBQBCqS9EJJidJLqYVRVe3m7YOtOfFySvvSX2gJA9/aQ8
oFqYaITrrayYhsGrZ1RgNoGYYbNOKL0dXEXyzSAmPgPkEJaam+RHVZZaPr1vLFDvtvu+0Ybr1/wU
muQIlHkoygii+JJxdpmLdxnqvB+aBDRVJuHVfAcOo2tVpPb5uXX6o367lPrD+rVb5LdwsogIaobf
iJNGABHIiVPBOo39svsuYlJpOcJ/32sxM6ppaHh2Gp/lhCtNwJ46as/n5DqTgI3CkqJzIO5NgqFa
RpOqp2QYn1AiIf94oJ9wr78PzowyRUldeVcDvzQi/ok+tKsxuJwgqaF67rzrd/VwfA+TMd7Eel6S
g9cHOdnS5MD80fKS928c2nMQxa2gR/F0cgR+JaFjxMtC2F8OJOiRgEdxxbxD5S2FaPPcpohu1dYY
7zruGtnYEzCFcHzt1tn/o8OnspJU7TkyQ+oRB7KeLwqVZMQ5by6IkVHlL6XVrA3Ad+efF65aUHTY
vfHFOxMCs/3KR/r/LtNO8ZGuYE+6m6xJQQJUMV81fgRVAs18LWQ+LWTnPhzr+YIAYHNIz9AFJx69
Rwah02hggGcMJEopDU0zEuVgiGgVB5ls1gi4hteqyttxfqFYI1/DDgjXqrdZRCHJxUy20CX9cXvr
OpxlEGvkbJizj2xzV58nNu7B7qeQoaArBXI9L8YRYsqN2mOUnNMGteTspzUZwctQPkLOiobveAvm
bieQizF/oqbHuNOrMb/zatGUTiQyMYAxWWiNlDL0PMuHU6NHuDgzjYfYs6eHEL2p/1NN2LNyhAKv
PfrM52OqI8YBuvhsOJ3RB5TMiP3tDo8KFzfYqdx4MHwxAMUaQj3kR8XdB50xsBKv6gIlNtl101WK
L7lrqvazp5552PwYomt9rFB64H/E5gFTkMEugFVJyNKiNEXe0nZtYrf6BHdV7nYBkbmxkG56GhwG
bGon5210vhIb0LCahFzPPLgZWZuZf/9jC5V2W13wSZhQYv+MFlfg06gPB1MH0lSI9bKJ5SV6meFt
Drrqx//+uHzcm0D9J00d6PXuaX3gikYrnO3kdcxcr9IRIWTHNzfM/dt1ls3wVu1OjzkhRWmJwLqC
VaNwPu/8vMwabq0DIsZnuvacqE0eFPi+1deQmWmkZrb7KhZReNS/yRYn1CP7mAldNKRTWWmx87S2
8GyYUZDvNbrm9BTHVRLyHlGMfH6bbIHhlTSm8HNj1r9gp6bAKm0h+KL3RstBbWii1T86BPJbbGJs
/sqdI5mkLzJoF2WIXry8FpTuu1WGeSIC9MOF3lB/fUxdKD0VqgXXzoYUt4XaXsworsuzyyOygFqd
q097DJ5yS0KO+3/M08vIOtouNraTtA4wqA6iR7L8jJMx2XI4foelwQLsFmkDYjdEGrGixUGYebN9
szw3RLlK0/1cnk7n7e+BQOK38hYXxUR49PJ3fRVyZDQOwUCIg0VQe8j4rlsZJ2+dkVHLNyvhpvdo
nS/ghmnOvgprkGxsqefBT4Kb6WcS8PUS4Dse8WrEsuxzF0nGcgw2Wla9V6GF5uiGE7j4hnYXUhRN
YZctPD3k1Wd98qMBS59u60KyN/cfYf0RSm2vYvvsFTVFUcYDOdaIS5g+duo7YhseT3hLXkW5ezO4
x5S4cQD/6PscYZO9CsvQzcAfTsvqmc5slMtZ9720nGXwHEhkbQgkC0Qet4q2TcSYrhiN2OerxVXf
RpF8TzX23TPN7MItUY+OCjCS/yrAJYNjbuNKroIvUZKE38ZvlnraF+6Y5OCQh/mCcwFWFlvhBjw8
+kaFBVu1ko8mpA9vgmIyj4/VWf9otc2wVM0ksMXyE9kYNS7VKFQfikV5d+8Mx1/dstDJll2giFxw
rB0vvdQFmECh1cdmRZ9SQsEIPM7Ku70sDBJFpbTZSR2AZIcQjTZyZhUP6H+/mtLLbqladkvxTyzA
b54WWLUe+9N6kUVTcrtLSG3V7kqAzvL6by7RYI6ZM9H0WceA+5zc+OHEoLPTftaVne++4NA1E1rv
A8bkJnHwiZTSasaWSlHFTmwzPW5Q3wPmGodxNUdp3aPkTL48i1UF0ucgXjW19gUyharmRR9GVDW6
l5zr0mO4Jz46i57p+Jeh+CVYb/SF/oG7SNRduF07iBrLpYuknL7N9AQmQz2lFZFRCisUtrVxBWdf
g87ReSnyCD5Ca9EXIDBkrYhSdHmiS/gz+QViPinP09TnvzZJbWMpq1eVUbWODYnLuk9vGkOFVLnl
U+kNoOy26kXf4/297hto/UD28O2pWOByLuayLrdX1LTolKKDp7ejmqtH0usPtY6Hhxe531IxhvrH
o5ncm0iR+v5Yn2Ry0TOSweLFINXCSsol+FnaIkVtt1Hs0btYWe8Bf4mbJy8IiKJPFMnv9M+WSQch
HEx+2nS1dJ5CPpgV3699/e79I85eU6K+FEfBMELweEup+RDNGMrL4ASXl59DWIkJLBS3EGosil2E
jvAiqYypXY17A4PVu9Hk1G9hsWvYGlISc6gpmzMS5btlt4PFioJHOxleOmLvA3VaUsXR575Mprac
mNqQiUDafLD2aTvqDDEc6AbCqaJxc2L4xfwEye4eDgvc8R4bEo2QMcOdhg/ePz8+iMLw+qAKN/yZ
bwk2qj87hbyMxo7JbezwQsAYhk9WtMCJNusbcFgDX0ER2HP34bhOzYwnBYrQ13nSXdjxCGdLvNgy
oWEGAyXphsFxuMTCNwQm34Y7Eax0hyvGHmuz6rwkj7c7EsNQJhUfnkZNqZPYzDhqqaxjrASqxEgO
tlkvUC+I+VuUhn0nsImJPllRkdFvL9esefTvj4gJDyKWiiPzQLINuFJkZGP6hR/3D3sLj3iHz3g2
5TxH4ORomvAtqjQfvGiK34pJIWU5SL5PGHUX7fubdAN3hJdP6Qh1O+HKQwv51sHiW5RubR7FIbmm
A0s4nVJdS73iNka+WtZSzLdccbzSV30B/GN18ZxF7ApsdxhLe+MtEpBvKVs5rheACHEp9iya6jJP
5jVWWUpB+LATWLaMi6xSWCAJS+9oo7Tp/hhc3lpYZinGs2qn5Qm63pSHh4S3V8xIbr541Hu93/7q
gIruJjkdPl2VYAQvNtFTZsy9zlLVGifyJPPL6wwq6VC1+5RkLhq29ppCWhy+B/UBRlhlxdkD0CVt
M3UhyrOkCQC3KRmGc4BY5VMHOfscf1vi0+D89Zn4md2Q1iCglKRDyMpVjNo5z7EJI0fJORLlhlz+
yda/IgUkhjI0qCVS0JI/ILV7A7AXjpeDkto5rUQgiTz+uSwSk/wqwpUArtobDdT7zZF2d+lr8QdZ
13ri53wKrlKOrwxsu+DOZk3PSI66FK23mH9ctWYhdV7Z3lQuIvzPf20K2AbyPKmkJ54ymgcxmI32
5QUlrJs6V1QGa0rbMxekvEUPAV5tN6Tbax0T1wmkgkKEUT9r11MOcW3YUG26pNQqs/6ylzL4EYbK
7NiCh9f/LYRbMaq0oMFxG1gR9LjMjA/FjAl/qUhVkOYUclKpX9XscXye8QWkn1+1gVqPdszRfEeZ
+UCf4iPuydoEncCefeM/iJJ8GzGepUVP4syc1J2T7L3OgA7w5e/Uk4kD/W4tSx8Kk+JR6/uD9qzG
BZ8HW5ZOQKxbd7sDPfm23mHGoCxtRJ7sof93AlTpeVHgCIHtcyThxbRlf7Rhabe/Nm/5kaqczm5T
V0+GsQ2RaKTgnu6sboecfvP2YfHnnXnv1GM/lEZR3z3fT098D5UvPAlatXeILVHURbPC4/7DNF8R
RCOYJwLUF8aQ8+2frrb3hjmxVdQaR/51AmsvXKmkJFV1HimHSiayAcNbL3sHFJ6++/aBI9yhVPw5
YH91cEnWmKYTphzk5GV07RhDEpWVxQ4VgMPcMoH+gxcKVYiafbc7oa4YRHlFNUpc7tdzJTlAdaCU
FeO/IPXyDNnfvSqK2XzmbSLyk4zNFem5oZTbejQUENPhQd9qmh641Gn+stwFRQpS2KljVCJYfvhK
LdjtEhfsWZpZHA1NmBYQUd9w3Oo+g+OTS1fnzdJ3EKnHjCojffPMaa0brZcjxIB34/SebcpwAh/Q
m1yhuLxJwAziw4UsbdLU9cpdktehf8ImVz5oWZU17eS5d8HsbWtisNrfug380JCUm0/B7hfKiWWN
1GvDUlUIbwPJqxq8NP/hzv9LTeJItQIib9ZifYGZVLvqZm9IRDCqCUPObsY1EIP0OBl0G/VzTyBT
GZFdVtGxBloIiETV61IMHmBUSUTJWrWx07/w2xrKfHrU3P5dlIx1nMLZCqA2a4b0ybu1UGEXKYJE
dDTH+UWJl8nqw9yWc55IYWPoGteCju0UMaOly2OxNn+uCx4Eh8iYuakIfuxYUHz/R15XjTNn3pH+
9NqDbUc7d73L16cv5ReZg8Ph4H8HneVrCd8lr1eZF3MvQ4B+7np30TMYKNTJo4GsVIJD649xjSFf
UIDyAHE9r2NAaTGJz+wAO+Z+fG0buyMu4QRoTRAGlTFGRIMhZMH0JkdJRL3bdFUVQ5XPlel/kPda
LnMWPDWQT5dWz+jHmJOu7TArPsRdDhq+I8mTqRvJETT2WDlAOMWGXn/FUctFW5IO9GMAhpXYPwDi
G3Tsz8g4xIFJRrIuOtJcAy8MvSOHVmAA92cp5/SDzh6cg8k+j2iQ2wfBXPO0cFDjj6xket7R7Zic
n1sXneOf2O/GXH7xTYp6wVZkHy6Zcw8KXg00az/xvGaX7pu3uhxCH6t0C6l/vW7yBzDyCgQhKXFW
37rFSSHy1kfxOADYETHiDUpEXHhnogcVsQiyR3JvWvQhodLmHL7iSeaWof094nD5lEncXQFnmp64
0xEu/ZCB114yzYFJs6ERVVPjrwI5TPbOh9uzYMzRPUPvUOqAt2dNVLFS0Y2PbXK9FgYhmHz0ZQ2g
G3SfsTfyBfwZi92YNnhGnhg5sT//4eEo269bBJ37WmkG6lChUVQPIkUp/LorJMm1zBtxxwqSQNgz
jAtfh2tcl6lgA99MonDxlUSGXoQdicTv4tGsJfbUSiFGzc/xFqLP6krORLpHlmW14chaYewwwJr5
bvmQlFrVFLEy5EBJVDh4LLkGOBzkPHHlHLVAaNQYpXZUqK2I8OYJzy0M28S+HHLSTI9yoVrZ/AXg
EXuzXyfbIbWXHAMCYgpax/BloYzDXfkpfE/PDEPAK8y3nHbqM6+PPnCiX/Hr5A4p0ruEinY7to1U
RHWqUfZuc59jwyRzdX8eYSmfweWUdPogfy9gltKFA2P5q14o4xTH91tgz+B5k7vFWyt7DoTz/tq0
vW1U0HFB3N2uMIJjUHiXODycz6mHUeYZ3wnvQxaC0IkV5pCkQK+gp33lMwpnBbmlh6jtM96qqCH/
IUsdYY3K7pYF0i3kfSrtgTOrxTPUy4pjuZ0bBKwWcGif04Mot4cIA9McaFn8sEDoLqplhSQvnZvG
fDkvinMzfMRLQwR7K5e59g2IJJLPqEsUtwUeoBQaEfqFvKT/ot/m9MQQLto/V1RcqIDHvzsRsj64
fpWpKeNL+Dk6k6PWP39sQZlL4HC7+9gKWIxvZHhXU9W0ui7JVmiQt0fiyWVvIudPGA1L8z1KBK4D
pj/w+2vA8t0RcRNogjEceozfDQvDpuu0El99ezGvkf5cqcpP/VuXHziZOkweJvquFJO6QLaAull9
iLsBN3xAcztJTk+19W97a/QB3p8dvbf38hii6e7LhzONR2KTxXXKHKdkqt6IesW80o8mp0LMCpH5
+aYwfn4J58hrC9bxZPQ9C8KhqS7Be4/sSGCd8h3MVvDofTeolQQsjS87xsBWrJvotQwmwqAjzTGO
fPqmpzrd0T2WonPvzE4CFXe3+UlZStlQBboHddaqV2NMYJ0K0ohWTt/k3bQrP4pYb3rHrNF5uJ6C
qDnX21Sx7R71GDfKjNb7z4d3BhfU+FDX3ZGTkcWYcCrWfU7/awqRovN1FSIJuc4P+fZlVrXPgLz5
Z5ZYtuyJfL9H6dXvWXunreLRJqNvuBcKbntsw1wUT30f810RU0SF1oa11NGpyDdiPXyUSi2c+E7R
HWn17/8NZHlKH1FRDl2VhzxPRfG/pCswFrhrnZ53nXfaSLiGYrdrZdMIKRSNCE+MNAG/aKbcX4XC
LGgr3uoWweRmXJ6jd1TIzicxMVLOqu3lfso2HuLvTBca8NegrpBaF1gpVcGAL6V7f/1WW/aegKVQ
vvEGLVOeMdOfB/DLTls9xvJZvxYBBYPpXxRpZap8yfIZPLuV1QBF0scR/D4TRYRo2qyrxXTgIWPx
wf7FSms1Ne3VoLk9sOrSuYzEXF9ZzzIVGV2/M2gossj0xyvhJxj6+v9OK3qr96TAcSTexx/EaQJc
K+HwCPrPv/oWqS6FnTP1IUwplWGtUvEL9bAJyzIv4cnbw53s+qFASGmSwvKc0Ph0bgaKsIS2r7n4
bu3ixAJk+dp6ChyCisOC/pb9WlDYK+LUL6UlJHYbXgIHtOo+qpG1Ry0Z8/ZrEBHG8b+1RbXfdnvr
CePCXDs9697m6oagOe9vmOJqjKkj9kdcZw3vktYuE3N9PmTFe9ty0Wze8OJoXEl1sQJ0KqfRaSkd
wy+SNOMCALXvQeMouOZKVD8gqJCEJLIp5NKVFGcIMoOct7juUT84eBd15N2ahZUD0Br/uGjnAk0f
/HJB0Ij+9e2FY5RiJjyb7eELG7X3+qebCPjy3hVq2DarrhYC/xdrT/t2IokFMeVqrm/+dRih3V8x
Y0YbFxU+d8BrOtI187QOnw5MWS6W4rkeRQXQRlQj5dTCgyuEAFMB3Om9FIuTgRvS7cpS6uTqr+ga
yRfZUldi3MF7OJur0w6Ko2cc+B6QjkghTQdHlukYuNXn8OMDbKduPOeSlx3fwNDsjzQqCZrVrze3
v9Ag1zhVnWilCYNBUZ9Gx2SEAzE8Im/Va6Xz4JqCkIammYBZX6Gap2anTlO9W6c/7D/93mIVsFkf
2bcwnDumdDsWXC4aVruCRhDezd/9U3YU9NpguN/RIHAKz7KrjH0TuvDhZNDWRvJG+UihKhwhd3Iy
Qh7zkXFjkrJkT14Jhr7AXVXGLcLUTOuRvx3IHFCnnIbEpX7kPqwCYt8jk6VMo5EeTmLVyjnmIB7V
dVhq8nfSGyF04zr3l4Dt17H3BW6+AhLZRgB2Zdwh2ae16ImoZf3ZT+jMFYsiPmGVaxB6UC23f/DJ
hEPJ8LDA0ieEJU9Bw9AWzSEbxIAthtWCD6raPT+0wZ9j9xrtWkMkxM70X3znAZi+PnDSOv936fYT
Y0389+PWEBBfYj4thPcGb1odStob4g/J+sow6qeqWP1aMIZhJr1qr9x74EpV2Bel0Mvad5EkZ7uO
kKPLMFGsPNpC1Iw8minuCUOcpjRvqIEhjNOXVF6rvsDROgP9qO+4jZDMoUB1CdZ/8jzEuDNg1rd6
JC7ZKWMF7mkY8OPhipy8UyR0NA/iuPrfCuMykQwTl+PWNKOS7mhBtCJAER4ap239z+9cM47Kbkgx
KutYKOvtzwxUYXcEUYe2b4P1ZZk1ubHQJYQ7GpMUy1P5byOlJj95ACydEMDu+vHWKZUFfGkZmirz
NbcVOxZ1BY/PM16ZLrQQMm7g7BN4yxXW/vhwE2X3+wQqV2UeBISY0G02wtALj/LKwkFL6CsQMExy
6mAIqPxaZIBETUC+sP/JOs6bp1GXijqftC9skuLcoFzEh4ybhr7n++HUQ0XfSrmiiGJVVyUri7vX
u7JUZyJAIXfQ7BikxFjKojZnfahJsoKB8eeOK9sb3BXbtuHQOvBPaaB8VQijgjUcGgQrHwJELx1L
dxiUcIuoDQLGZIG8s5MwZ81TMb5VPj8wN3iCFGBGhLP+XlVcle9tfbUvsRcnMhVL2/iFl3K/RQ7k
Wm+tgwJelwYTsfOkXuOzTwgIxgGmT9n1jBAuIP+ZXD5nchRvbaCmTjBfNz18TOCyGYiSqXEgQQVx
hrEBGqCj3DVB8Ixna7SqeJRkzcd+EBYphG9z6T7wLEP/w594JzrzDmzERGcQxumZixjtdpzHrpg3
dvokBknrVTQdVg021bBFTi1mKxkn+PjCnTphI1Fbtb926Y/aTb3VKG3SUXINoJOpwF2BMWYzGahf
LNQFrusjaDpVzw+vZ6L3r2D2UongHJu9ymQkETFeK+ukEweDFV6IxAm21pDLab9yfkxYXG4Sh5S8
nFj8Maw9y1bQigEY4sS6psCCFvErJ4Z5e+CYfw8+J21kYKbsaF7bPt6nD4+spwsk537BineMfRqW
ZmdyQhdjGgUUQ/RKupXvm40B2GkPdlpq2F1+NofHFpUzmhWYC8fHood4rZZQv/Y7WAEeXeZRH7Ij
wN5XvruYVbPp6EWPpF5imYwWmFGv1gOXpT1IhGpbUpfE5y6BTeKX921/apCOZbhVUquBc01g6XZe
cxmpaVvtHGd610FfC2qmfavkkjYOas8ErAqroLSaKdIUkLnxVLoF5tiDD3cecvZuvgvq5wO14Q86
m2mz1V8dJtiBsUlkPQ7mszrnSJVWgCGyRxpbjADwKURT7VO9AdmclnfUV5+VzYeQjlQQV6tfyEPF
O5kZjsorOrjMPHdLs8N4p+Vdh+k3kfQaDxWIPHGhGdRYJYzK4mvrRol0chA38CDfthQGhsTMAn2y
C9h8hbJuI0ABvag0T6x80hwikBJ8XWAvK1KQYDSdUwTif79lzZ1X9DVhUkXtQMhoTx+yxQm/IECc
K0dS20hFGabb2/oypvP+2PVV/HtfnHzlqBxct36QwP9OK62dx04XjI6mnrZHXKJ8FdVw4ow9Y9KO
tmoHeXmnvQJ+Igl1DikoBY8bxH36z2QRw+yPm8+E5EZ5OF5SmxZIkIN+FoflmPP/7cXE+Xw1BQFv
KybVSZWyoxswXcTIFO0nw39Tc6bvarw8wWLxhOqQKAxQMoGUQY/JxFYnChPd09rTZjHAj+gGvgYr
+iD2bS+ojZIlS3GPh9wnI8VAItWtLTv6oppvOl1wCELPBT+V2d9X55XAaeTEIxRCNrhfXUTXPbXP
OWYC/BFimMeqA8UHvsjQcxZIVLkqPc0Oth0aPUk2Pj0U7+NDplLxgHBnWyMnN6h+gOUcaEk31kpt
YSO7E/VShX3+js7e5a+jE5ZwNfElKth8ABjhQjoUBQ4Crl5AP3MdNDAeJteOkEa2SYLUBK9es6Tm
ugReCA/zOl8VqHGvCAxTBDDCCvC967xJCX082IFbiCNxpok7IfKLzw9Q1LNgOIBq2M3ridJ2aqLy
X2juXS8GHNQT+jAO58AZVehytmXljAElziSSNx/8VtvHKFzm0tNCL9CMlJk6dIaMAocgkmR6U3Bt
eOxQ4MXQaYnL2f64fgte8bMv9SI0jg8Juv9syTI4BrhldP0j1PtSrjmQ1AdzieEW9gXFXBGadNFB
c3p3oXNeP1MpSKOQlTCyfQAEMZv5x1EB8CrDeMGDLscvdz4ZB/WOLErnAkj0SBiiuInlSGGaCeSz
jbpvPe2G6jzXG4VeFMwKirY2azx3CC6J9YxiXDVj2bR0ZxNgOgQXoyVIOxqvMQQ3DvyhIXcnvsny
TXrxFWdP+xw+Hid2LpkXwQGSBamQLsE0bcFE8fduwZTyOhmIiX94ythAmfmnL3PyiaLNWOw1Fz3b
n2Fo+wdKPNSe7H/5J2/Xj1UNs09d5CwUgpJXVONwZcdvhZ2h7v4nGtV9VzrqKpes1Nj3neIEnMFH
3cQbjBgrV0ru9yNGUdBI6f4+iKvQvFVG1Z6ASrLsFpskv3lTEbbZnkpUbd4OoD7HmzwtAvBprBoj
lck0h+5z9RSUB2vpC2MQsahIxVFZYbCtaY9Jy/6ad8RPE6h8GGrPjWMib8EVTHHFFeRbLZnJD8XI
p2I7StU/I7hQvnFA9C2Pod1Qhel0nPUUKfcadppQ6eNLRbo2O1e6DEaqg9/nCaz/ejpbyEYpadlB
qMLSJipUkuGufwfV2l9wOVjiwTEepHI1f00axPz0wz/LDRkIF2Scm/hJkPXPHwKiv9ML0cFq/AfZ
rmZDbZfKJQQj9E2RCl36b7dtdn7pkQQOv3YL6HvEtgLl07TPltbyAXYfDMMbBqtBwEufWGxvw7n7
u7NWtu2sqUpjFhmDMp9KhL4+U0GDAA/axz99ltJTh4T19OpcCjWLWLqJRWaFrXdyzgI77Hq5PF/V
KIzvJx9st5ma6b/iA4iKifaIu4P70ccXQ1ZlVwGNwyqFJ7weAt1k2Ey2KvuXgwBrHSG4YSeF9o91
iakmii4yZuEpfUHtb3eOh4ZeFd4wumPmZNYQuQF6xQzdCCajNRlLt7FpqOx4nWHJhEuYQmdPjqJr
6gR7xqOxlljPXE0zDKGl65prZbN0rcqOlXNT4uJxOS5DSjnaMxbrXlmmE1HV5Y8/8bpIj4Z7JTGY
4JtbaZ6rOTohK+/JrrO7QSIblRrPffxn1WnftibNZ+HCGO/N+xq9Z69cR6vIqnLiF+OXpD1Q9O9f
6jJRJhItyL86XSbbHdOkw6Xl85V0sl1tgqMf/7SFXeu71vDXsY/Mbr5gCyx57KBOQvX6+GTujjkh
orjCfh72pABnrVxY9vPyXjRUBQNQZ4yqKIKiVz0m6tncpf3XJ+35nRflIP0BM/zH6n2auuVwWi4E
SZsxtzi4Ei1v3GDJb314Ul7eiNRoH9DfX8ibpJVzUFfnEBSKriCkNumpXyzeJz0PKupn/GzoLL39
soUJ5tBGN8fJgIvxhDadtS87PbzbArI8ZDHQvS+J0ztuIqFNdc2Rx0maoDQd83ZhXSx8Z78cVmKj
L9r/1pj+oLjY5i3T6HXl/9ukPLLftnriHnKU4Djl8qhCwcKVxSUwMbH/WDiE3nSqzOUIZOMOFwD+
uSiQQtuEOJwZoSi8wMKt+C6R7FR6WoE75lKO1TlDkk1oWmpZxOmMDNvKvdxfrOppaCJv1gdQ4KK1
/YyOHElHwExx28l971ydiGhOOU8Tc6cRz0xdQmx7PTIbdCNp27lgsHwedMV+RExqfQYOPLDlEuUB
tzkl7ZrqmlbHr6TpdYdtmnVz+ht/4fheiubKcc71QHR7rmJudTmppudpTV5D52TQfrxvDgF9hmfs
qxBQ3Bw8PMIOYrdbX7nmDEvUp4p13APItZ94ShbSVIcX/p+Sue010WcySS10HjDxVpjMfr1L3+Kc
CU/2uqq6n5B1mefYrE2KDSDrHrWMG+bpiYYQf2+2s7WqVX+cKDStuYMh0Zlv+o2h+OORo8xx7v4K
gPrxiTGO2XpYphgApcbixols6lT8zrUadlJVZ+I7/HnRVuyY0ezTbWZD3AyI7auINJNhYZwXOVLB
a4+TXV3CdeRNlk6ztZYInQz7GoXiIq75E1vYyfaeyOqUeYewO8pWolE1wZmOYZQNjJ4oCcfo61o5
uRn38g1KJ15PSrDVwLNrp9XVmRHggpBOpwTq70K55qmTHGGkX6OE0F/RP6F1VqT7Iq0gIs50Vxgo
CCjsXQ/2JkM8jbSr9SV7VaPtH9gnyJOMkVA6b5eZwPs0PXNcIFWXPv7A5RnZ+qETXVHxVJN0t/rj
ru/w+MrkYwUDhyL1cqeE9K8JP5aN5doYEBDIeUw2Dhi+wASrzJwlo6Sj8nc/Z3q13q5Rxdk0NpUz
V0zFL1PTE/GSMPIZCgBQhRTAen5ibaA79sE6VCni29kMub2rvH7Axin+USpc+q1woI9v7QwDh7iD
+pxCSBoAJzvDASG0nRloLyX4U9QwApIK88qiTVp1V5gDV30g08X7VwosIj2HxaBVtc9AJUVqYku3
BizeeiDohWogfStV/5RPuLiPa1DkwIeTWbhU2FlTNinO4qoHr8phxn82j8v6dhriq8JUEfhteieZ
7oY2ckEqudLRJvDRX8J8q/5QqmUUIMyqjfknfwuhQha77zqloMLmEKxurDpmiWA9MAH8FLVD6gsL
tNDZW5XUsJdZd7xH/SrKBiww6AMvp45SQswwMhSd+IxDcpaEtNHemRsrjQv5KMr2jotSXTsSh65d
zyx8hIzgK/9nWJmErPxTr2vroYh1JVNxAAgQKjCSQ2kPdgKoqEdrEPv2JJbAWXVIV/Fo/1EV3U4i
TDL19yoZUJTk6RvtWwKa5zK33UuXJp2w+yLcT3Ec9NKLghA/IUgN45GkFJHc7TU1aXWXhVfatV0o
AMrK3e7kN70VEtU95MDOfIxNgZ0cT1rahToMTUU3LQz8oXcoXfaWlUrDbHnYQRqmAY3wSA4wMn2p
MrP4Tv1krAr5F0IUJEL89rbXROyZ5n5TXDRLZoVBj8az+fPbiDvrJivTVa1jad/OB2y1I6lRj7jf
xIyPSlg9njMzAZKxuKUXu6GQXA6zBmmHILSpDAS28AUjDnKxGNUWCsVQ2e1D6dPjNRFCytxKIaFw
ZAnooQb9lRj3+o9LuXs2QvYu09CqV6b8uyprrlbJgxAFDHqy2V2py33czw+rTt6kVAhgrSsl8dFx
9Dbo/gSv4q887IE377sJVO26pGcEAHt4pTALTOIkKyE8/9U9+5o1gNa0OKj4kDwdtwIP0CRcz9RO
Jxm/Xm+MvcaZnl3Ve5D8VtMSRLT/O1i0HXMaRwa4X14SpYDE74CnHWpPs82Hl/GvJ3oZ5Rh3GS7k
7nI/5NVacOr1UK1hNI+mHaPANxlkYrga0wsJqEiHN19O7o65JaLMnT06xjCQxspkOLY86MlVS+qO
4WJVzAC4Rw7sAswZ4WZXS+e++nAucK/bWRRVnLEmavURdUezmxrffcv7NeaQIR+BlIZn+ogu9xRQ
DJufmX3K/g1g1I0KHBHoiDgZwBzQV+HUIi2mG0WXSvXqnAOzzrgxSJESeAAOH7y8lF4JXnwHAsnU
nwTyUk1BkiQQKifQO11pChy2Nw+NCutl7skGVrS01a/F6Fh1A3Uq9mW3E8d5raKt++RVx6l/xetr
UfM+a+97+/yQpeiCPRCtQBwfHBEsaKQQiUt0khGqAHM+Rq03ZTBjZNWwS1qx7IgSfL3Jm/3Gz/Uh
HR02HqhyUdrm6SPdd8E9ry33d9jRxztCNkffXO95d+CPWSNk/gQRMoVbH2onqXHZyrhiPTn5yjYP
bLLKximvGgXVpDfCN6D00Nhh+thl/8/B1iDLq2D0Sxn7Kpj7Q+fxD/nXOa3ef/dy5ON2Nfj+zK+y
1Yn7C7xWpK5jAgQJI3IxIZ5YrL/D6HwFjkMJeO0DuWmGb0dcCP1SWaQ3jS5dCzVV6vmuiDY41+nc
AGLjfCJte7k1yQq9ZZSeVKN3Ulp/1weiNpKpITO11TRt1NtdZ8PA7jV632KgzEMEzNB7JtcFZlAU
TrHlC7NwcbXhS8syo/kY1YUYsQxqmRXu5YmfFDlI7FtPTkQfOR1ZWJg5H3wnNXwYiskFq6ZmkcHU
cW4FvifLhMUytOnxAz16Kv53SoN4lEGVEn6ANr8upcj8M9L71qTGUOpXvuEgZ8Jr3ibAepplFyOi
owITqsLZFkvfSrmUbiMNDryg+6e4WT/0dX3niYtRNhYqLb/6XXIaKD6VvKZJeOGXGTNdxvyTrgVt
dMaoJiwJmSX8ThPYS/9B3B232KCZmXpYxQ84/PYYpjBO06gHxq1iFAXPimAY7VMO0Nlqib1SMa8L
agSOFWC3xbAoMj60zqfeqHRFmKISH9527eQTeAQHD3j7Ejc3UMb8i/okLgrFx2WNqAahxMrKL5RQ
Oilm7Z8P3rmKLcm0kbBiwCp+7KIIOpNsw0HPFFgfuLjVjXeeQXyBk44A6he7rR9+c4Sx3mWehg2H
MWPU98+MzBwjlxvoGLtDmikGDkCkQW+UmDeqDrffWHGxOsHRWhMY+BFYVrl7QOBV9tU8+knYRNd6
k5sYfvSGC0HsQ+zBo9Eofp/XMjh72UAzDuiuPdqfNMwHq1bN3Qu/05adQi+nkD95jgkC4IH9aNO7
jUYXsZTjX9IGqVj2a948FRbpR02JnWcj6gi3JT+xYJgxXG/yo77gZm0PEfVx+sxJgS+gXx1RdPQk
D+cwrI0GSazRzMknwCgyon9y9ChodXkkga4uxub1TX7ygQ4Bzuh6vNPFGZey1Kllb9pUipurllkl
GReMAgZ0ldQunyL9rKn0mLows4YjyhWvnVS0mzbgBPPGceBhJMVhwFKyD+D7cTYEB6UUung2Exwd
w45xcWRk3eZ/NjXBxV2Cd42DVaSQ61xe81cnVDTN8sLZ3Y1Qhavj1nRdcrh5o712BEUWUcq6u6Rw
v++vZyZLxJkh0wH8lF9aqpNyGA+3oXJR/SVGf0iA5Yg8wpUosUzC2TD4DZ9KYYg9bb6IAWMi+QE5
pAHUGTxkSUUCgqu/dL2jQkvNuFwb59CNBGJLzX2/SCIZYQf8g9sgMxPlI2yv+nmJLLjlgUmXC+Kt
5IvBWy0FgT83Ktzbs2EYB2dpS/6sXIJkR59pbPg2T3th0WLzRL6wZ0bpbpRJlPHcKwCeCIxGn4Sd
9UVZTO9XGJ+eZtSrTFvrMUEjOGnfAvwNvJVluwJswmDqq5CAcdkxWMz5mo0etXcpUZ65BNnoGDNr
sZDPlZ9LhH0W001v5ZcykZKJ2oGCem3WyE+8Ypt7gjcimvkOHSQlDwNfg5AI3opHuH1EGIExSzbc
YC3XFMMGb8CxngJsBud3YgpUtlv2OlzoH4ovLk9F18m6mQAcW0nQTPAPaFA2RGDZyCFx0kQLgTCJ
Q0uT1DYKdVfq5J6kKlnFRxi7juqTRVAe3ZBPuE3C/eRR778ZaGi3kI/ieMPYWQ52/iNxnuwVfcnP
MXLptAHENRBwotaaDqHY43/DRDAXXfZlQdJNt7lcgvWjVIi0X1s345dDCufmQ9fP20mTsJXKAXQD
lxgO92ZDIk6gh9PTJvd6fdY2bLwRwklZ89udkfutlY5BLcy47JJ9m3+rdezoepy7/dIBqf3Bt3yV
7DChS/9QKNGfM3yxDqWwNwFs2gsBBMaxUA7KJhpJA6Q2Ap9oF51DMX3qA/N8v+auYKSXqqoo8Y+7
xayxwM9OxOZeQT0n9BcZTEEjmOqk1J2XyB2ZukyLvPecLyzIAeyuAtweHzkUUecASggx4/47cAko
IC0Veim7MHmkUuZwqUgZ1Bb5nWrX6yB6ZjPdmQVWRRBZ1T7OoF788tZUnp56/5t1kKXQ9WMvE/04
SIjN9gMr+0UphXlM0qf65I7WKfhC3Qh7qFWi/GhLJ46Em9MkHaDs590ndZKwVMXH/Tw75SwYD4nm
MlgXkx99YMidNbAe0XCDzSaFtMVPy9zL8HKIvjgJ6TkOHXknnaXKyLlMecSzv5o8IynaZJKot2e5
D4NYwn+vCtmvQm9mk3cn6Ja+DhohRdzAPzUB+ZOELXpw+UAdmw/qH1kUE+SaeEq/4UUB0Xv8tJ2w
pq0ecPVfhfgkcSD7GnhsH6FK46aDGv5Xymk5N6frcQRy6SCDMBUxGC0H3iWwK4e9WpTwE6fyYwg1
0IoLOnuXQGehLeJBH9yvXrhy5IKl2y32pS8RMUaiGDUhNfJmTVAHNkOe8d0guHkjuPdy3AfYv+XU
msasi72gMSPE/+PlVKrpGwOqhpB55R7eY6DYPrhotvMKqFcpkS/1BKHdVX1TGUiEEW1ZH60HkUHI
sNSUEHHYTIjM4nSPw60RfPQ5SBPg0Vkhi9WLjwUADPJlsR9/1J0AtW3XqvAOGnhM+U8zrePB44sm
ihSwkz3aFxkCJOIVY0dkwL9HzB6bmDPwwCoNl7GkaFxuRR/AtRj05JAqT1qbXPR2itnaqqygOQqe
02uOgC4onVdCqhDPoYzOUqGEpcV7j5WFf5kYtPZNWbZVcchb/ymCuydunw8ndrjNaYG6VOkJxsQz
1CY7oE2nElz0zQp5LuV0ZxZEjXicpcJVf4MqBYr+GMbUIaGfJOoHW/fERpt2UmKzsxGpXriuqKI+
u+KrYOnbG32DUJDY3aaoIRNmXejmpJjhThhUhRvLhqsPqutBLPEkMrnJNN6F+sekdgW0/hdKqkM+
Eq8O6uEDD5NYFTqkYr1536VwBaCXoKJTAi0tIAgVDnQKC9LapgtpSpiU56Yu9FZU2UAzpkkbsbhY
G54EIR4hQJulOOSbkIeLMiuxtJ/iCL/6xrc+eS3jO3GbX9m/OJ6r5VPQJtqzVE1qMK8xScsyvFoy
6T8OqjD10INqc5r/Cj0zdkIdNEMND5cFdsgu9K1OjDyJi20LnTtXA4dBZdFq65oK4NX+sE+31YeR
GQ867GM1hEo03BY4uftK1mYoT49F5bKrlCj0vR1t7ew9rrVkPsT7cG3QVRX1j14e0YJ/KWIy9rIo
09rVWklggr9T1MXIbABQNAI4Y1iQyc+7yJjo8oiSUAePBa177s/+GUIKdCDSSst8z87g3+3SquS8
o4artnciGC2uJrrJxGgk6DIeK5aLWykm8I8ejqcU2LXVcuUAmqaaVaWxR1TVN4pqCBBfV72W1Gey
h4m/9p18zB9q4gKFKrV6VNnI3eC62CQ0hOxIlcbL2SP06xos/Rp1EbDStSks9CoOhS4dUaKjd8FY
3FUcQxpOa7KaigOciOSfpoPoMPl+aRsfpGzJUTdCPOUaIEVCrL9fe33YAEkNbwDQYdp6Lez3NH9m
xUAuM248CRTRukwr6k3PshRg/XECvC5aoCgF8mMdCyw4eTyCIm2bDZy1ges6OaNe5zStcIzXPzv8
GMuuukHPWYuZXEfFM37yMzCS2h29m+ff8jun+MDqiPB4lUjWU+axDyd+jD8fl2JpcjrMqxiCua40
4i1Int8h339JKMTgRomSJgWVGMZwICu5xNNGtuXCKjGgY5HqWZTN92iI6WghQAtDHSde1RoUX4Lj
5BqTul0hl93XU5dabQ35FdeHts9kxMx249Z8z5EvbsEXkGXnRRrI0goS4k49wjpClqplfZb5E8lF
Z02beRF4MfDoifxX2lZcw2hyjICUSvWPT9UGnakRY7vbTAxNB99t0owNQtVop+KG9gX2pw5a7sWY
uFFj1k4hBheTcg0C/hOUwx+pa1ILt+EYbqN+B3YHCc25Vqak0oC0KSUL91QqKVbnw4zzqEDOhO1/
lJzwYqEiObOqGbcoTCAwdrmfFb4II108DVdsUCoSKMH58Jwm/EOPUUxkY05mCnfTY9VPCauHEMs/
4qr4g0ZKlb5eqsMZ+oGJq1fifYX6PPO8fD26SKiXMxwMDTCCh5qWMJHT5YTm8PESglGORbpcepuc
aE2ED46jzQd7hh+5ep6lLahPqgTED9ECDGgfeINZ+pBFy83K1ZsfNKXOxvtFfGBvnN8jmpqoUdVR
Op6IDvR403z3qKsetBNZXfGsIpRVCFTyIRLyxy+4Rmxzlodsf4QPNd3KLR9D08620VELBXzDzzIo
9WbpJi70TbPvqQ9y4DXFRLFwnKqJ3fUp3llc2c1842cQ+nIr8qRkYCG3ixekDXsGUsMxL7EwGrXn
M+hMJGFnITPx5pjgdyImzGslunv975Rdc0p0yZw8RvXuJZ+oGZf/lTpu8q/v23h4nYYnuLoOTsUo
SDQ7F1Qlex700EPtQ95Odh/e8q5lF3pGhwQrkp/pUPsCo4UFEIRhKg4gufA31EJWrS0EjNifi6VX
QZclXl/Eq1BZ5u2YjQuH2vlRzwIgjPf0R1mTynyIeu2UrBhR4YeHlEmx7kmDeyOsSbc0DQT90KAj
5Xk4fIzm18nyY2ZQJoTFx/VtbAhhaLj9kgFUdIROOcpCrEMfd5HR/DC5M3qwnvKEohM11Jki5LtF
l5fDC45xiRJtUMuEQXNuI4Vt1gJD8aSGS00ApFLIs6MN9O6vPl+J1ZuidRUrAR95sf9sb+vPMq5C
mGUxBwNLInKh6YYqNm6c4tBIfOcB3bhtEDtLXwWtCASM6ZDtEf32Tr7hQqn13FsBIopUGc9UKxTs
4qkRY3iQ/AMPaFLTKZpCjHdRIMXELLUXoEv8gmrvK4HykJEbrRhYptcGeXTguFCdWaKlhD5SZGcm
ZszaqpPYZjOhbvlZTF2xjMYTpxY3MaAyZIAo2qBIE+zOXdlyvyH7hRtHGC6b1JwGSckyogCnt4xK
5LtF0OeXhf6FJL5LNvTgw9HcqNaJw1D1fYuoXC6u8uX0NtjAmM9hUkUKbBBBGSFygKUC1x2nbuud
siYbvQWky4IVC50OPloVcKUK1Phf3J9X9EL8LlvfpN+Rjg5d9yxrqI8ytRrukEIx2Ca5EOwJ2aI1
CPDP1FYNqYkdAps2Q2ErXi8bJq81gQHcGS57dSviuxXtM2vtF9CfjaUIN0fCPjmV+NNiOvP8kwdI
QXi2lXO23iXj5yh7+s1ROS3/nW37N/yv7HQeLSQdRwiW9TvQ/sxhpZyohitS9WBxAWxMiYfNNoRn
oV9wd2d3BrxJEKsCMkCLCEEzLvx2Tpa4mCIKSwjFwlI/Tnz0OUyn/V9lDkgrvUphUIjAnCeGypKK
xfdtHpjRYLPxZAd/BphZWM2Qy6Fmwvxjn8Upmc8AU2De9Nj2xU8+s0mbOPFTZ9WB/thcQDqEJG2Y
vFRrML7h3Av8Y76OICrK3kLNzj4ltNgRV6SVEw91oMaS19YwzvQe4/fNIP1be+qeA+RExF5UJ61D
CtLbWWZVWyFWoXaRPm6Gudv+legd8tUivmRBnW8PlhT0SRV8JwqdWjNvjPO+he+BcHg+gB6Fwhg4
AkXIvRGEfV5y4AfcJG4+iZE5MGHLp5NaeqPYfYetg8aG3K8y76uUs85OPpN0pne7RGgYG/ER1161
se/cCxKijRhgbKRV3PdDyDOfJUW3p/iY3CDCaV3VNvyu/Rkz+Pfx91+J5DdksNQg23QRWk6ARyxZ
WaF+58C4P3m8zwiGTCvu7QDdOnMPpfAPdnJPoBYlFP7Y4YWxHa2YVtClSV5cNGA+zIIKLQK1UU/j
FTTKPQy3biS0yU1i/k81mGrzAJph5vEDV4nbP9L3NtwePgXP3C6c+7xGuPaqCtoWa9vAMhEH/aj3
/yd5iIDfVsjsMbYUeKEs21pIJo6R++Aa1/jTz0ZtQEIqoKI33PHSs91NT+5MisORk2GwnRbTIwp8
XVdoDIjYoi/q8A4XATYfn09zRHGj/rmeZ2cBZi3Q/Zh43Cu70J7UODLneQg0xFriZKfS+1g9A2tJ
jCXH6gUbWmYyyISDaoZmLa6wQcAZJEJScnVtqOJrpC+0mgzpEkjPpqJLXmUSr1NQthQPGpQEYenq
f7Cfp8EujpGkSeAisaJm1ZYkoUl/H7j4PnoO634QG9l/wJVfK9L/TldSXIzgc/OC7LHrjBEmvwSE
nVhwWBBhymXoJ9/dtmcSpvu5DSiopYZwZbJQ4sKVeuA2HMFBrfU309JTOsjur80xLAoB8pu9ceJQ
4MRJi5rWTnAY2j5Ra8PDFfYF8kB7axV7CS1YVqwa48UaOaj1v0Pp7c9IWVDWRWBbupjLbLupEIAW
uD8LqU53waMPvrckFeOkHCB4msybaQlKr5scA9j1ZJzYlM14fRXB6vmi2NHJtvd7q7qfn/RKJQOX
pu0qXHXyFWFXq0jpm6b8bGbBCOgTvNLyf5164Cj66z4Fe0JnqzGy0d0WZhhjH8nFYriMS1yKEVYl
kZTWmyW5/KdwJdimsDwg1h72AdLKaikgcRUKEDt6XtSJmhZ5o2PaYj9oYQJHG9AK86GN2wTASG17
kHAnl9+XXUEPjBmY1v3APSHzKIu0Xo5HGnXkPT1Hkc+tO1dTlW4ifwa1iZ8qf8KT31LbTWHvZ6pR
QXhDc60NLDwhlTsaIFJF8g2iVVhHGGqz2cSs8/Dvlk2UNqx6DIwGmrCzPRVx2f4/verVnsuKtLY2
2MrmEsNhEsfU+43UPUyJiWnbSC4J/rjbnTUowSCILdz3mMG6vQ6fWq5CfL481ECb9Fk7K7BgP5w6
VGWbrcu4FkZZSeB3Wfh0H2QZCjiIHBljI3BoShCmCQYhdD1mjxQkjNbuYhT14PODu9KOzoQLaJ1N
DOYh3qvuC6q+b90dMHRrrzYdYqA3Z5PtY91nkvH2b27n0jLPLP/m2tLTD10b1kOjz2xeMSTPbll3
y8ISqdd23Uc2H/cbw8HI4b6ogPNwkori4fZaqRNTOAoMW/IR3Us5z25SZtbveB3UQ+SQ/wej4yFR
AvpmdG1DWp3pr6TFou16KIKpUSOBOp1MVwwdFUslrkT9f9E0IFQqjCaA4JxpEYjfq0Hy5CWDZkow
GR992Yzs2/dkc0BWhIFpnLkEQWmP3Wl+NcLp25LFn/T8dDfqe/HznszVPTMjkGfWgWxN9u9geYYT
0Bgcem4vMV7sRd7Rn94zzBZ+v/YXg8e1Smavxj0fGoiNG6l0vDx7DqyzKsX8XwXcrashRIHLyp8C
IO0Jp+hljzjt3MURJc4p3t8k4rcWs3ijYwKHSj9bi3sJEKberFPgD035W69tmSEpw/+SYIbHCBs9
HBiZAWMODBbX/aGs6h3J8jzo6unwhP7b5Z8BZLLfpzGQPU9Lmovw1gg+mw+wWNeBAAA5CLQvK1bv
Q+FDbUrTvRIRqtwvTRIflEolVeGG4sKY/aKMini9lWxtywTl3L8BBMBjXKiLzMBcG9h4Dgn6VEu2
FuOw5H72DM46EjQ9QcTJcrXplwitkwjatCBK4ii2IXTrVaB3Y5lJb2/JPgWJx6z6+cwqqPQel2r1
VexBkqfQjYbfz7/jjII+Pgi0qqUPQeiodhYEjG0KKiv7ajJ3lTdOzwzXPjtYVdW0hqLWibbMTnNb
/eod41KX0qO6xHPtXX+Il5PUjqTAYu/wx8wWcPzhkswhq3GM6NrR13qkdJrAFb4cEzT7+2hW09dg
iUL3u9jZXLAhFVbUbgDfKoA8ftxUmTep6lbzNVEz8NXdGVfZhSRHhfoD9sumLHTA/MDhZ+HFO0Ee
7u+rCIZqWknykzCsA/qVvhjCio5zZZ1i8rSJQHnDHQkfbcbrBTQRzIhcTnaYE1FBhIfdhqk6OkIY
lr7Q66zpwANZe4bfI3ZCHCDHFVqM0NEYXu8MVGlJ0Qmx/uRYO2l2yehqn0x2jNLIG55lffaNXgHy
waloSfCPT7nx6tI8HivEDas9L3h6mJyOTK8j2If3Xntr2cn9IJwXESXkF+hOCmWEmd8iAdKKGk2q
iGpjgplkUt6ppsEUNhw0dNm/qr11v7EmdTYmt56ASmeVHWp3wHBYqYjAHO0RrBXFCgeWxqpUGsJ6
GkYn0Ayzj11eiTMOmIDzWzFjAUudwYn5Q9EuWOcC0lx8qdymmNDeL3vvTw3W5HeWUOqYlcOk/lin
B1sS7TMNq2mrzC58nfZBwvIdecSbOF5mSC0udh6tdDjQMfzlr61YHafT4Yv13DTDFatol/yKVk+x
Ht44DTZmwghCBxY0ubAIhcoUoCk2EOOIpVC8Vl/yV6ZGtjfl82vCdd9ZdiAMblEZm+umI6zP/wKf
tWPxvZuY8GM0JQJ5b1DjhY094L0FB2HZpe3l9chBai0TNPvqfc0HgiorgIhdC5WnydOALLMQMrXH
5tY3jxfIt6BQL9vSbzfnD0wpQC2Zcg4rwFU5BQ13BLZXPosPUTkErVPOtd63rCfFp2Vz9Oc53AwO
eHATH8Scw481Lnnhkk1NhThQ1o5R4Un6iSjMZD3lm+VrZwvkGD1YtGCHC3DtV38KF+qPGsJizS3U
FF1CT/QCXczWf1+XH0LCWWujmZQ9SPoyHKOsKsLSBjVpYGDQ6E7YLCCqAxG0Z/j9uFry06E7dPmF
C2amPuG87MDzz0P0Jc5VMR/jZfOtUylGPsxUoRzibhrKEmvUJTJBS7xBU6CwsI/oqCVUl444jVDh
cTWDSj2P9mhcuo2EIguGzqZAgfvFHFxpPhjYDsgh5u7eRT22+eKxYQodE85ppKW3IZfuhIkWIxR+
Jk8OMIlAsM7gToB3peqiY8iEhDKvmjaHEKgowi0Yt9iP9vDwMkitTwNR4Pj6k47vzft4I8kWo4Zy
bDyCf+pLwVQoRMlEMrCC8CmenTt5QZaRjsegdeRSfwi9bXT2T3zQHRFK84JXaHg/46rJB+/3b8Li
ybl9g4fDmxuskge4ALc3ta7Q+zXI82u1uuM/X3pbETaFLuf57ArieVeIfvlSE1S9chk8R/4+fW3S
aZnIsBxk3B6uiHgWwkSYqJ0qH80G/FOTWiEoput4KZasSkBq4UFK9gn4nPT5N0flGkaoNYjy6bYs
2RXLjqzrsO8idyuR809W0VrDFZt7OkqTHom/8IBy+oafeLjYvf9JouXJAGFAYlfxGJSIgDV0APfM
LCSCmbeN7zwu8s62t1JlIiXAkPBVm3yzRS0pHOlpO7hd/jQM4w9nNHQDHaY5rn5c88asmQEYQPNw
/89KHIeL7Q65LVc7Xusyhe5VHsBVG6ArktpNGOBaIC7yncDoWR72WtCdLkw6hBV2/xMwS2R2qivj
BnuNFNKwUCcCDhd3yfPqDLC7xb5q2fjQIMjbjehcBzN197vh6jhRq2r/FvxmuMIGUpHegCWXfPhm
RevS9qWhGA1FZc3hBJktJRN4H8OWpXlz/ZU1J1r3jFLvsITu1/DmQu9ku8gNEZ6CqY1L2NcDsg8T
N5WkAO2s2xTo/HjfaZRUQvh5Pk3HCLNQSx7JEXFcM/vPCE3tVnTWq7TQwOeHJe2gnjNkQ5rGt7fd
gBNnDMH/M8kkGP5bDYqE+BrmBzL+lXo89ah9uJDc3GfGOIJSY89RXDy1n+vFC8E9HnFeYC7ox2e4
dqbaR5QHNzLjhjDsUKqojiobrdLZHa75GGkHAr8DA4lZRB1KDB8L47jBwkhcybttj38xrUt9MI65
jJ+FhYlDgCH24gYKxgE61Fvg0iX161WS0j7OWygRcq/TE7Jeer2IkoPv9dcnXh4+o7mrI4ijXhA8
rT8rplY88i4wijvGldvsSQgYRBOm3LBDvivW8uDWFTc/PpuAcn9cEHxc2DIE+IGNX3OILW6OJW3B
6AwcZJ1HzBIrS8lD7B0FKXhCElQjqwE4X5+cmIVE3nkf4U3htHeEQ55LCbvz9ftW0lhvOfDeLXYh
pMurYOJMt/wLt7hy55sBQl87iYuH04V2jgl9/tsngt5cp8p1BdAUbZtCA/bzC9ugrpx7tukFlXDv
KkQWrYCfN65mxUEgHD/nsKMBkFylRSUCOFTcDHAkCrS2dd37UES9pC8lNE+Sgif2UoGmMS47GXxZ
83xJztvJi70R7oIPvze3tBKPif6bmMbHBKwiopAj0gpsCeBxd2ezvhLRR9sm42FrUemZlpa44LBm
4vWctP/OY64ZrVe3l6VVoKmWuUT3DJhdtXkiMviGrMOrj7QQFF2O4/WV0kPs1dZnZ0kNdbl/GiAn
7lEDzahbONQnQkAGhnmitj0pjupfj68zQDNxy7PkzUznQdVJ3vnczUrj0xCXBIPX+xrghb2cUYtA
/B5cupdaaZAYBWxAiqtO7/k0Nkho7ybSwqWMTkXsxJBmte8YUzMAtOxVbd0MbAGkj37DGzkrPGkP
y4yrjBD4MrdwWqk9EDx6u3J8NircXwHUlfoKFYDz1CQmDdUf5P4DYhGS6k3dfof4TwE67dl/ONvM
5dPIdqXVHTDRSbLxr+RtllvP4eXJX1Wynea7zK4IQF5cGMR2m0cUiC6K0Jmtv1cguqmFNGttWC2/
Og4FKoh6G1P2KgYoZ5RY/b5YHFkcMD+iRZ94sCJXfcnw9fjZrHmjZUvYDxJfjC/cC1tLOT6cZjod
xOtRkRXV3zZqoo/QwXHMqaEalQPZxHr4casQdmMYyCr4TAg/DYBCYXuz+wx//1RDs6L1eAkAAbzP
QnKt40Z/j32m0rCs57Cs047qUWF763+rSBtzfMCzmxexgw4wwDpCuNn+K4UUqVKA1f8OHEqUIKBa
EoVD/GrmReejrXC4oajQRtc8rA4+AJ7D5IeUUKi4rPx5rkVB178FIhKcbqVhIO1o6tkoG1IdaR3B
Jq9IOO3zTyyu3gNZ1Jab5gbEhJ0Po7NNr5hjTT+tQHt3cjTSJgwVlPqwHagh3uaqbgzeQCRZmeuR
kgKSiLIgqigjueQcAVKK5dEpA2RmZQz/ZCwdlTYCHD7v2i+B9RLXRYiLMQZpAvxs0W/xcsIA4dEM
3wiAWGhDMq1J0AY4ltAuaxlnjJKir3EP03Ap1ImzK+ISLDgzPNvf0okiazKiOxQ+LoSff4D6tO8+
TFTcuM1BHKSDYjLIUcuscxzgtoJQpM4Qi/XF1eD2P46fL7Dn9+czo3rxiP4k4rRbu59UWWFXfVlB
1p8VRkBHRHe5e8HOXnpfKSUYfUkW94DH+Ih71OfBvfwwGCJzwzWF+VGxdGnOeufkmoyRimSrW0E6
PO2FE9A2lVRtSIcfFC5t11XxaddJunbmkvG+mRGqBhmVwmNV/zJ5CjkGPTte5zsz9v6ab3yXwSpz
Gr/rElZeT+lT7yuEheEFajVirx5rIeczTlChpIhC+NN4fQQe6gY5j/pL3g3BHUC4FMrKhH32zgBK
49mYsABjwoKT6TIm4IKn2bDk4obYOXUcl9Jj1/yPMvfmShdUF2+DG9vKEWr0tE4b2ZATakvGJ/dK
H689T1+IfONZ/jUuR2b+zPwaekgjv/fid4PGZDVAam6WMplRtfNPNgc3wpdOiiBp59XDVZAJRkA4
slPqWXe+TE7/jh1QSg2tgyJlAj9cfhiRVf4s3LTnTG/1ltanTOqz2i0ijYt8JW4SPIIVB0GGIkp/
/4R4KX80YPYHcaJMOZNL4LyAl7+tszLRuKWVPg5G9jVZjPo/CRImXWRJs98SSkiXCDYiewW7kMyc
WX93zeApwpq2f0yQzNMsnZ5Hr5NaoV3tXBzeFicbfNQLR0V4tqhiYymxeDKl0Tj/EKPgv9QZ/SYf
KN3ydITogImPXLvww/+YfJQC7ICRzgYNtr3y59YA79s5p+47Cfv9s5Ltg1MBrMvhT78pwm1MsfGD
AdjZVDUAicWoFcqlfoZdeZQw/KFmb9f2DgkvFKJJ8kSsNlwLmGv4awKVKHxN4reKqEkkemzPTJSb
bTjQfN/wYCxJ2P7sYalXwaszuGF0LhXK2ITjWS4FVWbtT/5OOXp2ZKs9uTBtuhtI5tV144uRyFqs
DtqC2pnyAGs+Y8eu6vFlDvD/m50jEzb6o/xkHnk6Hg1haND191eEkmjsNlPizBa+GTupjc61CYju
1unj9eu8VLiYcL21ZJXFhuBdU5dCejOXImZSdocs+tnhWwvajeSjKju6iPQnB6MQQ2lRtTuYUTmp
EBEFOYl8vwIjFltHl2Nw1dBdn4dI/sZS01BMozOP+clXHvLBGUV9r2CQNzanp6aub3fZu8/yNI7F
wiXdmyEGXKxl3CNGIBvQ3yMgJBBSfl8wNTjVi+K2PLq0uORTYOtRmgRt8FEXYE0fq3/85DKV5c0W
UCUIq65V3a8+B01iGpn3V20RfObezmY4/YpMuiyMsKeT7IOToHSzOpavho53ZpLJlurRiPvcXCgH
2n0frkEPiPFbRHZ9UaHd0PecO2i9VMvQdvnp8aZoosh13/iZ/QSKdjZIknzfHRI8h5tY4R3PhlOb
qZ3x/jtBh826LggkQfMYCR5qh92kXx8fXNjV2cS4fMGhayLZtpLkQ9nws4I1KONwzzwGxXSCfaFZ
8ZC4x9h9WvHvwaWOSB0NiJ0tVCc/VubRTJ03bKJa7G/A1yqtMGK/DOS18pFQRD7/bUXFEk6VfEUG
IFx4V76Fg8F+sIz2ixOqxSpB/CpTkLcizCZRvQEIcwQ2vV869NAKk/VkjWdvlzt3mnOCdtxnaIts
fsB/ZbHchsyUOiVEGdCuScB5qg7StdGqteu5+x2ZfvUCNgUKdi4i0Ibi3l14IL1Pt8SoEfGaEs3x
eIRAn/wXln7UIv5ZdnHE3d/othjDait3WKGGeLE3WKsFQHoLWF0w/m+o098hzfCwBXDZRH2XHpkt
Qsc/iJISP1hcCFl+JH8yvW7WwdA09i6kkrzW3T7ZvYMrDJ8JfRHL6jwS0u/GqEac4T2bwI6zVzvG
GPxmLGq6QokXul0x1FZpfKAzcIwyvGzXwA0eUxb1hyxpg91cfVl8YlGLY4EkJmvviG30QNGUMSuR
lypD5xyvAHWYTy8vn/l2Lgg/XpkY/Ldbh3q5/yEuUAHRoOI5IkoUh84hrTI60nsc3FinDjmFaOuZ
5E+nFTYO0g7r43aklZLQ0dHbEYlLpUfjQhSxr5I8Fgo2xonKpCiNpGTC2UjnjmOWp3nolbP8GJbJ
aAkvNPRgtUpadCd4PoQz+6kp8fNHcjj146SMHsR6wPyRWVBGcS5OhxwBaUvpWjxJ+natZ5M9Bptj
m2+PLQfTMKgnYwCvJCAZco0A0LAeevWLn5+pL/6Jg/G5D0psoym7RCQmAZVphtLIKIXs/sNNHpoy
PUTW7k66szsTVjfeJe0M9bcSu7+4Jg5pcOj307mykwxFB/LpSNg/k9V7y5jrEtz10D7sO6IAgBUO
jZ4e4A+IgAOSyQbZ9uSJxoahf3phh/ST7KEfEkFdIfkCr3wbuLEMcJ/Xsj4fmlCyAuxRep28su5G
pfpwFPhSgzM/E3BlUmaIRvEUcasktrAQemuf3+qu5PTH/XiTAZOIXNQBsJ6wrx6Moe6jMB33RijB
58KEzwXoVVTOPqtJJ3TXo7SnLJv2Pzc538clg95YfnICNOZiXXRY5FOZWqDuc3NUVJRib8h7+Vnz
iJMUq5ABlrJM/xHIcnUpDrz5S3qYhG2g9dx0qRTEdVEA51NxRgmaoqdW1bq1zLlikeDrevZbTfd1
JdjYwq9LH2Cf2nJlxATTxQu48gv8fT4VDT0077/C0qAz5jNp4vvCfuQwj8AxgBiaiEL7mcv/zSI+
2Gp8ZQwS4qFJh5uSYyzlF+BXgep0figp/WnxgT4JHeP7g54FVTYu5vgxpexN4fzr8AMfaXnrDMy2
tlqhp0+5lOIzQPr0pipYtdTnD9k1Gxf9evSPs1FrelS79shbaLNciUsyTMEMH6ZETKRXEctPHTHL
iaNfhzH8IkjWzGnegD9MDFhFFA0G5eEvgD2MEV6AN9CR45Keppsplb/5PPWhXypYGaxPzAsbvaEO
c5ETOvYJIWs7ZZMVdGSxrK2F6yfsu9qaWa1EMd5xgfLLcifvw1LT6OJUYwjfTDeQrMvkaRAKvvSC
w2lCRyRQpvYnTpeKGw6asfxMail8u6fi30BNnS5xabpupR/P5RXlmVXkt4d1aV6W1kbdyca9+iLN
N1rpRrjul/ZrGT3ogMP+K06FslXom3PsqSGLghl+1mcPH0eOcJdytbxR2aIrfocshc2hnQQkLC5t
pHvsYaLxvaY5wphYVGIQMQTRpme98a7W4boufRwFs9mEG4PxQr3/fc0oa7tyDB5gPu8tKgLp19pb
X9kOC+m/rWHAEXNgwEZCgO/4uWCyVSVTSEE3MHlyoHojidmNV/6cSiJzBib0PTv4yQn4G+IHYaRx
KAuJSKKTWwHxxVm6eAM/YD5Y24WI45YLGsjD98RZsiNEdS5WrIIvhAxYo1QnwnrvCGhCk1sqs67/
zS6n3rYnsnrh2QK48v71nTE/c1x3/LZvwoUzIeQ37PPewvWhktbaDSgh2fWHQfcZPvmA2fzBRXWf
+j0BTkB97mG3U1UeCCTtMDs2as9/EZr6ErB6mijzRFLLOajkWFsNEWzXKEudgFOB8xv1lbR4uVSO
MMWBisqPBAtgkuY218n4sIfAssBz95P1P8BXOARakARmUAW3/Q6msMPOw4cMwpQJj3x+f4KFX4vX
HwiCFe8md+47kJV6xyGmrbM/nj4ljME84eSkmEpLE6Y/Z5qE9ByPcmoCOu6SENevHGppiL4h0OND
YUQBSMhzwvcMmNblHi1MBw2AOSDUf9Pd7vuuG4Mu8Ti90KRuvlpamOpt4lGdRl/TAQ77dIuo5W5b
l7Lb7ARiqVtxs2HEMnk5qXH7z1qZ4zNJMqXMhGtoEoWCkCYXCrBBK0nDKn5ZjZH44RG52a9JK4q3
p9DF2xXlhEV+KoazUkIwEFTF1YUSSzpswKszm2inJgO3JuZRJm1q+yCJxHC0Y6YHrG8Nh8mfWkg5
Qx51lmvPFUqWid5xVb4bkbHfgmoiHqHG5py7i/X70Q1wsG1/XDd5UC/5fDh8BqJIu0CKrvH6fXjg
xkSllTDRLGJnFURINbtfeHGJS7LFBGkwPTf/PaCqqyYg22OnKTZf31xfigrOdpeC1NJhmWfZn9KK
hQ0YNeeqaUFITbdWbcFu+BBEsJd9NKpNRZEC4r3ogS96OypzWMWcfOO9WPCbnsf6bbZ+pwDuhtcd
Vu9Sqc30DPUBmsuqxUyCK66YJyhXrGSAnXdekOQ6i4IpaEPAn7g5HFwCBFgHDKuFfx+bKlhyL9BW
EDLRv00JcEqQILBnCnjtVh1Jce9W/11pp49TY5z9AYJhH9FeTzZrKt1o1+Lynpla6/HREkZtwKzN
2hySixdLVx/zRgb92cBbRx6UiIjP39sgBj4M5NOTDSUJt1GC50fVKzvJFSQzcGw3ZMCBNT7uuEhg
e0BVZm2DYv7mNKPO7ysZmWuXE+O62vXhUsEnnyHY2aMQYG57BqGeyvvuGwl2cQGNzP5EaRx+X7CW
IoSoAPx2Sf+P0ZZEnIalgS3SeSPZYpxxcol6/eaXezwnp5wD9Dl8HGvBwdLiES2KCz/kON+UTEUM
SUSv38u9PqzUWkSveXMNmN0bV6z1+KsL/+ldsYE3grZpKz+/f7gm5ZNUd33QHjX5i17TAmE2Efw2
Bwsh++9MjbjXhudMTtCpBV4Bc0Ak88JG8o4Y6aKeps1i5Mii+zzqQe1iIC3JacSSxEvjGpB6TIXK
X5vMHf/iGzdf7RPZqPXZcivCqhxcRHS4uLvtojTFfruRcyeqO/h6MfRc1Ci49r37ZdLzKW1yeJ9B
uv7887IHS8eECdMFQ4FQ2vtw35z0LfGxaL+gcub4B1R/FjB0rhNSz920iCGiERxcTZi0oMvS+Q97
ntM7yfjGCu5lE7PiQge2OKk8tuc5vYqO9mZqt0Cnd1nkcyhrmua5QYkjDP1jVtQEarTEuer7RDR1
fTR3CaXnuuN1QngDUp2d0XByi+af38ye2SKWuwf5sIFL9LDPj3MlrtfyEARcXUy0lWY2riZUMmDU
cm4nfu81hqX14kidYfC4t4H+0vO/hL3dccoC/qanx5p/Ezbp6QRQUQ02L+oMfl4tMmPrWA0jSRkz
kCAie3wEc2KZPG5w0Og39ARaFHp5bJkfW/9r4EdgYSuJxZMCdhjMDCpFRvijgtZ5SGRQ81xSLrKc
TzDGc+wPwtz2JGz7upJaoIlriEV5bVfmlnIbKS/mbLJRZecjRiWT129v6BRB32Fz9aO5M0EkkGgE
wI6VnybtZgMAr1dBenO6V9r4PbmdCpATX5xonfx5mjqTQ8cw1purZ3KF8oLzHBRkwIrw1o7KFOJ0
2DuSoXv3ed+UA38fw/gAFYkA+TZj3lH6vO5MkK+ah8BVaM6/zct+gXTBjxqAtomoQOoaYi0v5mb5
/xD41zj1fcRqR41NQVuzeXp9WclPL8Z8xzmWCJkenl/oqK976IF/f9K+wF6BcegAt1PFR5JO6+0V
I/+PNFuSFnX7q04Q4OkXMkKlTO5IvgNjg8lIfBeKjPFi1IbGy7TeGFVj35pMZ4qFSpJTljbBKO8v
Iy9UoYTAV03QOnLgikwEtbrhOtFPLKR0QJzxOe0JCRDmUyiPWmO8O7DRz3b8pY/apT56ZEBvlU9k
N95bMm5QiDWQtFPRhKz5Ue2oVPkrjxDTfT/4wB/PCRQxM/ZQK0m/UbEd+kR92w3MSV0wlIelAyYF
aDyjxY661CPLAJh+XpgAqFXACUlquqdeLEKdDQOM8+eMIrYOXrxaHlGgjQuyTFT2lYMlk7zZFmH0
xw0yLaDPOIxwfJBF4jlJl8hEmPGwHzKzyzm1Vs4vOhs7UVzOCEkknwWL71hzKoyjCaerJ/1NkeEx
ZDOtxZJWw3a2zqSLH1IpiqgIz1rEm8ROm86uY82TebzIlEnZiYka4ccCWWgDjJHDQp0bVROKqAqk
Nj4lDWuiP4okWB+prqynp0aCUT7MBE+DDlZIL0XwcmMmozyNmHEBSkl5o0V4Lc26AhgEsRenZFfY
BfF01D9HCs2Gd2Rpt9RXgXDBQ90jcxzEPiVCt0eaSs+7Mx195j4lPw1t9hJhzjC7KmGaivGe+Xnd
g/oqqzX1rp0kV+QVgCwO15yMjuKl3D2qgIbsHsaRfm7Qq8TkJZ7JOdlcsMWNOlmtV0qzTszNTwnS
GxRvAhDr4EbfYZ8pNzdrSDvvUBuw+nMzVhgvRcwye4BoglRVLiuxWHA/aKRdx237MtSS+EExvvdG
M1dTDZO4DLOtVt3sFHi0ZHX97WiY6a7Iyml2bojur+RvkLwRW6OOUPtFH5DOIfCKJFgK0YH15W0o
AVxM/Qh5ErsQPcK7CsN7vnFi4ek2ym5jPHJv4i2woR+q/eAFWY+9UAgJLLWt/EdVa/e24A2d8F6d
DuqUOIVqyZxP00nUUaakranVLIFgpN0qB6qJtY1eGZG+ZPxtOg7Zs9W3k/J8eL34vAn1DZ4GACeW
3p1izmirSBwHKInGM1OXkmBTsgyPjFNdZfhuSvTA3aRJ1AVlIgggGqgpQkHGemzgrbXS/ummlYCH
fkVjyaDnrgNgso+zAxnD/IOr+zKoVQH2ALGINldmB58Bczw/axq1bmf30lFcBKJwBtz8Ug/L64p9
mbi0G/E7zo7dGbSYC4G7A7kJUe75nTRAlhbjuLXCehmv11LOvfm3EiBs9rBBzsx2ZPgqW8sMpj1+
PbWSrW0V6LxqT5UPbiJDV+mtKpRBlInvoSDIPXy29c8lGfGXFJI12VX5oQ16O6hNxFEsTQwB/M2r
7XTLL7RJmvbt1IQkdElqDMHPnD+6gMBbAH1I+Roskc/I3R7YKg4fTaG45Ksa0IjXqJwV3Jqc9lJw
dl2YIsDl97Ih4732SEPwSzCcqGJk0Od05EacfJhiujZooDbIBxC+M1H1uqlqLeTQ34i8ichU1I6+
q10xhfENrTWMEO6CUW//QU9Dcpx7Prvy/8C4jerldus/LPFx8hE8QJ9YH8ROsOVceM0xIRgjc+eo
hQmM6GGoH3RBpdZRkBKpK0ZfNDhVjIE7UW3CYByhUPVMECjcUye9JrkJRUt9uIuQonK/HLHsY2/K
U+io4Ur/HPpsaR3jmuAvUTcyQoAanx8XnaYjFNk3Mrbnvv58OVgnQX6yhsqO4ZeSjNFadmQmB0eK
8W8I0+13wV6lrmQMPA8oaGsW20Y7A/uNd/GyDlnLOD8jQR+tBP6NEBfzJt+gy1kV6JsNYGkirR4z
lzLBzKqC7uCxartLCxlowFA9a3mLNKhNkexzh9GxZtRdePYrRvUJ/6XgwIh+l0uWbxCxI1KWYqrS
NPagBVxyq7sPW62o0zx4PFNDLqyWZDen5gt5Lk4FuZY1fFOJ4WlrWQjFV42eqw6qNXIyvznmefiC
4J/1mBc0xwW2IJ4Iqrae8Q6h/CszdHqKtY6NmWkD4SaSX9ELM1U5x56s5vufECwlOgMWG+bbfWyr
hlqbVKhtGyJcL7ddBoYQ+JS5umtMiSECDjFpBBZtzRiY2ZUkEuKPprhExwNbTAcWkRcnJwrSAyvt
V1FZA/+KPMJdB2MXrxkGf/2mKuHUoFxwCby9LJRjozuc/Z7uZ3Tti9m6vH0ORiu/bCmCGdEykun1
a2VIYO91+FWoJx6nMVimVcEDW7ai6PQr/WPM5pcL8b1fCmBqjATtDMseLHzL7ydiVFLcTqWGWxVP
OoRI2l0WIa3z8U1Pt2mmwsOI9C0/7ThDesM/jPElbB38CGRZOxj/UgZyuqIWoUWMvdnyb+Zf+g3E
knhXlxwUT//47opoc+Ap+kaJlB/+zBaRjE57v3vzINkKqRiylqALO+f88GyEqNoEPKTi53hjvu//
I3mt6YoV4oYIW5mEnKmr1usfKLIIt3yPKMjNNzM6w8FxKWcLA8mjWQ5TXE8/gXmbKptJqlQJkEyQ
FnBiV/JnhaROitKDQrKGBZB/80lfDy7Qhm77CAJs6DtgvNaE8NagM+R6NtxW8ui5lPDPudVlnIR0
T95LQEyRwgzBdOED+5Xy/C/s//h8BqIpVogoUAMsvjnw1Rnon3uioNVzsguO+Z6ytBxshwTQzGEz
vUCRMrrj/ASYOKNW37L0uppFw2N3Zz6jcqJ33YVD3YsumGljNWjJ612GYzhLwgAmNa1lIe4gFGyr
CdFhp9QyiQ6k+Z58Mz3LEVIE4XredXTQ1tkIjb+iUT2moso8rpdAWOLc0tVxYTz+dPmTM44Z4pOQ
PpP29MXVdwV/EHnPv7jzVFVKb0irGWZWzABrUAGgdrQElAudeqFjYPjOZ4s5nsmY7TSIY7UxOLhU
6apPEKXcyPQ0yMs+WcaJvey8sZylDohhB6rKHpLi3fF3LSyHkUrvoWFafcDHv9KkUjYr9uY/1lBh
M1cgDsQj22N/dpTiAdeuSXBGHzs/0flnFdz7vw/czaTHju9vL4dOVVNof6qO9laLW8ralhzvlo3w
TcaT4Gz+Tz+SN094NGlEGHfRgi0hmdW0HJCs8TX++riGGF1SkKG/4R7f9VYzw5xfWC9E3hN3KP7m
ypTwSElsgM38dttDXnZvUnWGZSFRnZM08CGh5U+wzJqFJeybTjyR1gFMLt8hkbvmQ3m4sxG1Pt7/
pytzOpBOOzCUtDPhdGGOtquqo21B6TBCWszQRWcYFurEPOR+b2b5orXnAi28ncnkmnPgXb669PGF
TulmN9yvda1mxhKstbkNe4qs+FWbgcj//Jc0AQs0ZnmM53uPL0Gkv+jfKGG1OsBnW8NdmeiaXUWi
DKrgrC2u1qBnOZm1nCOM+4+/02NXeidHR6CkJV1SzVM1Lc+zsD3IYv8VZeXLJ6Vvey1amp2EJqZe
XCf9JObQ/Ucw8PO5KzUKlr2sJujQcMTvxWA0qxLSu1TiGSQy2szEQK+VZQrl7nusM9AuwaK/qGfu
ss10KUuGnS7DzFwQcR0mt9I1SSePLJW+KxfmWDd+cgU4d+Jq5XMSeVjUi9E17L2SGsPxJproVg8g
DxPPhDHyW5wNupE1ftM1SXyrUFJtAeNMBUWP4x0lhSjXR9Br/1HrnqkAXeZ4GhBBB4bh8di0aIn3
KxXKRO17HOT+egJuFqEoLo3qZesUH6gyWXfCbjw84Gsp6n/Uf18gomTfVcHXQFeDY3q3crJZefDd
vbs5GPcLZLWtMzbOSFujGeqRQF/wjExvSOmOv/76bKioOQ4UFSWVdnRKl5m9W1Em2iRgXfFUnTLZ
5OnJZVvBKeIdFRbSt8QB+pzWBBaxXbDomUYIEyp/FCrxQuIF6k4hp/k4l0HkWjdbXQJeDATVQdbj
QiPgZey0pLWsFUzUx565cJNxd+N624ZjVdYzbA5ZAh7sg0UfFH14fpNR1RMv0Nj3VY9qhcJpBTMD
9pXlysicjrQz3+6jYHKSYucv6pc9uyJyfSs679LrdCXfpMrinKOWHhehF+IF1T6kQYjrDzTNg527
BHbbvMcXjbEU3T9xHIpsLFbl5304bBOt0O6EkMSoLad1jB/nFDIfw6Tot2LO9xJwkDRB/Ovd1kJY
E2emnUA+2F7ARDbQNnHcWS2yQ0flBG10E23YWoUy5blOJ/ArGGo8oxmU53BkAPv8nLa2g9tQM9WM
68bJzUiiIWro3UlQ88vRDlPBDCqQ4tdH1T53E2dTg2S1j7utZKuN5aN4T051WN1+EViQnL+znXKE
1GqiL4rkrzCmRcAzmpRgsIGjKPRhIzIJwvwFsOVbJw0iV8SIoqpp5Hwta9JHRGnFmQz7L3zGF7dJ
PNaWm44Bl9jP3R70vB5E/iy2fuRGb7YaFfEHxmEIuLAigsUPLbkppTpRHmVj3niwRfyHA6AxfK98
OSo3mdsAXkyeEtfGdCZS8QB1NsmLsWCb3Iyb23Nrk/E28B9tHWeKpIqMNbH+GbA7sftMbvoiENER
maCgo9sGrphAxGshlLuucajxP6OWgUpcDiljEnFL7txcjM0OVkl9UMFVpFhxKQ23Cs3/Ghj+b3B/
4K8PlIm+NFSiQoscFxYWRDeOHIB8R21geot4jt46b2J3aBoR70jGwWSmJ9v24KdR695H5kf0LsUG
jqQ0weGGbHXaFj7hSoj8V3h6YdiVQaPuFAizb8JtIuQ21gbW510iUXvqpRXFFXUv0Zba79yD0ve9
Q/4exwjev+fBMvJ1XCbEEc1u+fD2ffnnb16jzBf9O3n9EjxoQjNPDKMKHCsmWBxYQ/VX1DcaE43K
xN8z7Gmm4Hr+xxBY+7bsX5wi6sYQAB3yKVws6hPC+3QHrhoMt4aD+2gWlbs0DKAmbU5l5W/bv8l3
AAZlgtSAi1L+0AGLqMixZ6gnA4nVf59WVQESAXbpuqpaiBnloJLVRTRjELzhnRj44uWo6fWXHPVA
3c+mX2V0hNHvFpDkl5txK1yVy3A+FhyBKE46hg1qXkjIGglPIBu8qHhbuTuqV9JWH9tDiAzy8Aa7
KAoS0y9tWhkZkufZ4FgIIe7pPp/I96IvMBp9rljkOZiq1+ltpHOs8rkCYbDAg0ftl8vDxJ7fJin5
RV2bXGVSqTDqkXCx6UeKpWE+miS6vov/24LfJ4fBekAL+T60VL8vUjRZiDf2EvyHFaDuu0bkaWcF
ULB6639vMhtamMHbQYiJUHB+FBBMP4gO3MYb6lKM3v3qGrUr/pAdBSgbKUe7WDgZQ+nUiljuvPH8
/L55bsbNeUkaIHYgV0VcHVnxgLgnCJMQ1joqXTU1OmnJWSmVtGbgZoBEikNElY2llpBG7ldoGzA+
ijSQaIH0geJHmWGlOdUVhrHjhkgygb07wZHlDnoomzxJnqwA8wtu20gRoMR7FAS7XqUe//4xQmAi
qf1Uf/nXd+qgsx7BjPHK90ug/PhsG9iqBnMvF/ksEOYK3iNPrYrMsaOw1C/6uJoGE2MtuK4R4qI3
ZxuFrbwT9HbCpTIstRmvp6K3juRgWraLpGfv3XflNYafpXohj4lTC87CWkSYpkCnY3YluppEdIxU
SEyhWC44LzO/cbMrW4Qk2Q3BYOyZEw1CovJqmfdLUJJY780pur9zctIG7Cw9m4Z+Yh/KA/6lf2nJ
1ndYRaukua5MUphdoVBhVFjxZtFbhbHNfdD0mx6L4VvcPp/CR+v2Gn6JOdSVzoC7ladwLEIXA/ck
IgQyB/2TyxaeU4w7DUcjRPtwvbZJ0WAAVxr4q8hLDAFTittsJf4TGX0rNd878LlKegkAwxSSkC8r
QOXxld2+44Tn65x5OqMrME87IM9hHuhICx7iC4Tsvbuqu1Y+AmYREhQW+PiAqr/gGdYI60Iwk74Y
RLQHJZvmZq0QVEGqAVVvJiCEVBEyDWg+9ktaO3uZch4TKWI5JD/xSKbpT/Br+LD9sq93j5QroZyE
wD2KjqMjYod7+gZ2wipbUQTqoEegkOlKJRC01egPzGOctNUz+qKTYFfFMTlBpngLyOQ/t3sXwpu7
X0tDnG0yCVV+vrkZmNDrgwMTaeqxcTE/0vQVj7EuRg7h7bJetPB7NMkvHYEEZ0C6Xfw81r/cNUCX
WE7N03oYr1JsY693MZXpvu5IoeaiVNjMoJKwwHo9Sro39NC5Hb2121DDW/qhE/LyC7o7bLrCiClD
T+u+fcCBTXrkX+Bd8WSXh7d7r45zXneIFN4vcAkaBHJlff+9OXgdSCsjwSFTGQXs+yySPGWzxJQr
kq7D82wGOA71Jd+D53l9hj1uGeI+ozV+mXW3X7J2x2g0rLgU70EP2dwYkO+AoYPJXYkHp4ZKHnqm
3MtlkDYhrPZ1NsiVchwrwtlYd6JX3me3wXzcXS+whmskEUF7hHkXaqhRmajVNS0P+wBWgHsMPQ7s
cZSX1HhQ8C0XAkbfs+NGcr573JG1tIMqttDf9ZoAcnaKS1OB/+xD+qx3HrAthRtGQEhu9aCwHbmf
E6un5O9AAnRaJbTUh2pM0oLcgKBplHuLUAmrPA+RzX5gBmhN1cedqB7mQrjaY1dIyQPWJkSbjSsh
GbXb7gi3spQzhEjDo1Kk/iqJRkzmrGuoYiTEWMPag3bKkx4n5RwX8ggjc9M+8QI/DND1V30sxNSu
YtjkpD3IgAbYYlkb4L/xZBQHVSBjwSl/GZCuS2h+4m+2vEkKxnbu9KV8YssOeAFndXeXU4LsnFBv
V+MT25FcJP4cI9slpFOUiO9uhSHjKZWSboV2+5N9i308U2YGK2s9BUfXgwqSsaF2x2uRErwKmETc
cFvAAUneZj+O6t04MB//URodYkGgWuxYaBbK73U78z7sWbasQAyCTeLuH/it0kMh3ufxjc+tPItx
HnstvLq5lkNyAhKZ22iLzr8zOgf+FY/ldfi5tfbmokpppdV/xf8W6/utu66XsXP3ZnF8hlCVAL/j
QTO4eJaKlhEOO7qMUDLZeQrFjQBXJ3KWxOr2hEGGOTxRGYsgecfnB9oTC080vvVjL1MkC2PsyFWh
oVYKoj2RUhUkwmzQDiCol1FmeC/AG2DCmSTVt4wAzo7tODM28biJIDF52DMgi6fA2eFiSH9us0gi
/CskNk4WMKrQ8wP7i8v2JBgoIpvf5+g0a/8iDVZyj8ExOOsnrnQJqQ0/U8ZpW7983FBDowfzfQ9N
GujSDjO7zohiwK35qiNAUycPVhxuEIcYz0XkZfyKU5xdt1os4QFXyh3KMcYZMcUBgb48TasS7yJB
7QW2TftyVo4MVHnTzB5A+7jW/PeNUdx2ig2d5HPfGcaZAGwIsb0a/C+pqWw1K+iMSI0qQAW8NV14
05Wsh9upWqFhfEWkcZ1oXepf/CZ60G+rHGiq6+JfOIWlcfiKBg2FE6N5bgYqyAlFG/PMP0GUaoo0
Kk5KtlWSiQEFmWyHuNoKc/z76G03zYOuB6jTs+5/5+d7dvZRbvbRSxZ170uj9GrgjdSP6ddeVCgQ
a9Ve3Dwcx6UzffLiGp9SEweI2MkgttOkeucAYiCogN9iL/gL3cUGFe+2PtIXyZz0wywfeVjnEisN
Ye66I5e8FAVCu0nL5wpLanaS3WirjBBii7Hh+VhZO1A9Ll5+M9cdJtSc6WqOJ9iPN7OaBT9ttXxU
mWUbcEl07QJqS7jkMYL7d5iUzaFhWxm0OdFV9OeeIMwBWLEhs9tTnNW0YvQPzIvBLfPh4u4/rYs5
1iRnPZaS1hOL6KNxiX8vK0pOxvual4Bar+uptn0ssEBJwlJ0Hsu8ROw0AdrVKu57EqQuvdb6HjZn
d1WolRx7PijxVvCCRxU8QiOkB9yQcQ9e68AihXr2vtvtkc6icVO97RlNMXNqz/8bi+NyUoLEk5M8
agp5AOd0C8Ri8rr66wxjbWzuU1hxeNidVOgTabYwSXBoSRfrk74VemyWbLEdugYA/kFBrlFs1c1G
Z2CO8pNWG4Rx7qWjRvWwUTfwxBVupuzqFIT2suyE0+D81RoG2M2wR3x8pfMwBKdc4hzKQ5i5q5ry
c4CoZJXQB2BAi5BG14VKBqKQugHU/bb5yTmI/ti080hkcjxcqJJBRvCmeWzTVS+E5IeAppPQsY3R
1pRj8+81KSmv5SbbC5/5FF59QggSfvCt1cytbjga70EVb5bCbZKqRhBDsLfmLh4fiLSQznBiT2Ju
zK7q4Y/8ksa/V1RIpdZ183RYDmAGMTTmWYb8BrFWGArsdCWd2k2/5OcjVvMb27IFkHg62YIvUuAC
Kpnb4AueolydOgnXdScnQiV5txTbE+UWVMUKs6k+oIo7+a7leWJHQqdydgqqYYp7k4Ub2R44OtDd
CsE+8JMYKzqaw5/Nwv+8KMNENC64lMWfac8fQVl+9S2a9u+AebxfRQRyf8NEa1QoPq2m69cHDd0/
KPNKH+8xdlQwhQVy9x5quULz9UPXC2bSUdw9tZJ868pMc3q8qdekbUTRrQjZ5KXETjNc7PuDcaFB
Ez7zQl5yVw9tw4aJH1V6auajltSNji4bhTnEYbOOrvQnhfrJpfmWyuYueBG7KjghQbQnkzroWCt7
JGDWAZRNiSW/Ty6nC4ua/7YSo5Hd+1HrO2tFrPK9zGO1QTc+ecwIMvg9Zvd8zddl1z9tWBugWoPn
ZIPevqRZXDan9kmSmidUe3I471Rjk3Ztxf1wqLsm5Wf1yDuCWIYGTRecdk/M1W3TdHP4UAvWIZFp
ToehU7/54w8v4+5Xorr+/TGUz31XYShSA2hiAKgNwWc1n+9aoXdjuM21VbYqeWAnDV1+nRnu8puz
4xIu61f7MG/tvNYpDYCr63DvMKG6DDPyU4yXU+9j7xQtxnfCgnBwWRUCibpk8plVrpvyzRcHbaWK
yHqLrvfH3duhci0/LM8pGhyyzT6x9pB5O9VvVCm4TIRYehii6ecp7BfAY96k0DTjMGYXzlr7TD5f
xrzNGzo7QgdpOs28SPaQfuOALvDpRttDCkXwV/8NMLFiWuwtuOyRpQvXR7LYoVyTgHTpMupZYL9V
uYOElsapZlQ4DxBJ1EJmMVQlN0GR3oHzp8caZ2t169VulLYg1F+nLlu6nSrmFxxcHQS4oMDHNSx3
yFBP3PD8YeQPmdMHkp/rLgOOk7029YA3wOZ0avBKXNi9U3t2OS0cfZVJXpoLpjRP1dMnXq6NUgex
Hja4lxINFcAT5BDv2HldFfnNXOEXM8Ue79bSaK+fdxhRnBwBGpuRKcz7NStPIoU3mxyDMfox0y2+
9XQ3U7KPVgVqEHKfda+eEIIcHnD4GnpvlHebAUwy0dBH+EgeBAh+wH0Ca4o50uB8B2SxQ53oMiJJ
ue5f6Rziu7G2VVS6eltzlcxa1HIOPDZscVOO+WzEhoPP0VSqBbpQoP1d28lNSAhTSMQliwyvaDpj
J6bY1jIuW3yRHmyge3AGkjWgh+hvjT+mgLVTrhP7SdaNIJznJkeQcJRfzL0W3a9mLpbl4p4Fwroa
N6DWy9MIk5irLMaxnHQUe3mvyUg2ioBG5i81rP681Q8s5/Q2FauQ9DV/izC8DH1QGh0TkCdFfSdx
92vAWDIi184pijtyJFUpSPncVozPdmLynoQFwr4b229jtJyKmWTfxHHLQbJf/zkT7i4qnSDQdySl
+e5ekJGNY0vEjlFVToSaiMeEx7W7cpIAHFW652FBP+DZ2dau041YRFjqsP3cam/pM0KwS+7YqTT8
+AkwZVExQkuRAIvdPzFrBeR5LU3AQbLHO2QKcagIYsDWuub5jfgG4QjlHn6mylYeWaei2PJUuEiE
BU1rcKutcT7TJIbmjtBxwOLfKv178rTL29gK1cS+Znpz0PsKR3S0bhMywoshTwDlc58x2BXSiIiY
ze95sWY0MZng3c1kZyXjVwvPg2vKGxALYmD2AaEus+1nTeq0e5ewVhJQpV6bHtMNhHgRUwOels+O
mLgGDRxJqC0FsKQb5s1XRot+wafLZDjWrW/0aSYy3St4rzz3olQmPRlUSVghAjMUmUsM4gIGxq2z
61CCgoBbjtacdrCSLOdSZKwcKO0znJtXdHb33NetMn+UVw7ahBHguBAGjEUeDQmWoCSOuD5CE6ey
wrc6cX53SKNJCDO+6eD/QgeL4em1oPg6Xubk0A79PMaCOaC0+q2O91nax/Z4lkM6sKMgvfqv6Mqh
F2ybBIsI6JlCvHsBWdxrNM434r/iXqAp/FqEUyRcg/E8h0HYW+S/vah8gT/ZnmYqe1WWuhSwtjMm
CxlwfBCdX4R8UN6JHBZ7KBoz8WX6/+3h+kn/6OO2hDYjx6e0Uykw78hmCWdRDJT7L2zRW0a4VDc6
SHaz7HB8iIBpwwtPPMBcDcIpkBoQr0h535K34TTp9VAPazkB8A3hUjaNh92R2Ozt7l2Fo/xsj6TR
eFDPa0LiCLngeU6VvW7h9OIaRuXFCG7211cAXKIzNsFvh1CcDfAzHLKE9NMyjcpK/EEofEXM1NFO
DeLQYRmZfsTckvCtuv3m1503INfFoB6c1vyu8f0Rwn5L1tvDm8mQFDdV5TZcvIXhYEo58lF8akzb
0jb3x20Saa4GADwZL2JbqiCOall9GzYHKyrwQFwC8zhQnONFqDDbTLHZfL7dRtOdzmpzvYOVOcYv
HRLVk/vQv+jrXPyZPfwrllL3JvM39uW4N2fzpQzsiU+SfpM0o90eVT6WxuJ5pqfjglN+Cw29Jicp
oPKJv6VK64xfn6rwcxllL+0rEMWVS5CWKmkBZR3ypkiKb3iVoxuQB3He1BqvrSRvXkyv4EzDS6Y1
t2wirPfQpygGv1m63oyBErQoilTYfW1nSVv5kksdMYavKGFGT8VaaUqeXX/nLR+At9ntjZVCnmUw
dZvjmoAGHxj7OWjmbxXCnBB0SkcJ/iHzXTqnOecPMWcDmfNAlaXkhOTkcN8dwfAvW/WS3jt6cR3i
sicX5EJaGuF55tWn8GHEwguPW7rIrb7iY2jXIu2bS1YROWAdwx2PKW3KLzibYgMR+/NFNdsYdr7h
EMA8uQ8k0PIwZ/8WER79gKWhvAkNMCkwJDB4nFhqUDCldKl94XyYYH0aIo+S+ywFM0MnyCYSHHJr
EgtmJpqMVYGZ0VYMNFjQmsqhDhDeoO4fLFlM/A6AzptlIALHP+IjXUNlb5dbNhxyzVGRKTnWNO25
9ILtIiB4yumwzU6SrKU2R7K/Wo/Wxut+TqPqdYqA4oDv9yYARtmv3IBuaoEze2R7audx/rL0OXCG
xN8ZnyJq8q66AZayJ5ykDwSuUXl/7tQJAust2rai/q0OR7sfGTcLSWnca3Mf413Y1z25RiY84+XL
5N6+A6wzvY5UZ77w49HuHeMOjLF4iWIMAMsVJahVm33PmM9aLLeLuPzYYF1xwfarmam62rWlnqBt
naM0SRNr1nX3SoRNnBW+P7bBIcSzCC+qQjrIPcQGZ5kGBQ+4YQdJGcO377F5M5U9e8KHti12nlq7
VMazjT31Q/nd/T5Febfd6b2QCtjFE3TWsAFBFmKvx06YjGYVMWQpTpg/VMeYQVpg2vKVMWx+igaU
qJdzUPPesEYnVPyHTrxk/JSBxNtb95gFlO5xCc71QA93IF3TgahRvQqv9iu3p6f+2weWZGjRwLUS
zTHJH5lQKkg9IbwXiT9EUCBrUmrJVVWeAXMXIv5Sr4vSQ38SZIjb44h4kZE6XxomoqJBwl4MyUQx
A6U8NZyI8dnhL3yUP5plAweXT4TH3OdGLA2EOS+uEK2HsWpG4/qqsdWa2yJlGXl5G7SBkxjb1+CC
OG2f/XIztvbRu4kFe786TiPfo6I7VgdVy6E73B0+PztKBGfg0L+M4Le9qUSoZgQ6klj6Ou70aKcO
vb6vjGvp7cId/WjyCvsbF+cuQHsmLz1nQlhkdFywRKleEhrZ2n1xR3ELTS03/CL9gX6h/8dENy2x
yrZHdv6khB7kZB94sMNrBrghkutIV7vHuaaroFKkkDCzVm7p/I2UQWkXuxEg8t29sLOjulR7tqLS
3FYX3iTrSJ29ya/PvqsYZ7cocaGRPwugbcPtoBF3uLZihKTGxpDrNTzsjQMffoU6TGkJP3mJQ9M6
t+wrunrqOvU5Ox21fgH1BHPwVZcvdERl59YrliO6hm5nOcwejbhDokKvA5PThtYsy+jyOFngXtoe
gw+wPFOUORV43tszlxIpeEDPj37Rf+abU8lToC2EnB5k8tOl6EbXHb2nrgIUAFlfck6tQVb75B4D
VSkJ8mdp29vwHmn6ZVc3O4sW01lE/7dimYVSOWJV31lcbmhUD2VjuGRwEIdfncUApCE1jHL+1Up4
uVwSk/enP3dkFuKLolrcYt2KpmeMKEr2uISRBL6BNwQNz/FBYNZawWwy6h0KHJe2ZLLeINzoH0yo
63ipoNpNLzU9hyktvTKTniP9Kbwc4SLeUjHaceDDcvSPrOTCWpncQtomnOstkgbUUceMDqbnV1Fs
SyIIS4YuAPng/f7Px1te7UgLptt+AeCY3dFyNvp7fxrLVDrTVTM9NxwTzHuvkWM5ZYu/wHLUjMJ6
0KlbLRyaeLFZv2goMFcPVTfeGjiwJGz+LRxXBc2wQE1VRWmTb9gk6zRxc//UCFoyqg/8GpFdupAe
0XcBwt/t5x7GAacfgCmWOp+jJnu4bheIAdmTYmPWWYQJoKBSkdnjlVuy2mwSxAcG3ZUTFoK/Wgc+
2v/TfiuOxV948LDh2SYGws8UBKPqHLqnW0jJOqsuRzqA6U7lwqU1WkvxoqRU8SX3TLTRPGlVFUJC
3XmwS5eBrvp+bzePHJ617hULmqv1T99/SNlQ1Y+ZW06nkxml7AtMm35HMifoF+7NeHfc8ImD1RkL
sjh4la0FX8WSIEIzH6U1NkizbE9mTcDYI2x1v9SM3RUmU5hW/NgZZXgqiW94s//2DrcwpuGLYwSe
pHRnpr/tTIkX52JTAnIIEr4qk9IgJ9XdRXkwk87BHwpb9cTH4bE0S8qvg+30EX4LDQ5VDU70oKL+
dqjUALh4mO2xXBrk7VnExDlSmFlq0bRYF7sKEWhib8GSLwEVpsIJ0COvtE5n1JMVtKmIf84JuhQi
OZpo7+fabmcUaD1Pv6vaOTRw+G6UY4kjNqbbqPeyJwpwyqg/ciuzbtJt7GrILK7QEPb4Oe25+8o0
8JJfbB5UZk2yi+bCwzXV1Mx81VTA5FfOZheBCnMRuzep51akYy6JgflOvYONxkTMjnAP6IvpHniD
omhKFXYuXbSDg6Jn695CJtF4fsq1cvNPtVrSOuuKkfkZf2dtAioCi5jMs/EPGYoo0NPkjCdvjXN6
29gV5M9HeH5kLGBUEIqdWX05Ck2GwXIa8HqxUFO36bdHL3fauYeVYDpxzQ27z+7b1dOpAeVIJnM8
NYyVV3nyA6k3c/wmcb5MvkJ278IewFEuJUyYSWgTymRz3KkZh3Dnj6WU9l8C0tsSk0513qh83cgT
XNPdrMG3PvUzC246n/ICwff34MiIMHrndPsfa9zJQSaQZZixYGlLMsFSHSwRI4ER2nSPLnBbGk+0
TyJgGyDIDIrvkgGUqA3axibv473wEKLWOt8iql/uFhy80XstOl3r62xIoaRJzgsSSm6F9BYb9+nx
NkMWYEBjfVj0yWN307Fzj6V7GYUQK3tUobTiHwMSwRpvN/FW3WaXKtErRtpH2VF7p0JbHbadkcHh
S8CyPqBQm0WCUSg97WlYpVXhib6JVX2nxCSxIulD5XydpUlhlrPaZKWwPczSnRV1UgczMXKMJyyR
WZx4bmMGUv28zHk1qROjBTbZT/B4+0NUzj51eHrib9f8v2MhHqg+BVR+nYCDAj9ePiIqpqLvaVHq
9mWHlHNcR8UBA8dF3ZaU/0JbbPn2t1+SwX/hXbM3uBHLHGbo3BiI71a+Q0Ccy1wuxQSvOZ99T3HE
VuTR43IxFjGO/7zCS1V1YgeHJ9ZWiWnOJvWCsEKbpS9p00BLZt5He4bUlb4UDtol/MkCwWyv6B38
YY6gQUwcGU5axwCCIIC3nyZhiGh8M06J7tXkB8GATQDrq4La4fypOmzkhyC9j+GWaedOxMXRBsrK
GVAnz2EeAtqaNiO2yvz2+xBOAcJvacNyrsfjfmu1sks7hBXnJbkE+Q0L5J9v9Bmxy4cxb1QWOSMV
Wr9V9AhAXjdQIBfJ8KqPbQvVu6DMKc4bdLuFRlHZ7JTuEVvdwuqhsd6XauCMAu63F4BobVU49yXO
OlWF9OZ1AOD1VYBWdO2IQfqBfB7PlnAasgQuTvqmfUNK54wVlQv1BufUtK6sOEXwD/1VMmgzCYc/
Qzn43xwidLiWWQVlw7AStTNq7X9fISS7vQeQzCzpoIeRdkkOd9oATE5g4a3rQte/hXLgKpfThpVV
0sO8rqQ605lMh5r2ugXE8eFTuCEkB5OjTq+PxRsGCDtS5H0pcWLWZcML9xCN6DbDHZfPwCOrG2Cx
gczbXYa1US3BOiu1L8DuUYyUSqldPce0krRC9m8qyCGOdb+kNWVVh0kIQKGXalw1R/w0d6R+FR+J
DybhxlUBR5oajo/+Tj/bZlc98BUAB1qYWsaBRZQ6K1YFf6fpgAiTOCVG0Qvgn0s7GU0CZdPAZgS/
1VtjblYeM6vkByxsFAJ/LBgmLkMvk5adLQ7YgDP6HY6wNjXy+r7kbLc+612XkR6aHtCNSGB27RMw
4jsXezXCmbmE+O99eQvfjPNYVEn4S4apOSXbqm2PrNVV1DkOCkQwIzzcRKPTeH6wrgVWPHvoW3I2
xqsP3F4O6GBxFz/c1r/qd0r6s5Ux32n+o0u1iYPji80c4Kd+YJoKyEJkq0xFwQpX9WC7WST2k0IS
Z9qJuxN+OZZcZK6vvh+kacUWk9Gv/ai+ZHlZ/y0ElZF7NUIgJBPFJBVIAJd5qcotbDEKSq4eQ+N9
EoYEmRppoM/12/EeM3dfdberRGmlt56wrj3eyMlrQ6JbXqWlIHSfKdvR9RCHzwuvMvVjxVX3MRUB
TMO3JYC3UqAI4CSvs2iN3SUt84RNunGCyUxbUzg3Mz08ukl3exzu/N2um38VOZ4N9oqpEY4RBjQ/
RlcfMsv8kJysRVu832gC18c4A0L80XYvCgT/Az6PL0WGTvdHSD5ZDv1Xl0BqqhKPlxpqLc8Wq+V5
xgDyMZcGubbcg/x+yXf7+JMQtCyUMz+VJR9CIOHVro0aN9t4hrS/r2V74LoAt2MBBSQWXSAs7/Q+
CYzXSRrx4AWSet1KMzeM4Eu1qAKFRv+cKFPmCXaOmtYsiV9cpfnHa7afP5072kTKpC5ZT7RO7eau
KxpTRT4bYLP2xLJ11IEetEZnH7LZXyIvDtodaVzR17t0xuGt4dgNjdXkscDo8Y0io0sg82evcvwz
+g0m/0zvFktaJqdjhB932rnqJvrKPaP/n5nConxrf0s2VUBUZYOsTx8IWs+kHUpz0qIcmhYF5X9r
4ghA74d0tOJdIqcpkkUgwaF4MDDdQ1X9FJehSx/JUFkFk/U1OQMg5xVa42rZMsgatKGX0KNytbva
u12Vj8vZ4RDDBRifECg8MlKZJkbqMaNN4mx6UT9O8aLYPr4JuCVTYNASQC70bGTs6MsTUSi7mJ2l
6vJs7cCuuHftYFAymwaQqiSR4p0E20U4SKGKSwvMAbwl6CajqQUXWfsVe/RFv9ygMzbE66bFZwQE
N1IVSOQGk38GlAcP78hYj8b5iXmmIhFZjI/YdsIteaY2cHhxbnBE+C32Q3kHzVefIP2VR9t7KF+d
fR95biaOytmVh0EgdScXvuV5xdSsh/8IFwYYHOauzyYXx4PTzd19NZ2buih7QwT4AEjC1VoClllF
aVpDWb17ymtDq0JL6GpJKM1pFQN0LMrmDciWCv8jTaNnDD8UoHCgLCaoEtaZnsa1JfL45LsJBrcm
UG/Fia2CP3E4W4/rPM6JyXSXCpQuQixsBZLYm756wV/o87W/RPbeEKPtXdhNi7wcqeW1ULwR8qaF
4/yXuT8eENboEDVyYnKa3gauQ8tFSAs8ego6THYfK68kE0ckeVL6K6ijtSI3oC1dVNinsa+G1dXl
UJr8L3bR83ODE1RgnfJjVOqSZWIG5jmSDAHwClErQeS5e8LJdBJc44kMpX/KbN81zzB5pRUBNq1l
H84pT8IUskH+PU34ncrJ5P8JFPdXNKpDO+1TdNZJWEzlqYo8k03LUQnu2yqheZWoOKK2g5yYIL1T
NS1HX6nTMtlEO/+gUwaUoUj4GyFmgOMsSlVe5ovPLQGGnivNcrdWZo9U6W/KGkCnWYdlKPDDlHXi
qrIwA2tmvsda6Km1RJ+tckFJHuGbmkA984VoXjI0AQmTNj5bGYn3MQAnbu3I9rlU06F9sN6iN205
jWFw6pZZg621TvYAnjX4ViNOR47Jz0+LMb7jdemRx6E5B15Vnh3GMVy9Qobjo8GNskjelHJgdhbR
6Con8nAp0xRC4GbF4/+ovaKc9PLeC/szJzfJorXHpU/p4kWkb4oggUC3ThHcK4iEsPMUovv8CGUp
1C5sZPlP0QwUz/UyIMnTHpSEQwxvtZcj4IW3NYCmPIdGEv9mva3/cooF4QnTkeUeq/7KlkYi2SKT
0ziFbDOykfob/IYafoDeCETi6L/xUcTNY+f9giYm56LIe2nirrAI7TpEt0K52nM9SU/km9wfM3sy
jWQ5g9z471a7IB0NFiejDEZcN26WXbSnFE0jjX6Q03ur1AdJGNjeno2hdkhtsED00IRb0iQstH7L
omJXyBH+K+5MhLBPpHqIttxk8YmIUFtI9pD9tztqIfc+GuaRgsmJbfsdQIB2pVQi+8EE5I394H11
j6tU30KyCaJI9CK3VM0LSOiSKpgEaNxw9qv8Z0i+SteBcnOxXYEuxaeHJBk0sZI0eLUR402ui9vk
uJwgm8cGRRx/dnNuvFH5bCypn+jcO+ZDAFvD5y2kZbLkrQLLBVR7Co5gNmZQB3YWvj5H7jsW/Inb
0+fKKWjeOTlLRNdHnzvirVWXA71pRB8Ss0eAtGqkWBVENIS5fnEnRGGx1F5Z991BNmvCsE6wBfRg
FnusWVY83giaRCl70z+nJM+sgJioqBMoTMAKxCHp+6suaiYez8uNVlrkbGf8HJZQb/TBDfbti/4d
5q9KIv35bnRCpdr70wqJeLbzU61Nb9ybag323xkdmTHzgag9HXOKn0KdkB1SnwkeHBr9b0PxAY2g
H4dmJCnX8ieOXfxzp/8ONHdPdnVZQDOLSFXtxTk5GInL92Jtbd6/8jyj6V1HdDlsL2C4pUsmlMDM
wHJuIh1gQQD4xpQoYVhZt4svq3Nf9EcNigAzKyU38WiEh7v8rz1AhvP0FyfODqbbI+++W42S8Pb7
0NGF/Vd4gkKIoPY8p/V037DzpbGr0Zh9fmaYNOOphsnUi1rwEf3EObCrz5aEL5hX5C5YfsjvV5kN
71FYwbLUHZX4pDowJmhuhA9ejCYjJ45OFjyvy0mfKYwPHDJnRZ0dTSvg7tgGFJOTAyk1HqtJA3Ka
1eX8GqI1K5dkXMcA02oCoBMgxnJ99om1fzM8V584i1A7pE7uLE9AdX1nUuZrrn2KRbalCsx7DQZm
l5UwmwORHlSvYBe4U3/xpOxNn7wwsz9EN/Sk26Os1vok6rIY2vnAxyYpsAzAW9xx/oL00AovR+Vz
1BEAN8svbiuskOXTE/857bfN0t6AXb2Y3qzgCxFdXjw1Msbale7dYt9HlT/m7y6JemFpM2avkTXo
R4rx+wUu5Ht/Xy1tT7MaYUhW2GBQAkwiMFMvdUF+5kQs+7RoVSbXNRndfdv9nRB4vJ8xlZK+95ZT
FYRbcPtaKGUMpojlfVlhdJaPJ3/j1Bfcx585GCfda0WE7mJ96IXwHjgLVV1ngH8iwExD2lt38yRo
GO0zzffPjVAZS92Di8xFDRq/wO1UDKVJskgvzBS7aKTKJ8asxtfdrtSwoc31+cuob5eliwyS7a3s
l7yO14z9CchvqLkO/JfX0OX1BJMGQ0VXxBOJ3w+S/4sqx7WW7MRtJN8kSfPWavizbruZeej7H9TT
0YJHP3fWFvDDzVpXcrNpxXfaa3PrwqcPN3JQckV51ywrUiIYKBy8Ge4fAAO6g6mITPnFaVnT5huY
xmnXXyHB+7ftwZHwxj02toczveoWZDR0ntiHbrKkyflBpNy/1ZRykGCDXwCPa4rKLblIM2UIaMR5
i6H3ZUQaawTJrPsP3jq2JiRUPuwWketWASySHzMsfUlQ0VptpqePyBx1wp+jKDDwkRpsGVShB2sX
kP2tmEWCUD32PiYoLVbtHpRcBbjr4tIiF9OepEMhA/4319+8UwgFI0iqGd/PB7lS/UHDdnQU60R5
eIP9My+C9ex8kXu7/mFNw//NTeycMmKnTZCyUab82C57bspZh+kYDRGLM7NwN85neR/w/gK7Wrtk
WmwyhWURRCikou8N9J9nTR2sFqi5dNDwKm/3+FZBOA0SVxHPjuhkcX7ybTEaGDmVVsYbeywylIH3
Zrx8STSGhG+BXHkJcdmlxBAFRcoDZex6MGSlcOOv1W7Dx2N+EcUNZX+T9SjYpxLA6atrYptQeDhv
8EYRmrx9tJX+MTmcnUHA5nXG7GV/t60dqD1T1D4s6sq58vtfZYvVW8VNPcryo/c+vK9bIT7QyxaD
tw5W//zwnCblJcy1Q0XYTjmiXc+r/nk9qtRvWFKP5GPASp+v/Yz8CC38so70LpEFGgfhlJrO0MVi
v9JyOyn61TN17miPazmL3lcYtrxk9N0YATp9nGoiG9YWL+6hfTAiLOZhnzVpgVy5ZMdwpLSobRAf
y6sFuy/g7ZzmdkFBRGyt5P7QG54pLrmKCq+Nz7cXljlBKEYS+2DjHYLnrXIlmpzaQzdB2sckbdqY
YikuCJJ60xPdxjBKvLgKWkNXnIolBflF4/O/CTt8FAxnZibSw2In0qB8J1xSneqkTqf5pup6F2mM
M/0Hpv50UjXZ6zi1tsRDIV9VMuW3TZXO5aQaBfkS8PTPdVLHhPIpged+lYAF28gNL9kaoU1QfRzz
yJACCXvzbDmqQNW/iDcOpIDxZ78jhtZRULzFzfBp7l7RxnwBMyVYc0mAF3l5KesW2Pv5oCLWDqbm
UdsM2JBqY4zh+gt3LmFWG/rrpL2TPQJVNcGOJh613vMbWy46R289dZG3i+rooilfb7Yr7xiscVXj
+U9GKsLaDgIOK7xK7BJrtfeo0d2AT1mbP6tF9/Z7l+KsJ/4HU2MfNEwqbGqnHvsvs3slNn3R4uzB
2u2BlJUvDUz6+HcwnonfUZL4eLMH5k6hzxD9pINGausNlNqect7KQW2nZS113OSDCFwKXZwVrklm
FkoyH/pEfbZnUOTd6cvXw41PeuRFWX64V5RJ8xaCzxQq1kQj4MwRZjNlc7wkDETXjfYE8az3HtDE
BCAt4E1pHYRbmxP1Dfwu8znZQR8NPJHWyecSX8Q3VrvCcg6mc/PVRgWIwnXUV/KruqTpOchDpwXm
5FHhz5BD6ke3alFdJNu93Zz1m8tXP0AsQ0eBH171ZtW+7h7LsyJiGcR5AneioVHJLUbjWbaIz7K2
A0PiJbNjCQcAF9+SV0Ixs9TJHOYFp9nvLM5WpsPfwFz/AxJaPMCeAgdG7ezSigWTtDi0e6OXeCbd
BUi3mVnBRK8CfXk3oF5zmWXdWVEnxavQRfrKnEbj+0HFVYDx32hlduCyeOR24uej/GQsWBS3pIvN
7F1nwgT1yskc02innJWVNYJXi+X9rfwY2B5moGi021NskWZa9UF0h8QNWLdCsblZ7CpMkpfmYs2g
XmsFv3jMdstcCo9GTrLKFOdUD9TBLULSZgkzOt7tkQC3qClVArh9FwnhHaJTgX9iWnUSb6uhrh9T
OQjFlzdiewbXmylCly9mUx0J57reBt45foWheWq3Eby/hbqv/xeYofp4tbgEmTvz24epYfyXmCzd
xm4mGr2owZ+q3MboBqhCyLbNQboSfP5y0UKjth/seponFJEN/5aME6rwePstzSrcKks2pEc2HrXQ
Gb3+3rlKKD3BbFChTtPPdf49mRm2UBgwrrvoM/SWyumFkZiSjqmAKgElEJkg7MujD9MlQKiQh6Q6
fWDoXzLO4ACglMqIGHNRkn8cC4uGYgnR4BokDQ5QS0ChTmB/9fQbUj7DaQWbgqQTNHRr/OiqTGOO
L2Z/McXtJh/PuGrFMZmh0/SpsCXU7LzUhKdR72ty8B8QSfdrxpMZhqmDQ2Q3ycvQiUoJhdXbd7XA
VHhKFuKm8iuTbkjZMe2wSuqNhcrv4/w0WLY0Jmdi+grCefqPx/vDGgKsCKBX88pQK7n4Fc93wRIl
n96F3sps+TbWcIC1g6GJZGZAkSQ3ZNZXBMw6qkQASNEPgXCF/2ZfGWWiMJHJdzrGU73jX4V9uOTv
SbCYw3L2nZPsfoIqRrEGs5EBPNQSjhbESp64w9xNusQNQQLqz5PnbT9EMYhEMO8u+r5Wk69thgN7
TYpAjqB9slK/O7g8FiHFhQrEMx1/X6yYDp35WV3RaCBHA9ut/HN+6lu5j4TXIby/X2kl9FLvE70t
+xNI0TDFBLUGEUf9NoFfI2sICcNAtD8J2RMsvVSjih+GaiSb89cOiOVLqrGhPtvEYazEaKd+LdgH
tHNqU9agSGTT25+9FIOiNsjAVsylznFwFq+BRY7HEn5oreGPZPzl7Qlyi47wlg+D3n/L1kcvL42F
8v6nG++Azxfi8DxRRIWXEcWbFRlGurqjeKyclwppe4Y854Ae7EvOgzJdf+guxvfVitycVYY5PvVu
DcxCzFm+4QsGFVkJKm7g5ov8ijo/CWHCX3GKCzr4umUns5AKn+pS8DxbYlTpcczwOa22iNv5HHVg
kCXw4s7VNjRbDVS7X6uW7IvMUS22XeJA2ap3/WBq9A7XUJeZVDjy1J+HhKyeUH91Ujbo3HBRe3pD
noxaBRugpUu1rDBt/j3tlZr++qnhulLl1NMEpHsM++9jjdJn8aATXr5OVldVsnCtWRcYMnHLYiSD
rhHmRQKCPEL0XKw5/qDqN469YGanq5scjy5CKy6uJSlgnxZKwFv790OOcFdEgf4baES4jeNavn94
jPsYzvTr/Wj5809xfDAfOZczMvwhbP0fh82BrEJxGrPoXdSsdtVAUJ8Vt14xwnVE9B+ASMDxMYTM
Omi+qhupU7zpVd/d+ljjWGiQ9rU1bWS8cz9vymIIl/oBv1F/LzgXBNb0LFc/abkuiKVXfykvT9da
/Ma7AZdI/O+MIU26XbnHIUZQYaMXPVk5xhYeDU5AGE/nrQ/vV7eeZJK7xX9ewGWWjki74Cz1SL/6
gL/BBRx/QPI2WbrcMzc1VuhuwYZRB8jOJZom0bouWO0BPH5gbfFyxB13VYs1rxSFLyBR+ooNnMAG
eIyG9ghoe7A7Ntal+UdM5c97erqcuHAVzYVRVMDI0Rn7sVKKu9wyQIYMnjGthhpj56URUcX2hAWe
uGL1bvPWPSdqreEERBzSbGN5LVZsfjaQ3feH6/ijkwXUNUs0uGCEpHx5IFmPiBUC6MzIrVZ6TwZC
JIaWPCxU1wJswQFPvaJg6ZsFfqcCX3xbl4b5P2NAWeJRIBZfdGX74vZWLnADQZDzKQBoXMk6X+HZ
vbEUuFpuSzfcpP/LBD0NXJehNGCUo/iItcFJ2lQJh8jNhrX4cHivVrzjN3u6eRTtLR7RBDTYfzuC
cTB8QQKOWqaUNwtJFppGPjMfrpA4uPht2DGD7hhL1nsPPIHwHvewAsBdpNrUinipTTLbGZXiHn2m
zE+DqAZY6i1DJCJO32jGoQDl7E7uWEdkBP3Q9+b52GEpIlrkRTCcMWV9TMut+LvOFRJDhy/Dkeqn
bdvtE9vq1ovOGDzH/MbYG4zU4/i+BvvIpWVfcRgAu1H4BYfIcth8TvjWFa0AsI7Z0acPmuZjyDnn
nMFygoeu1RX4ex7djGDsI9yjTl2Zek8xIWS1ssL3JW0p3QEt4Q/3n+aQokIjae+1Bcl3oG4HZSQz
RhmvZB8ItDaKvf+RImpji6qUoUJ7t9bguZiY+CzR2JfWu+6NYCxiDrdEgrt/9jaL3LIu+CJNlVXu
SG6Px7wVkWRNkIJgcrieINxPmuh6DVy9rnGN+O+D5nF2gByzvQlY6IhJnr5fC0rpPq+azWms0PST
HMrjueVVGpnEc1yNcHi7EWvue71RQlIvRqXBT3lLB+MrhlNxEbWxsbtsff38nh3eybtzoLAjOEFz
6NEoWHCFvTun0w/qN9YfrHcG0TyjZ4EZqcwmLOsAGyqBLXH6m3PLqvXIrfq1iDO/KpDkgvIkIoAV
Q1V8iELazSpqAgBKHn2YV1B0Rjls0n5CxNaSAYT53TVgS0Q74jMz01fbjJEhsOGbxJVFPBXXdw+o
KY6u5nOkyRoaPBKViWEQSmjZJCGHxev19mjn7gtRUVGEDmGRe0Xwe7ffjq8QfIo4zPfzHBXSZnV1
LW9Ph8gJ/IBouyat93VEaxF5bsPjp0uMJbdBx7iCF3s6AAZNw8t2pHyV4fCbAImtsGVY/odTGZqK
SI1b967f61zjyCjef9a36ebqbBTDAE7JJQgV5JgZSGkWoGzV1ZHp3JJq9Ifz9MdPwDMIJDuXu3Pa
FGbaVGO40bObW0DQ50oopf+IO8A10QM7jcCM1naqhYgvZENKQUfBRqIJ/eZBwE9N7x1nZ8K3YT7f
2W2UPeR+QVWudJRkGV+GLsSNWt+vnksVbH9hE/8XcrQJWDS126BXCoo7b4Gy8a37DMWugdlzrCxr
NJH5p7lJLV90BI3NRd3bJXhXQ5bq1IMRcLQDIL/qUlkpUoG6qgljDJE+aeaDKSfTNHlP6z0jlMsY
339U/BABV0U6E+OJr+596Sh7Pkuhx/X/XHDuRfO7Beoxl94IlNjBd6NwNhAzrO7+ofaU+FYNb/un
Z4kSGVbqkRuqbt8/X2wAgYQEZOSm+abCb+seBKGWAfZMtkMIF2km3FnL3JbSaoGDMFNsu2zcRON2
LWeKNFyp2TsLZknjXPqePnGove4yvueecyvMCUpB4RBF0ljeivGa3JNU/1P/ltB4WWmOTqoVzl9B
XEPh60x8HARQBicWhm+sTYbpyjgg+G/l3LOgy+RbNC2P12nTCfe/Hgc7apfCZXpNxt9Poal12Enf
4mD9tjiaLVm5klXAx3SB8EveEKjM87NnioYnHVcwq3I8Qq3bQhGOXSdyA/9l7sMrRm0JRZyTH7EG
dwYPNGpy0uw7Gwb3BhLmAfBXbIaZl2c1E02kmAdG73UdrOd+f/KlMvuK+Hf3OIw7eJuQ7/giOx4E
fka4dc4I4Giao+VWckvSwW6lhqXfkFvk7M9SaPBAp9s3lo4F/gkg+L1Ci1uiP8p2IF72nILi1X79
XTlbfQP8ubf8Y9yDSqV7GXGddIvN2aasKOfuDyBdAdVr6TjKXPdFHdMsCGZhdJy+RFEMni1cfQ5h
+RS7L8OSFbMHS44QW55ReWD4VzOyPocCorLPypfifpePTzG6Q9qPA+zmYj2Pukwee0r7JTKfQqnk
jmizIxKI3cfZ1Mcnr9dP0Dprv7yeWb3m6y42eD7eP+NgVNXeOi05cRKo2TJ/2/+SMNq3TyvPK1n0
dWiZo4i2mPHqmdWNUzIyp/rYEWXK3faPeQPJylNj02mE/ozCTUCLosl/i9ZmoMyfgMDUukvkYkP6
Qy90UZJFBLX+qz6hOl6OmFFMLOoczomxGw9plpuvClhv9O0YWONdjlR26qqn7qMUbhxsEfU8DotJ
A46kpb4c1jW5rYAhWIWKaFOQtQBZE7VU387Q93ZxR2EAYim8WcSXzO6JPZR4rJGFlBBqS3dep4SW
jEzL+Es0O3dkPgjhS02YMAmMjFO4vwUBx+Euiq33Pp5y2RwuBEQI4GqrmioEkh+DODeoze/fQOQk
18JY/v/5S0OitZ0vySlKa01VwruuHA2C6IhVSHzch0y9yRKKmijjsp8JBolrz1eO8pS2pXmCUHhU
RowgrHllBvqkZJlYedLR29r+TfFjkQ/izm9WPNO81CdurFbYovo1coJmQ2iHVIk6fyd3V97Q5ooD
tRLMAX4uxcdEHOFjsA9ZxTXyzSG6tyRLz6sro0qf0sjOXd+k7wYj7/gwUCwY+AcxeqadBxgFDhDs
xXQzXBVHVJiDJ3U0vmq/9VHSrSjWkAO5RVPSA7BgAD51Kvr9w5Co1l/8J4oxQQQTShFL2ESNZra4
VySaN4FSAxaho14qLmhHNsz0sjbt0bHdKk6PRF0Lf6n2xgI3cAvfaOOkOZDqRoqHLGHfaeqodlRX
vCEUrMLt3SxUCcAF3sa2LS7xu9lPQHKuk1sfqjqcdcTEC7KSbz4jbpR3D248KdL6/rAW6E/5x/bF
HHqHFlndCd/n2Kq21bsHnMyqHyAIm8rpFNy1bGlZEBTmhDW6SmeDakZ62iTNTvK5ZcNM/zdH3QUo
6jy3Xl0z/aNMwPXiwsLWJW7rWvNxZgPNZsIJ7EFShMjc94c2KeF3vBCu4x56e1UBkY6899+++4Go
Ion9UkJVcxDdVtpJ9t3wlrTudcnvIaH3p33mkmwuB+fDhUaA5OusJ95Su98zqvv8TBoSJ9qNv4AN
tnLUBg15tZoVVOkyDyi2tYLOmt0R+7iLXvxigxlLxM7fM+Xfz4h2xwoPXyJTNLiKXq6BjErwsX0h
6ZdAidaT67XV6vASdfFtcVBEuEnQ+gRbZMfh5JexOp6bVVcmc1Sbh15EZXNj2vO806W+hlvNQb1f
QFsMbmKExoqLh4By1yGsxXoTnX2GMReCwMt/asvvIKhzKTP90ZpWal5qp22NTLTA2nL8PRYG2WcX
dY6AxipPZQsih33wHZLPRDbWCtJLj/QVMgnwCH7Ml0ANqLf7O4vJiGMxc8LesC0XbtIIUd+lCya/
+O7nB8FMBffk4YjTcWjN9HAiGbaUjRwKaa6wWA/oXtHwnJ/vX4vbpsAFtlgERYMSgwo1V3vKVbdM
4RcNOdez4wdX8II4uAEfzVKsBPqGhrm26aFUOWbWFUkkTfyfTzfiLFZXnCyW80+CDlR9eGNasxqS
N/vh3Y4ep55grEdt4cA6q2RFj+s3jLWwom9vmPYKJOENLC96LPuC3MNe1keq2FlibDy3DbLK3pnM
8n3VVWCkuXxvyzegkn7MXHcWL/dYQGDq7WcX7hXIMNrpw6lwc6kiNgb7cqTn04sQPgeerYTXOx5g
sy9x7LNdQS3EV6o+UNHH1rZ/89gWKm8nWVt1Fvq2HsuCkYU4JrDwdC9olXA0N/5ZemnsEW5a4dIy
DzLH1M9McOeRW5CN7NIOsOpKwu/AOOguKB8jXtRQ106z3MkEs3ncuBCBP+7P+vxUH8EZ+CAKiE5P
SUfwnEEUxm/tSyl0gtqvdKELklM3UoLbkA1abTEngi2lfkM6XTQHOMe7w0oA0MOGukvkln+ilmT9
GZLgk2N3t9h843QBcR3UZhH+7srFw8xxFW0JOxHS7pL3O0lat6ysY5PBg51r4g0btvcmQZ383I9e
vSJCthxYmBR0qCWnqPTHlgZJWv24CTBT2x4/CjPuSQyoUs6PDvfQxlihtTE+PjfXJ458d7AugZvI
3pldcihqcc3Z7pvlPaPD8GH4td8cInTp+1TWDWGEuMr79+8lE8rq9KJ7pVL+rmKow+5FPvrD/dHL
aWXAJjD/B4kcTX/FK9StjYMvfcU1ZiwMpG62llxRZY5kDeTjLdASVyb5ShxVrH9/N7j7RaJrlYln
QejiQen6bm6sEAezaBiPOTAh8Q2lS2z6nzxnGvzCf/tnjPYCjGc/huLrI+TuGLOT6Bgadjx9pmsB
vHS7URYCxaAuOVmhjtNjXN4JX9unTNfna+VueDdbw/hYxDqcfnV5yE7nPhYr6YaJuBKxdnF7j6xo
vWx7x8e70fO3DPPZZiaH0qE24e7t15ZVSXVzwH9Boi7HkMHfaaKDxOXUTFMtHf+MAnbXs132aQCe
dZRmjNLKwA1nqFJZZc8c4xVwJSI72l5IwItzea3gsLkX9apiPjGk9BVkn2ja7SDm90EQZDp2kuHk
1Fvi4cF/r10o3hcyxGkyuZZAMJfRyexQ/lDqv/YSiQDvpjXPnSgICalx7oiuRVXKfmf/VmXQRVnp
+XFscB0TseBuLSoMwFwn0DWN0Zr8XLsgtQKFtXzmNGPCD1wMZzWfAlTXPUKzt7NFs9Q7fotYfoiq
FZ/a+qTUvfRL2wrBhFNhe6iD0uJDs0h3Mmt/UrpYfj6T8U44kSoIcgGI0cILkexB0KYlmzKdF/mG
1rBV6jFifclE+5xlsMBeRJEjqU9EyCIwFSvs2ePGJbCBP9PZq25Wf790C1CGwO0wu2Bbbdncf2Td
tzAxSaQr3mK7KDWfUNtcFt0yilqlkePvv/3oaf1XY7Q+zIhTnhFz4UEq1MoXeT8kX2uTqqK5TJOY
jxWBpospLwpBndoCZuTFe7qCp9WnTb0WRMWGJyHKtvy+DNEHMOcoLZOcBr03EYs/5t02jfQlrkuV
4gl6InqZszd3kxXAVbJnEOi60FZDrOxaA6nHRVwlg2b8j8FbYTvhfTZr428np/0BIXqTl5jGLSxl
RXxEXB82+WuqD0D0GlTiitzpnchAgywRYRd6NNvlyh0tJnaLgsEdWFk/i6vJNZKZERKCYVVL0ptN
nuahRnuiyuxBuWRHq5IlyBMlj9NMhj1GFt2iH+jyPbhtoKrWDTQU/Yr8WRVoVj11q0J/2vI8evfq
dR6sctS0mGPgvDtemAnFo+kqJ2darTtjPM8cJ8x1IMotJZw5j6/d9G5iUP3tOrXrB0X2lFUt7Oe+
/DA85btsxgecCy5xx3Jbct4Sp3O8BCFbJEAwqmklpteElQNH9lHD4f3kDt+FwOjeUEG1X8rkBHhL
Qf3z9QZ1t0tYKQ+k21Ac7qKjg2CIUPMq4mkz3+AtOLlTF+/9eQqwvxdVfPYztVdDTQe96QfttX0R
v7YzXd6u+FQ7N7tFZfIoSElxpjnF1jw6BGP8mXv6br1MDc1RufN7oBU9YcmzMpIVTMuUaJn91FBO
ZzFMex9adIMl+Gwi1Ue/3uXWkiS451q/Ip+ZgL8jHXlpNQtOzUrg9xiN8V/yGcbpLJyzt8dftbVx
CKImTTtqYIjo7vpEg2mvn/+8uyKeUjoH9ARC23K6My8p/oM27TMqG9Y5+Oc7fOGzwEA8nu103CEh
YETEHKZ4Wcqg8cGnHaDnCqdLpUzHCSEbHaBVzaIgqAvLrABrBcy+oEor0CD7GPFJHYYp0SzUWME8
fFO9btq6CCaw4n9IbDi3kOSvsdKNuIdhaZiCakBb5K6FeQr8qb1vTIJ/fVoRw8aDZg9cDIF/TVO3
DSODaCOgKM6H4D6iAUTUuBJpSPpsmcejwX3O4gkQY7A4YJg2N3bbT0DKclB7HbxH2D9TwkZceBaI
dNuRO5kNGR6NVk/CpaxB54dmsbT9VhRDgqWP8172gvQgrRZhbw+fM3FcTdIVy3Ol6wp2x7N7+nEi
MVfTuABOpWC7RVX7PNnYpH4CQkxqXM98BGYBc/CarA0o4lsPBb7+S/7Xff0SyBT2k0MptsZABVaL
7d4NOUUfNWj6xstCXkAU1jqLoZxlfI79/nqw9fexmxpLK5pkSsVxDR4KUtItSJYrGX0buAPn7p85
8f2bJBztu0Ep8r+FMyT8viRWEkkY80u3xdftgs9N0ariXWzpHfwni5KfIlYraWlqmlgBQNuOIyLq
TSfYwjgyZVmBqLkQnU2/zvfu36QaqmHudWjPnDuzoPauh8C4XwE4dgi9Dhw4IssIdTzKouKBABSL
rMFoL02V9B9GpvRF+Ekso09ggNFJyWNc3GMYZnzfs1CcdTsnnD9nWtConDh1+0FmM/rEUjcqtXkR
mBDTAcx1RqYNTpJVtTJxw0l2XHB7mKBYwioJszaiSH1rxOeJ4ooZXKI8WcZCSvvbTmI7/EYMxTGe
S+OXhbMxwEpDJTtl2DIK02iocdu0a1N/2zeubK4Z8MtjPLdTPdzJBSBcSeUHAVgg0xxm282AicvU
qc0FCx3Xsbhx++5/aezYTsz4aN5sltQ6uup43jDTyzxTHmFEkKTmTWkjJFYB1N1nsxpiSAPv3MnE
4KZlxMDuE9gnY6LTXl1pCBiWoGcrgN5FEgodF+O8doNVk51Yi9dz86kOfbi9ZEhvUfL1UWfNj9ZT
cB/2321DBUmlu21y0BWiH3M+Bcd0ymcuvOJUsZRQKrTwsALWJuRUiR4/RU/8TWdL2ANRf8hVAnK/
Kv9n1aDwgaOkE0FZMMn/Exr1+0ptTBFNyuw6I+MkX564hg1L4N+7zOc6gOA0JVRTQ0HtGLoD/niF
iuZzyIGPM7EhKcdvX+fy/xJKfE5aa17vDRATc7p3dNSugZEpABPN3XVdb2/+Gon+HOjDBv2J1QQx
SiaE7xcGPHJQRmKYmni7RbsKoHv8NC96Tz3DPz7oM7Me5/+6QEaRVo+acHPlFWvXQ/IHSpjdrnV+
1uNcyU0sgLhAn1P7z9z6CefWytXsM/r5i9MKmYI3Tey9lMVBfcLdRxmFKhianNi2Hxxzh4kF8Aeb
PKyO/j1iSR3MdfkHC+Uhch1zJs7FL7RlrnexVHo0x5W4k71YQd6VZySnMPXcGTkuT/RUoJHF9BYz
9c7n+1S9+7+vHUsKWQNflVAXAIgn8dq6gYipCt+I/tA55kJamqhwSOfPhUlOA8GGAkxDb/6Qeh8p
QETrUu1RY//BWIH1+S3bYjdfjQVg56PCfpR6Onf5yBdMxW7/VsfKhFgjc815vboHE4N2xuSh/oS5
uVeXJQXJq7bI/No4tmC5QPWhUQ5exxLdaME6Re5wJxdeGH8bn4vDFwQwVg29SZk6Wyn6Gq5rgl06
Mpcc8Ct8Xo4CPO4o9EMamfnK45j9apzy46zXmtcxLbr45vsQEWuZss7VQDrX+YleHZKcNk5pNeUI
EcOAALt8ywwC2DyBGYcMGZUfoZGtEy5zROJvS05gKvdWDVTk5hZH+kp/lGISRvG4tXlwKF9cQr7a
H8f+Tm9e0X0d+6cTqhsarn6uArs0HcGim9qJwKurWWt7I5bMNl1ooSWmMQfbhnM0EkQA4AfK4GNz
XNTfWXTMJ2WPK6xHtML3Bt5ROCAPERlBVT6QTz/PHme04W+MbFL+SvPqdf1kAEFi9phNlBKIIiw/
URB1h3rtW/Biay/1g854GAQgaglJZClNFKovnnvUo4y5zakKIvoT4L7ceENUPNbbGt4oDi2kcfC/
+6uTvN5fJB/DE8deWk3oKAsVOlTCxv0/vD3a9BlifRUatDqXWA44+guC9O4/U/Mh2MA252b2c7rY
DMMYO9DwhShwsF2tJ67Ekg7OOtqr0rkJFgTDag04WoZU5XN3aDm7bTaIPvnLe3XSQK965eWhFci3
RGz4xUMElpDYpO4HVeAODU1q5dEW11Xn7+i+b2pqpJrOukpxoxa4THb5f3mkOkZ0ipOEsaL0WbP/
gP7a0wCJZIStu4FYdMqpBRg6VSuEvMjvirICnaHFuRuMO0Hf8Fn/KyexxabciuQ8p2SmAlrQLqgT
q6EChVdS8OgpXmDhOhvPjKKV+UHkn6/ZfHWNQ39R2Tm0WRhI3s/HW5KMa4qWTt1buuQg4whOJNxV
A4DPopWX6y+lc1pbG5UcI+8N7Ky50WOqeCFPylV8GqQlpsZKikh7BHXWhLqsPu/O8L/Akgxn9hS+
VBxslnuu16yoRCgwJUOx2TY2/H+V86NW1wxcjncXr7e0lnfs7mZPb2LQOoeJWDCJDsYmFIFLzBzp
K9d8TP0ey03Z1gQhPj0RUNwHBhpN0o1OYohBvttNo8lx0ly7QtxFIPtoxdUEScSKe6beDv/6TGi1
Hasa8kas4ijqxouTwLom9aqYVmXddk1IpvJ0j/FJrOjhpa/FUT/IOCdyv8/+W/xF0pr//hQQuVCe
3LUeFuLhiq3ZvqPrSakIGRpYxMHbVNcZjt8GZqy8Yqb2XntR6KCZDGUAzWZ4gbRvOHmI+mmVukkC
Cdfaf60fT2y9Iqs4ZF75lSqKn6K8/Ig/x1c37Thi/qMrt+xhMgHrnDe1CMzW1wv+KABBaQly08rH
DnKbzNbPQ/W+wZPbB1TMbrLVvWF5fG4fSJRQJw6obHJpyLQrK8vcnzabK2GfLq0becgosWl5Lo2E
QVhPqzIFF8xc12zCK/W1R9ws2aW00xuTRTomo/DsDSXst1lCNhhGcrlS0ZgO8qVuArb63MuLRIkZ
21MzpGn2npcjUhKUpO1lAtqAl6F+lxxdCEq+XenRH7dxgvSQIEWkG6huGA6984oT7riabsnktOXR
aFyJ41U0pamuTOA9gL0h1CRtEChwiCEqAzrjyMJ/SDRzRVaoN6cE0wDVlBH6ydc5AyIP9V6MJEum
2LRkzYlhlBvfNYENOvshmBS5V9JPhRXWu5iee5BK/sVtJbjJXdc9rZ6GZIo6IAOPlKbq8h04xgb4
AmbaXjDMdc53Nx1MYtpKMl4GtuehzBI+HVmXQa8qgPYZy30Npuiv/CwfbNGTiwKpvxRpeR78Q6Fi
yvVZS6HTKOHsEZJXELWXdRXCPijWxN5ZsuairQzIWRaWRor1V5f/zGyR3sZQiJEzQsIe/GgPwD8H
LieHmfCkswlEIN5Oe8NnHcRaz2As6VYyIOcrZXfTPwmd7/ABWzIUP9DPsopiKe0qyPk9gf4Fd1CZ
xoFORsgzDAJNqMdCvaZ+OUIQDfL0MYr4//29gjC/VGSsKYfMjCPdOf7anX3jkYcSEvclcY3WfKij
x3Tm3Zav9OSLbvAqm8nhAWSjf9flI5/fGC8t/kSc/bDB9lNQn2To49R8AxOYq21aXdwLuVGePwfu
HuSXuwNLOs466AmSU2pyuUt05JvPAeV6aPU6VQSSWl5xxOj/bYuM5kBkmCDNHDFIaw/Lr6VvakSC
eBWkImqjHDEeKwvhLzQJZyLR7KzvFJgu+s89dwayfSLVI9cWcKczVabLiR0nTUEwgxIbFMZksAf4
2iesKc+ylcVTTDxljVP6M9uWV/KAaAHAmTHxLv2IQ3WQK9a6+DdkE+X7IAEY4CDWZBc5aJtPuoqH
BwV80M8c/nuZUvGZGJH2HnXH9ohE+YslFenI4ma5MDDlr36MX8rF5Zj3TxXVQoPcA2DjyZgzv9f2
o3nIb+5Ysaw794xGeNCn+vt6OlJLrdTF7pdLBG/JFZVrXJ/qfTGoDk5dcVJ6NEYEEKbglLTBWuIV
gOEr313eez2JVH7iGbjMET4i9II0dgLLN7sH2dUT52Rquv4N6O7xHz5KbYGZWm4srciFxKMssudP
JeEIfjsJ1wVriMn6sWeCUB8gnJFwqF/1AbmgVUexdyUPKFXhuSaJvvWzPVndVfSN9JYhVmG0CRYE
LUFhvwRYxUMbtb+XXjJTD/LYVmXVObpvvL4/taYc3afk5Kf0cCQrk4WfFyW20Cw0/oRILe+lpFQO
iFZZ831jUBGK0RhCFH8xwrIRJSTWQGJxdw/y9F0h2hUcnCky4Bt+XP+Wt4sTmHC9tI0ncf+Ua4F9
xykh4sw1/YhQYvH1doKC/EW1BaC7FCGktAQaR+CNI0h2HSk5wbkJj+yV+EOYBqMz18DWpniKs/Yd
JIn6Zgln9mRQtmFNPhMKqKmBDA1gWE9Ijy6NJdGMhDZ4niGYs2/09OYtwFEBNMWnn2Sf4sNObbK3
ni6zp8d0UvkPufqoRCY88+rNRx+F/pfWeCd6FTilnAs5kX7bd5ddVxxjIlYAqNHSt6KeTI8lf8ui
AuglQx+809F8mOEVCX2BarLJCK0EPtAiSZVYmni4HrorCGmX6fgV5OJZju8fsuxYMcJrf3TD8J+6
tEsjAOl4M7QNHcF4RrO7vsw0gMprjx0JKKJFCcLkEibWD7/7I2V/HivBjNqzQVSzEAhmprFE+sT5
mkG60kAkM7kYRctzYmc64Qp71CuxeTagmrjMuJy0uqo32T99pteYlCRTG1p1TYa6quqC0Slor3J7
e6/Tm8Z85qJmg01tHy7G2g8SD3UzLsXrIdRO+Oe1MdAowpmg6fwuwWMcYQizqvi65tLcHHsza+eU
uxT75aWl1g000kOooRwuRZ6/cnEFyKV0ezQEWcoZh3eisUlbRY+DadMlkTm9yvHoldWUnwQhp/zV
GajT4Q+BCBVooYFwGT929sJMvNUntGPSbBCrENpct7ZZVutuqLJQAkuZFGxGBd9TdB+lxPtb1+eu
OPqeTZ6N9mShvkHnmZJB0DBnkXUCNlIqyPjkF7wPPMo1cJLVZ6gBhbTdoCiMC2P5Q4HLuMQbaxNs
XbDzes1Pe6JAAiC7T6veud+Iql7prPF446xTk14I99FOM6jXVT8Jj1xMxeMmpf4VzdlNhePyHQKm
2iO30qWxnIJoWqcKA4Oh8YXYi5Ug4z8UdwFjt/+//Pt1BxbjL7MZsKoCTiwyR+i/ahUKfD3i/V+v
ZGlbE2q+OyUM3LSbaAuMFMWelV1U7ic2YmoODE4t4ffSZgLiJMfY13iaRmJhC1Od2T6kQ+A22CNe
F+cFs6HXxQD+1xbHjC6BxpQkMGYOby333+xEBmefB7vUhZvD4bx+fupdxfOr2gRgvR5PoQiQ4PR4
fZAWrztcXImM25iA1UKcDzdZUT4SvzRBRebF5N2S8ozy79JzD5pkAi9VwJaAs/pabsO2nFY3hiiS
cNT0Qoe9NErjnUQXrY2HBw/k3fFRQul5p2oQwDVftr78KMWz1DQpLOelNo5vRgCMuoporaARA6hi
eRJh7+EKmcVpPQrmPeEY7LjQgtNYbE/V5/lMiO2UjiTiFO/HQxu8u1cqSzQj208MbmieMM9xk0an
PPeVEDD6V6k44y74UGsy3UjK3GRMXQPDlegyMImQWxz/j/i9xqb3vSCZRVFtA1XT7jCJpnJ8CQLA
yU4GwBRCe06NH50PR3gKIYqPznPV4GRkayyswrBQL66ODhWIflX0QGdR2NBNNxIZF+w7rwDzDROi
gdwGtzBf/7Vu1MforDibuqdP/BaBD7Y1QDVXyG3IoKY2jeIKfF0vyjDKEue6RVJcglY4d2PP90CH
rmU41Q65+PwKQjHQOlpxpwhl7m+pLynLAtir31xUSJhYE3g71J1mOsHzUxK9BGDYCDt4bqoS3SC/
xxXugvfA7dfgIIr+gJ5dQ9jQVFQ4u19dQWd7vat4TyjlWxf7o65GJrpldTXCBEcbXq9QQ082XULu
qCo5ikwWfuhLqxvOWHG557avTTwxDpuc8qJaOkRpMCVNcw22Q9n/g6cKoMTkvg25RFeoob7t3MyO
mdBuOfxQ3QJRPYeEMlORGyVDZS/FwmRtzVt2nA7+gDIxmyQBu3K1oWPlYlm+b3w6uJmuoOMyvp2G
3n3nhPJFj6j7krXcbO3GAbhBzTeS8g/hApCxir07ggbJdxP2gZmdLx8DXfTuWicySmQFHOE9nv2Q
NYmf+gjrl7dLl/qzHXcg2lyXGez6bhnfRgJWryDIaDMxn9uSICa944qOsgt3l9rVfYfsm9oFty2u
//tK2j+l9RNmU/V6sTulu2d0CL82qQktS6/F0FOr9qjWHgI0bMfw82RTKLhC+7I21Kzrj/epev/n
yJZbZ4+JuZhaLri5w5oeCCrE8rpbGdkBdm7dN5y9ppt29VRA/AO2AjnbV3xqVTq5TQweVatol4UK
C/yjTBxy+fb+lpsswDQstEin+B6yTAkNfN71cwnf3XHK0R95uB7LxrJASbbdU99QLEITq5q8ngd9
shUbDgbYCF+yQHcKwU6az5uhZs4k9r//CyFSniD/MiWC9vbSgEmgBCwsxMfX8NmiCyxY87FYqJ0Z
TZluUL9pqb0mDSkydU9LBQVdSc8tfYUMcEfn7vP31kIDsNusQfwW1u0xq/4BZmMNCRYRoKPZIVlP
qMSsOzcxGivfaE0CWpYtjBIYVKskv/FKkJicRdMMGgo5IpT/2d4dejnIfYu0DNyLusMl32gnl/7h
cYVyG/fQLjA6ijsxXND9nbnVeY1F08rSBvJD7mx7X7gSoJpfovZdIAceLF89thno3bLZzyNnPJxn
xzdLsaVS8ag/FcO1mN0kC/SNcWpyEP3tK+O+l4i2JcvN8JATWodjXHb4aSi7l9MFFQvrDzCgBbGS
4ex/wvHTdtrcJimN3j6zr3u/lPfVam9hLU3qmJL9swSsHgM0xag0K0I7btF81sZD0pKVjQCggB0z
ZxSXTUq/TiHgKN9Go8DQjn+WjZG0jwVkAVNv3N9mYcdLDds5BnVnPSnficHmDMkTSf32gaMwl4HT
FznJiSTbTkCZd2qMHYvW28cd/2m1LqyjYu6lmGvueWckA9gtSFri8NQZ8ew+mBloTDwJAKfFSexI
M6Ztlo/V3Gj7GQYCt87LKqoliYW2rPU8MIuwM0ISOD55KNwfSu9MJrC2K8EOxKDL0lIkyG64mHoZ
ijhY1zlBc/yfXnnIuTF2Wz1s+BC+MiGkreVfQSbQSKcrJ5KPJT8Zdx8wKg3kBRsKqwalGA9QHyd6
meHc4eWfJwAil8rSG1hPprtmRaM7ryBjOgiLM4DpclfKLn71s1pTjIjnAvp9LIVEhkIIP9vI2A9S
uRARnM6Uu97MXDghem4b/H6psgAWmVkaxOc4o7v21D2y3JzCrxhTfo5VrcTXn3NuSkhDtp3o8BFB
YXp4lEwjt7vM2b6+i5QteGHz7LnyzGKXOpr36c741nZKM7SetcTE29nGFTnSTBodLS6UZVjonbeL
Xac1uibpSwP1iIR9VUI1zUtcRFr4vgFFrLorjBfV413GtTfz8kRrsyk8cRwFzbbk+sjeV4Uo028y
epngxm+O+jHolyvqYFeHJ8dmDDCOaUPIQSV2XmBBE25tQEzr4Bs5XMWz8esW556OmySbQXjl1+yk
xPUFPZDlT3Z4Niuc7XC1K64huVOxNpa9Pv0OEjA9V/qrUgzTNrn0hGLwcwVb371CDzPv530cBSr+
INlpdvkZkMpfn0pEAnFuxop5zyOI9d7N3T71pr1y+puSnHEU+yvmSKRCWBBvztSbwBI/7R76STNr
JfHpCSXQNpzHuCM18ZQ0KJRcgG7YdVMB67SY5+0CYJ2hgWksLDo2OtlL+cql45qgix0tqVykMuv6
uyZFRH3sguoUjms5EbCwoyIfoHSkzteqPSHVYCy4LtIEFlWCIeTQI23Wb/MxvqqUdDe2OsFX3xUD
3S8nIBlvHmErwjLudVr+StJyoWSbNau5+Wzlj7+C56/HWA2++WEInAXv5TIo7M27FgImQMZd6jQC
uuq3epddjwHLKLKopTWJpaUhdnwh8k4fDa0nSv7xV6HZM+kwhhUZj1OYO0jWeIqewOkDIazYU3M1
/fwkg7Er3qI2f9h23Fr6/mB2LlygQMIxxWbh964tV4kWfiuA6/gYhhmP5sxamsfHam+/UvS5KTB2
JNaVUNcf2YYtcjmyXGD3pxmqx7+IzojvcjYYAIHS3Op7H80h3PHLYfcmJLyWU1bQWhjt2Jl6Br3i
wcyfiGEVJJZdqCe47rAMJd3+iscmxe2JWfx35090R0LGStrkzCuBqCXRk3JCeHCJ4XCwy19sI4Hh
1rsK7Y0JiZYnIx+AW35/2jvbjh6PjDgF1UfxRttquZ7TFuASORYc3eDZqmNzQx2ygGIfA3Fd3Zxl
qOBhjJtrXf6gtYNO/bOoEb2V2N5f9EGIZZg2UWTcPLPR9IEL55606LoOBz4D57gW7thMKIH2PoJx
hy9MDaJfEFDJqzNjtTTGE4U/PvHPrGjcsLaKVhsu89dretF3Lu6tKPDU4vP5Vq7yI3+HpNxMrHk0
4ppNxPKw7C0as3Bw0C4Az59n/rYtmLA4YCSrstkLHqc3tLjwJw1YQJAUee6FZ9LvFMMkbVZaLpJ7
qmLHFapKTdWG62F1a6796HFYQIM/EySdsyl5yCL7qVXZhU+KJ5Bz07aMOUvSYgNfGuQOEJHuSCFf
NJWK9VVX3pcWfSpXaOCma66V+Q3k47Q3Jni7BT0P8U+d7wsqIg59hOQStX52TVXlT8lmtcrMy2om
ZplNtupRfjv660VTCw9tIFykFQrrsFk56VedovIZnxNYi7Dw2MxRhWN4hR3QRVyVXHJD/Lyc/ffQ
DKOSyG2IopJ131iyLepew0PM64We2Knznxc6TrNBgXKl5pQPOvDqKea/4tFUtAkNUAYDDEeD/cXf
mQOId7h9/lnlOHaA3kuxy1WqaEZi60htrps6J2zIlPakacyOyjE6KR8nhukPuVPVYGUJg0rIo/k7
wIy/SCJb7e6SgzRiQXYvQpwHvp/jGbqrVW2wBw2nkrnlPp0a2B1Z4yIzvp6EMWGFufQFBSPrvcuB
AhxXnVaVWCQb37nkxW2LrMQqC2C9NKl6xiCPCEqvy/9SZaQNINYD76K8WM2+r/vacYECRboc7iOn
wV9LHF6bb6mELCgHy13NrwipSah743NIwt2biia4h8D3fCgI7oU3RPL03qCs73BjRT9bmKzqvxqj
yzflWt3ekSWPaByXdsK2dimE9W5jL8HQUHtGtH8pPcanMEYiAibZsPffSYPD8QA73SShAN3g28HQ
RBzSzaIaXfcFQsNM/Jua8Ida+SjMoeBvUoLmg9dxorhk/gvWi5wx/5dfrveF3T40m4lNHpz2khBQ
lg+R6d/C6IRTU1Wu+AyDM5xlNCm3D7BKLry+1OJB3mXIScS/GHxaj6uVm85lVXDW6pGHCR5zKQkJ
/wki7MK0/0NI/qk69vYfhd2EVtEcWYBwm699pdlrjyWEAwZ7AwIjoOvgXiJL7TrYy/vs0n1ZRjf4
qb5NyTlYii/5ex67+XC8TreIjnz6TZUq84b1NjY1dJoUm2D+R4lY+vuHWlQ+KJ6/qlQmOXWRFfP+
AiSvuAml7dCCSywQaU7ebRlqZZHrEmnFv6mFePGV7bwmjtWRLcCvkv5naUtkth3z/Ty2xHSFPiLN
qbgt0/uyk5kCLKHjHk4uS4inXzDL7Hy5KEbmexoUkj4h/ySqQz21T5Dz+o51lvlORjz3qpc7gKL8
I473jKVagvoEeN18XJr9py2B/45wy/BPXbyQwqSXtX6Borolz3hA6OLeF3uruPtid/oP/nQ/6Nmk
T22IAT7zOdjXRbabk2auZ8c6UTdNmW8cuJgkxNw2FufAfG2WxRzYZfCrlBBFtg0yLRjocljsmbAp
88EwkKBy4+QTLlztLFLn7wbD8kbsmb2QwPwvpwk8vFFm58zfS3doN5u8vU0MD9Q0Xi60U05RhkJ1
UMPgbMuldu8GHpgGCYa9IRGiq25aQMefRWwKdcivr2fUGX30803gad0Lj5+GlgKAf0y/MMVv7Bvf
WIRYkjQCU4Pg5+RLOBSMfypKuTVOb2h2z0zyO/1Q07nd5+txBxNibmbHV4MQ0+nDuvphZypds079
6YHz+qn/GDdKF6CaUt6ovzC88m2b/wXatPpu+qsQDswJEvNIhkDtcQNkoDtNZoOmnRpQLb8FiqGD
9wyy2e7q/onFfQQ28ZMEvL01YoQI7dFw3m8QUYtO4Zyy+4746sK+evzZB43TpvfPcPoTHTjaTi5K
fdNk1iaoMam0XNdO7pKtVy5SXXGGw9JuvjipT/GOcjeNk3rVTJlpAIcN2WjpcgnifX5rxULpKh2g
kanD4rkz1knF5L168+u8EY6d0zMPT6WZTUA6bUP6yMJYN6TkLCCsyMv1IsiC3VzMy0jRR5JMj01G
GlLPwnrves/f0o9RlOcaVwmOdx71gFZIdd4mNvzY/SdShW4FpxaQUy/XglS/VbDhzGYftmTGhTCb
ZvD7uLjRUOhruTYSfZ4b27XG3W5ftCThSaZ43mthWIrhBlN5wTh84O9wX3IpEGn4f8VvzP9vkMRX
1PByhvzNHzsxmIyjCv25ERa3d1j2ZeE+p0P6FwJmzFFougVkcTJB/UaqkzNjEiu+oanZjatP0iyz
/9b3Hg63TMObWAbN9S/QCmkcJ5n+4tegXe5JtuBZ66+H+nBUlz9Df4Y0L+pyTacpK4XzdlDUP6st
MWPfXP54CPHHaRDt88KOejwNkoIXfkkwJJ2FK46Lj/R8QHAR3iANQNJ58UJrJInfk0Xo5yJ7HvEP
gzvLSOf/xfS7p98Ere9WBmYI0IYMI/FGoHEMcoGZ3IZcdTd3yvQg7pw/qTdIyER1sN5yblLNWUMd
1oNIxkk+344BpBKahQst+jGvSRSJoznL/RPpcQMMzw2t9bnTVrLFoQytQzOaE+NxNfXvLOTe3odz
Gm0n0MsKHB74UuuvF3WvzzVciBT0KC5Aock76UKFjcLFSp/RDg61T8MSdyFCgmdiMCDiSNTnMOR8
ePxuWcE8a1wFpZoZSRWRyGGof8Q/3hQt4Jn6NoG/Ucvzg/nDRqCeYyhyADqOHDtNN8Ob3y4uhMTx
zNhp6uSHuy9LLBj35N8xp6x4+VzDc9BvwYd5BB3HO16Ml9COQziAJrMkusOOtLW9NDXtMrD6Nkkw
qYGpKTKpGNhFhFbJ9/gyUAdzO9KZHQFBXNU35FkL5fO06xjawvdCmpPBCS51HponrY/u4PkvNRB8
pzMI0WvOqWUWDQxEsQfkG6OIzTmlQXn3juwC6k8ptOk1BbFRXizek60GjM3VY1I5dvqaVTYBHVyi
9wEctuwidR1svC0aHPFvg+8lVGieW4sN25CO7FlI7wHtfFe2vl20m+9WaycmMe2m0z+GzTY5eHCW
L+9pfp6a7UBtfu44gneUmesqK4nbm4QuFSQ4Yum1+fSfYT3MP6BR8MiCc0HTDYK88ZTZ9HIgC/Vz
I/ULIN4tOMST4NMQePt8WzoP3yiRYdISMmPQTik5JKp4CM71stf3Qqaz6fHXUJXfkfU69+0O9NnP
ENmxIsjfmG+8GNF5TXlgsFeXGzNod+4TuNQb3OWP3zlkDP5qU0GeVl92kjcHxeveZ7UcB9RGpoli
B9X0C8jpclukN31EYZv6XbatoLvZK8igN/Bof6g3GJ3ETlSj+aqL/B+JSLPfU9UBazvLhWoDAk9z
nrLQk8dlZInqpw/q2a6HeBGcB0KCt/GPezH4cKkJS57tro87HoEN/LPY0Xa2flB7e1ISXfCfo4eV
/QVf69X2fwF3GuG8lpvFeR/0oo7CnffiJSF9oho5b/daqFCUgCBwGuXXRBtXlBs+cQDswGXPbMeo
T99e4+EtOoVDlgoqsiZq6x84Dbg4G9ARDXXfRQqf7U1q1Iu6lbsZyxFfSKxiANLm+KW+7Z/hzhZD
+KxeNpqUmvtl78lqWlashCBsNcrObkO+EXtz4aGuxqOIODjKLmPDx60N4z8Zlm5a5eFogF4HFiHU
Hx4fD/ZnVvDTdoWWWUtRBVQi9IdIgL1Hl1nN0/rkbOsBiH6tCDShltrdGqx0bNtbI9vn1OhqhJfa
Fwl/wG/qmoLSiGD220f6mq0UViC4WFp4K2sSaK6SIf2uS3VogXhrNMDJAZIq9blMxSOVMmrrtc+j
AdedUF4u8XH4gv8Xz83yZzTeCFgyY5fHPTPyVP+79H6MdFl9Oy0/aIe5fxUUZ0qZioITMzdf6aqe
M78OiFbc3svTaQ74PTG4/qyS1VYbmHcpp9C5oWKgAooy6cdTaD5OW3G6mViwBq35TrU+YEN77Hm0
RmHaRbpR8fWCO8CrpM3/jUyomyWsGcQxe/UgXDHPqrq789u0QLRUv1ZBbJCJ1LXCu6/6A0wEb+Hd
4TOJEC4Anl4/JxFB+vWm35OlckVAbXXuodKZx7PVro2lS3P6G9NvovBhc1wdXeynw64mUU3KGUUD
2i4SXcrx6D5aaYjhw+QUzTLaBj1Es5bcwjmkSsH2V0qFoSh+6OB9JLvm41IX0nI1DsTHn1L30dDe
QOOFGcj2vQJy6Itv9yU8n2Ok7LTKfeIxkuvRev0dYn4jZCjQ7QvQ8enj5WxEha+sUeRz4CQuAPk3
/K3YTvnYXTt6Vv51vLIygLzH7v+KZEphNsfPnBvwB2qb6thIlVFI6NNm542dti+X3xu2nTYp+hwI
jgUTwHko6wxUSm50GPQK1C4M36bDenphzMefmOP/5GGLV3/xSBvKBSNj4O4u1j4gdo5VusTYTe/M
wkPtsDcT67qgl09hdEAzoByiCACaSeOhfGrYI7Zxh49uyYV6TNAbSdeilbHLh26vHT6a9frqtHA+
JXRkluoe7gn892BqaYNNYrJs0X077ByjF+Y9HJtm3ybo04swArqfV1oW1+3BoSZk7ZYHu8eFUpAW
4N3/y4rXGAqRdfBcb/MyyjZYy1yyH65lQhVojLUWAyQF2LXtRrOlfM/2RJKQhRwpdm/o3J0o8Ut3
V1h4Xv1mCkDMRUOoRYa9FGRnkJmuucHchWykhh84X8gdNtdbESkBIOxfqHLX3+1N5bSb1feAJmHX
YjA6OQWzj7RJyh44cDFVoskeoA38aPsrCzZBa7qjtv/abt/WrQOYUCu9WugG59P4Dvsvm8OL0oxX
86nGdPt8KlJaDwu418uDY9rVJVwhtjO++sVsEryb90Jvthn6i89GAtgXXIGJ79+HhFnBm896vj/S
Iksf4YvKiZt6GtuCiNK4yDuK65tZST/UyFbWloKEfCR7u0loZ/l6rtQDM9aA2WYdBC7R+X68/wUy
g1rWJn4B+NtJCQGWUkHHsrDRWirUiZiBJFWhRiew03hPRG7qmbd2k0f/a+uqQV+bvPoCFDaiSoU9
cIqeeRSL0EEXkI7NckF8knZwfNuDvyKvJQRWx+9KgpeFnL3bJhXPF3b0oeicymEp1y2coEBz1944
BNIXx9e+9xjZD73GJ5RKrsi/30+uoV/K7e0b6kE7kZzQtzMnj6CDouB1lzQmv6OdkLB96oi1mfv7
uuurcI3dFFWG3NeqldYerPevMOmsMYbRXpKEE0v9LbOrx8UFni+LJsCYCPe4aZ4stT41J73lbzKp
DulXlMvImo1BPbQLCDD8BylDHAXCCEFjnZuW4e2ui3ntzhK4TZiUEvcwIWf8MArb2A+Khf98P1/R
rPGQGQSp7Ne9UsGG+ECCh1SRllCgYYztG56uBOHbT2VeZI7foIOAmu6M0gtDGWut58mIu55Brnva
bn0KSl+H4DQ4Turd90lYYRx0jFOgREskaFkwbpar1GOpVDL3mBzzYG0Sg7p5XbUUgoS1c86eSlP2
mVqYLczESu4PUZeUWzYPZWlD8QBP5eZq8NDoFSJJaGS4MwtIoX3UBs2kiXLWhYdg4U9QStby/MXs
xWwEtQcoWDQWdJkgGoU1npFF7IRT4OknSLYNu65DcPkyrEDNCcIzCBBKOP8a1SkceL82eUflMXCb
DvdGRkP1n/H9j+Iez0PsxfYkkKly7QcPxLd784zhhZJA5ttWVyhiEUcPMP+O6EMe/UMBWr7FKnDq
ecLP1plxMN3a53GbgwT9xV+FJDOr11ZITmbsdMuW5hrAonDRs9qUpeWLQyfajsPqe0ziJUBar3/x
RIeJdg6QQs2mqHftqhOjzbFCQYFlU8UZJ5ura58QCLpIhbvQCkEgHsQr4bRbZ2r/ufm7d0MeON7G
OmlXdnmqTTPY0oUq1r6HlyZPRyBw51vNOqzthVasKEqdPPSEQzYnm4aw9QH+U+mwrvTX4ucVN3Qw
un55ZDxmY1gpJmm+ADnd6GhP8FVIDRWbLEGNYz4rK2xbN/c2LzZGEm1TXPUXsveSoVZQQT3MGNNd
UNeudOul4dj0k3SFTnimnXsXrr5vXouotw5C6WFTwgtWfI+cgABZaALBK9jn1AIQKBK8SQPyPHga
ipdQWBJbl+5y69WF5Y+sc9h319mRUczMIj0pFn4u4U+W9f9M6tjIurpYxU0vKIauZWV2BEsoj3/C
lwE2RNZBF26aTStfgd2FoFNAFTHo2V2ZXHi+ZWx3tCIdOIiy16Tf8BtUA0mlG1Lk3T0FcIKHd5we
3/xePQfYn4zsX9Iq5qs1niJhTQspDk2F9OKWQykXZdL345TrRgc9AIi6ggJXJMeR2E8042gilwWs
53HP+YIdTy/HWsmOBbb592zCZeDvF1u6rBMJhgDD2/ySLZFcfrr7eQAcr/crndGST8mUxYUMsh0U
4J07LRNIW0fWXjUiCg1piZM0YH0m+AK7JGzhHOcjiD5bsqJ0yF48TVvSyHo7/yLyIrYtXmTmjG2F
U6RjvPc3dpedwXpXIV3bjIdTY9PDYHKAZU9hmz9i7jLeANGxfcuI+uZji4nbM4vfp3VLSsyo3nkV
b4XfzyzUTFC//ki2aS8iLpfK4JrnZK4u5A/XbpNmtuxTRyvXcODRXUhF0FBIgJKTiNTiTVlnHg38
5/UV/fOsUoWd3YVLsCpdQYzCOGMt4YAlQPDORHYrxMO6gX40SQVSytQ7OXLbEWXPY1zWtt7Gg7Ne
nGeWzm+NqLVy2g4CyTRoa6MvqLXgWw1IYvHr8IXJCPDe/7aRC13fpexNHPp8c28aP+zYm/CK2ZjX
sRLzWjq/1yBUBdOfvDsOCqNy5f9jPKCK63E10cIHbM3Twzi+OXCOBd3vGjK/oyFhNrj2pfneZWkw
HINzIXKpXr4Z3/dGVNEp00TmOqRjPO3A2/xiytdpwKWhnrLC5QptDjUAeGP4Rgyb6UBw125ZMv/t
008V0sqoeotzshjvR/2/TLMclcQNFH8LF+EPddiOlbUS9hN3TlEXzZPTjJiPbHZaQ16EBvksRzHX
pHXWKLXfdPN3M8rPzVoxC/rVKbjblWBwaR+Pz+iBy/kOrFZSV0daFAoG9eKSZcL3BbaFgkgzvr9H
DKJScVjXPFbjfRQvwRCoHKT9rmqEflvA5Lp26etgIDZk3Pd/qr9uQIvxWnM1njzcnXYj9g+X8O6X
5rK62tvGYBgSj2FFOp5mOC/jnzfTxsDT/ghGgOYuNgyYdY6s0Wd7D2AYK54bCmx4D7O9InVzfcOW
Ag76gtBBCYrQo+UooBCjrFd/8HYo4JHgaM28twKCdyk7PhIO7DDhgp8gMQkTFakSrRWuUTI9LVGT
2O1YDFPw7t4w3rotuPBSbeRGn0eunaJABA1He9ajibnHas1/YttQDSSJPgcTdE/Ncn1WoijB8geG
7wEP0qWn9ld1TuXTI8N1lhVl+ecWBzRhNAZjBYpNJ9JTKRM9SRxP2Ol5qjfLPG6Vjt6/yagvWD+6
hYAB9DtqDpEPD0CaBHBpKuxHgGrmoA4RzFePGvD+ZIhKqh672JBnvGyMeC6ImT/oFkHWxRZ/6cQx
MLpPxFfg3z+HaDgH+vzGPKS3PId23WX961mulScBlClAF8bHbjEjqx6bgpmQON1Yc+BoOPmdtpp1
N4ZmrQJLTm2y/QV8+Pb5DxjHKmMq+ngsDIKTSKyc15rm3Qm6HQnYpQVrGlbXtT7nLGsEg6TiN3Cx
UzBONL7OtNGPYTJsZoKfvCvXtuil/zF3yDsWu04uA5vrJUVSSljFcFSgxF6cObiJGtAYjDcumSSU
dXRna2PmpYNqUo/mpvgL6z09ZwGPsJYfzVQza6rJmvC6RKRrHxCYYDtFwAyftGVs+lY20Gj0ocpt
RwXPjhp7TgPeufJQWWPoizJ5qK3JsJM3uzmRzS2YsZtgoH8/3DguzMhmZkavcOqdJQXqgd9dAxIB
UN0nG9TTMQcyBFEMOfB2KkukR4IXMihHhcz6/85qkV+yIeLdDAPnCl95kQxjYlhAVImpdYAR/3dO
+2MXx0J5JO1lVNoW3K5obXKonh980c8kQa4L/UHSdStGq4vnvYStPgfRP4jrDM9egbeIZm8Mv7ER
+ERzdNvd6/vJcS4W+pMsJ2aGhj0gqi1LlkaejWb1gIRx+yCbgVC67iJEJBpNGy1oZCl/4GJb6vhs
iBd9Mn4rx5TsX9oq2GapCy7+34G2QRkjC6kZCIzAWjHGlIlctPajxurXf2j+h0noc53zJ4W3QhGL
mqgvB2EH5/jDicZKCixsEXfRO7Yhzo0CORrobbOKZKu8tcfnyXvL0agVxjRCkApni5QRT+NfBYj8
Eicc+CPCxZsNn228WjuOx3rHr60H3qfowgNXNlDOWtOfjraN9zq1Hze9xTp/xzF4toXxb6LsfBlA
11pyb1aAZKXosFRPeecN5urFtcCTvV5fzovtO/F6U5g1Vkh18T/quuDCN3pBlNb+Cq2L67+tpl64
jBt9cWJTzO9PKy1t8AcLGVXScJo+75jmHVvlJeZwyZ6QLna3g+HQOsk2yRsMbIgOFV/HPlKuO3YY
fFqiygCUp6b3A7fY028ic7vFB5pmfIPlNhTxcElgGSF+vSlrk3ajQLFnYms23VUpgzb25jcJki0V
UIduBIuBae4EO2XZpgWNP+OlTDi5JtzBHQB6w7i9fyWspiO3DURQIcoKxh5kM5OVu9IaGBG3kD7d
Bhv/iwTRF1q/dP7tz7ygQzvz22GN7ABlt24Wbv7VMEa1Tz7s7Geiy925d7oantg6lfEiK3R0WuWg
0lrHR28M5RGt4qImI41vOrK/iRF04klhWUgd/fAjU9HWCFGIq9zGun4kP6MsS4qUHDTM+p+lwah7
h8E2+hWNL1Dj7aV01Sl4+tbu6hY8974C1pHkXEvfaUMCuR5DPdi+w+DpYhjLPJ3kydNYV9wydnPb
xbbRNcb/TRmIJrjR02zTTO+jBz9pyslkP+2owOAFVSlgUa+IFk7l6h/BQMefyQYVwEyQ2d8Tgi3a
UJQFqWs13bf/cYpGXmNawnT3udoOWJ8x+gMdhXq/93tXXP7cymnxawC8Lc1DNxQfpQ5c8YMNPmwj
wyCh7gtd+IiAuOwajj55Hlpo725x0f4951f+PZg7eGFFzRe4u4vLUs+kMZwplsIYLsFllb8GFVEl
dQSjreKJlrPANpmvf0taIcG0TIhf/dYtmw6fC5n5Iu5qFDKDJTU/4jsUXx3/PgiN4TEPcryfSRw3
K63XueE8GFwFzOoyh9tHaUDh+vnDs//HDF8XHV+4e+35mgGxAjSX1gWHLTpqxDecXPR1SIGbfloN
QHwvhN16Yj7OtHGiM9VEPO/Xga51sIO05vgambdLq6u77R/8V59mVBGnqHlXdSesFNUedNFEGMSJ
cUWYLbiNszaCc6CLI341Vtpfq/qIU+dZJF06qgXo+hznHWkMg2d6/uciX1Vo62OKoNydP470vFG8
dLUvMrIyeyT3kyGEFmNvChSwqX7pneLcSRDcQy9v8uRHoN/BlvaDWhKjK0wuhtUPN6oMgaPND0R0
ajtybIIv1jLxTrUTIJXXxT6WoozeL5iVuRuBNTegclFW5czXmqPYuXmFSPYUGBMs7XMWbhq8YTCp
XugjlGVWFG82H1oNyqK6//nfIJlOEeydXtWNFMMTrxRUc2qJ4LYqFPiFige4ClwdBg4ORhqtigbW
WxLkGiAyu9ilJOGGx0fIQaYwb7lle36BXT0Gzzz3w4bzmGGType8SAFmysD7omLrNOBtik6XY0+n
MekG5e6xHeu8fWDDGnK0zJzVHquqCf6Ge983q7KtaeBG/kRTtKFuHbqg2EsgixIe2j9LpG1vsd2V
5s1A8PcVljC98K6ShMgryycaROVqw0gL7UvljPy/eR52Z6Qi7aLA/r/BZrOkVR6bKm6BD/rb+a7O
odQGlgcTXtANiSbP/5DL7j0W1njOplZH0q5Tgl7Tf6hLsyyMjMPRLzgZm5cicfpcqTFiRsDRbyWa
ejkyFsG8XbRs1fEgBJf0iU4KyUW23Y/h3X5oRRl9FgzKTJuZ+jIRlJfetUGeGpQYJptVoBs+SUdl
XW9w9+7wgJpnd7ELdAlWVvfy+xXG/WNgQe5za60GUGB1fAM32b2qXOc0WG/3iPhC/6cGFEsorIP7
h4rcPMzdnmtfSBOizAL4JF6SQTuYeeibMaixHEWXu8Iy74YNzit+uHqeBC3v8KLJa25FHXCJ5XAc
+YyH0Z7/vi7+tSNdyRa6WOVZISN+aj5oPfkHqIded/Fy79Bu7gJSE477EviatrNDo/7w9dH6qVHz
+e4qYr5iAqVi3iYCDquVwfJeZDdMIQEslfSMSdbKj+OGnckIhoqPzoSX7AYASzfl1qdWBvxeEdXP
ZIf4wCHHQFhlw4AYQ8NSqVX/Jz7c/dSJRjMIYMKlYZr9SjWApaE55BJwoSAOh7j8B/3w7KvsGXxN
V752+X1+9NPDkXrEyu8gaT6U71yRGh5jpRQr6/bPDEc1jPdZGO7adLRnm5zqNY/pSh1aVXln/CRN
WRiESvvHc4Gr1ZAuJD7/MVT7P04lcmvZJxgFhMoJUq0mZsrlPT7zo1NS9ZO8VYTGHycyW2K3eoGr
gOhXhuGDWdWtvoPN4iBfwhVJ+TBjaFTq1fToivrUIRZf+QDN438kzhEfCL2KJfLZXMS/vT3jKe6Q
y97EpCUfH6x8FHdo6mr+ITGOuAUXWGAkdDsariIaHDTIrnO4tITLg5L5fks2DmpTuWmq85B//5C3
jkn7gFHuc+IDe+paSoT6++622aTu88HQdd4vXF0KsR87L8j1Tm02Bf776n73tny7Ku8pbniWjNHT
FEP36/+GTLtTuF8gWSYQ8+AD85uaMJ6Cn7RK2IN+wzkF2SbdZTI5DA2DOzGXlQ79MhXv1rQp8A6M
93FpaBIgh2PEfsT1rzGqdPIyBDTJT0G84uvHWX04k+c5ADFvVFFB0Gg+Z5BQNvvFl0gigcYEr2vX
iEL9+vPdIxn0COBsnIx6K/NT4Q5ECyX/SGSXSWidZ+y0ifzdShiX37MlafrQ/9XjZ8vKrt0nLSFh
7XGhde5T10/Nungvn1r9R0alz55T2btQHnsIWYffsxz862dpgMNrchDwHEx2s9qilaOJkvlw6Soi
tXYmd326wZFYHyAXSXBeoGebq+U+1AtBQJray5Aj+JlfkztrmacVSb6UFlUtTpf8oSAQ4+jiHI2T
vC8CXhP+jWyauBpPlTEGt+XipjeJJWRxFIF4ztU7hRBqg6lYjN5ILGqNGRzkiJmWN01b9JA7nRNc
pZCMqt56EVW6zx5YBXN7Z9C4L9Pecjrephyg6eYbor9/qaorr1vPSCq4BEAWB5Lk7I2Y+z47r/tC
66hwrC5AOwODWF92pMVNlP/DY6KOfn2ceb+6Qc6+qsA7jAQjEogA0drYR09Nyx0JMIqm+ocVsefp
o80R3Ravm/E2/lwON5uUPgmNVXoRumZ4a8LTInuVUmf1sNpq8HbBRkjYef+z+Ly7MXhkzWEq8+Wo
Q2HelfF/aibnJPmvZca7PFl1e8IxW4aFjqns1gewhjCpkcqUVkEiTx5eg+Lho2H6B5o+7nf6YsQJ
+KW9rYKx6rdhiFryEH5znxnNzZTp7YxZWRAkgduWgWBkkTZM0IDgn/xxI9T1dNMGo9oikTija+qQ
vQ9nODrAHOhoAaTlWdFivJrcw4ALPiZQBBJf1Zpim/nudd+T37/26y5UMzMJ1N22nE8N/PhFtpkP
hcIaMU5mG113kiwgkqM9/dV0YZbDj4UavkoaWfwc0l8b+vsdUmIB3gOP4DUxfyxGJ4ethT4aYSec
bfQkeaW0/agwLD+mE3Kz5EeqcvRotEPBsTkpmiUytNCfJxnO803Vg2VG84pu+cRjRRc6SB/NF0pP
Ix48b3IqrQZTVg9PEXSZ11NWjCbK0/4HjKjh9becl2gytIc27kVpCNTDdAUXnps8AFX6w4YxGRuQ
WfGwJxic3RWqDg/+j49nep0Yq71xDSFghDv+yxqbg/U6SdMJvIPCsA57hLV2V9a6qSskoksQZrZB
hgK/Dvw4AaJKgXRwVYnKEWyNKlieM691CnpFR87bHU2wDcdZrLNruVNEzvAZd6aVgMfU7OERDSSN
p+LcKRDLl/rS8TdR00Y0v5yaIh0CR1Th4JOUHMjgFJ3OnhHKoL6Iw/DKDCJeVlSJy17+9Kn7brNP
6rRFfLlQ6fNQA/wMI3WH3kP/MMIuoPQtOywwyHFtw4+hrYFYC4+vIolSjWf/GCb7SPGizuZdlH5j
0SG5aFgAl9t62464QLji+D7DpxiXMrrq4m6YVmWZge9h00zOHmiWVxS6V7JBHp5C/SJqui4K+GXA
bI3Fbu4f43EMSweqTRWy1p9cKBcC5EoM9vs82TxYcX3IQcM2vIhMicavNXIawO/wXLJ5F9s8nFGy
+emJO6hwckuPD6sTgPgtAsK5ETKk0294dRjl3ASiZu1rtGVhW0Jz+oBlQq/ivT5qheE49sS6WO+g
YLUpYwKDxXOlldNAzO5quaAeuZRRNHn8mtJjyiEEZlO/kaWH69X/Uvns5KrD7HpZ1D+O7m9B7d9k
f+ThG/ueBD9GygmJz+iSWp2F2H3i78oUhANVpGZ61GGJ9HP7vH4X9wIdSyl2wCsiu2zBt82uQALy
DF7yAkt4cZCyCTjfGHCKIDQg/M4vkpaJIYMfWcK1hlt5YiDfdTocxed0a9DGCTbc1K5VXo0Xtwzq
JnCSRWVowF4UCFbJgEsy9XThnfM5fd+yWDA1cN2O7C9Nlv/hOxP3zPhT/72Lre49plktF5ihrq1n
SNRyu0yijDPhEO0b8KmR5GFkYWEW61SkKl6WYeJWNKCwFe81ifbV4tayNWlX0cxW5Db/0VFt1wIn
HEEGgG7JUFNXgzhbFZQRypKoFh47/3vX1iWlIt76Ykcu6++q58Gcp571aqagnoh7tWKrtFAwbG7h
7HoAzmGe6yxHam7a+BcLMgUzIH83rIzALHl/EtGfHebHvGJ5qVdwb9PkshvGwCbUtZ3rqpoxlyOM
7igosX8gSXGcRQUYBfdwJCPnoHw3ICmG16/oR1JcKStZkov9FalNT1Wpr58HbhwlcHKRuSFgT5BO
0NwfHuIVF4bIU7dDPAFvasI6CBQ9mIhXbvE+HxkEsvXvIcDwJCIrfp0ZGOMx7yV7lugPczHnQN3I
Q00M1JDgJQJWqPaByyOSuXwo1lKNG0BG2ujmVQ37VlsK+uNfeQoaFSNPShIr6a95sOS1IiCoNBpl
LYhZLoRKq7pK7KqD6DU+8I/4NxR0h9xWZZJBiL9qt6S2dVbuDiNbFylLntlyzcZy0AqYtwzMAXp3
mvoNipi3TnNeatIacnzVF4CoukH3D1To+bO3I3eM2W9akYVNyjBe7eRAbLvoacUPrzFfFapuY9dH
qoNo6Fh2lIR7owHR2MCdhfshYWFgvAbuBo0CggGz4I7XKMicLL2LBKJKWRmvaG1dT2FGQUfEdPoB
NqTfXP9CYKILywTfoiScyL67hSHZE9mpo1Sda5aMmZUrUp6W+z7jjT7+/BAXui3+95TDaxKlT/eD
CHidT+psFyR5PjjZJuleaxVDHC1dDOlxZfMbbekpW9l60wFEWRckoxwsl6tNZnMv17Iaig1teLAM
jox82fC1uBItldIxEKQbAti0R7z4pGs4SDOfaJEIs5vAusHCNFoXRsh1js7rCJFR31uAgHqLMFjw
zxZXdCXZK2KSU43u7+SuUvCQO44Snmtb5cfbc4Vzkho8n433+ovtyGQHidKFtCU29uSuHAscUJTe
KRRjxVXuPmbRaWzuMSNIRJMqmwT6dZ51RnJTsrtKasZr7PLSreZ8q4ShBHKcWQhzIsQxrICLMm1w
Kx2o/FyXgs3BpFlseZUWCYMbru21XL5uaCdzzzvPEA00an71I1iiaGr49Tk188wr6Kiq0Gp2UPJn
qV4Y69NZ5ZnwEXdMfDj2IMbPB29cCE5+sht1Z+BUO3YOaAbIpcmaeni9wamGWg2er67WxPoE6HTw
FeG28VnPwi95OtHJEPDv+/jLX0ebwoWOsUUl99sW7j4g5BAEwLpsljl3LGHgKyAOcVhd91tKTSkc
Ox39vVxDzHQx2S2oLiJCp2HkKQ2e5Hed08sJrlccRyCHdWqZ6oWX7BHFtNukrWKHLLGVZ38N/arC
f+oSE/AUdP1tIczCyCnKZeZod/RD4U2kicJo7pQnCfbdrkFdRg3cOcOK+32Um9X8E1g6noBgvsnT
4p2srS0p88LXXkqegrxzIE/TJRU58uHAluDDWhD+gEr9NS5vzOtO45EGIdrbK6mrRYCJTdxOY7vw
BJYEgMZENZq1mMKVVzoNo7+Ca/u/BKLvkI9ec0jzB97kIS+599/5ngMeaeE3nSB1yafVG3/bP7uK
QGRQKVXj3rzSlgBLWwKFXl4DqYVJsKmgK7woLD8QEbCgyXwO8b2ZrUrPoU+YwG74A44QUJb2IBFX
qtLGYbjZ+EBQ/cZUPTF3pmnX7XlO3wtyLWFJj0GnhVdefk8vBn3lLOBXcLlUDMxuGRHFOHACj1nI
5UMvxQz0TH5oNDWfAXh3l7wfvvm5MZYdfs/sbu1ELfZqVjQCzWY40KhqdBJY0J2AG61FhmD04yQg
DIERytXfrag3GC+as/MCORMtc6ZYrh1KlHEqC3Mbg8udON77aegpvWg7ErPf9zufkGuATRKS6jGI
wtuvptJXOmasVMlIHP6lIRPwO+zdujpfWbNzUKcDrA4SrO3JDnkq333SpNrat4Z5w0XuFMLjAN3y
nZml7lZY06EQfx0b4iBHz4EC0FtnIslX26pW1i/iN90ImvH/bf2jhnWTuOgBh8vVUTiga0i79DUa
YZTUbFEf/iBhVnwYeM3oxqZhoKXaLwFAMFPLp1036Y8jIVlS6mdgSmc6uXUiIKbaw/E5zh124/9I
Zi6woeV0vcbUnuRtAcnMGhNu4NfS/KSZx0ydzl4vFRDavBScuW7qZe6CI8vWXm/MxdMqbEsdK48S
RJsugt/UbxE8JOOB1Z7Y87pBjFbcpTSpiwZnkAjjTjqlzzLmxtFR/I2uRyRmzSHC/brf6DHB3tCH
4UvSoW4lVzcT04Mgq2A+LutmoEzeMCBoMAa/xDxrWeyJasPXUoS+vbRtzKiuuqBQC6BWoK1J0Z+4
bDzBwkZb6c6tqnjOIqj4QkXU/T/fku9tkfW1hvFHmrKdBp0C2SnrTLbYOiea54YzNRf+Leb3kwfP
ioYQaBlQjQJ49UpEdP/N5jhvTjnS4BVqg9znP3xNfVZ/Sq6wBt9sCgh0DMc3ilTJPmnv6vODOYTF
NFyib8gcr1r26FRPZUGkcGPDGCOzynJ9KQa7+iEVQ2wtlNne6gQLR5APWrf1Cl17tkfPyKzKLn3D
Qh+6J4+75VJSgVkk1r79aga4d4m5OyrlaJ7Z9kuJFcvCdyKnuTJRbfm0i6sk755sysQyZJy6UkvU
Bo0mb4ZJ8jmcm4YVM8DzBsB8nkWQ2o3tW+n9Q5pglPm+i6zPV9mZrBs/APwgthvKJoyAzNnXpbvU
5x5iHgGOfQAsWFN5Xqc2z9QAuqXS9ca0qzwuvfglIDJbb/tBCuESnArh7iWVJ1CE6gzZBnsCLhRE
5n1hBid7Dlk0gSIaqHZ5BkA+BkPPBr8m/O/L/Noe+0HEqSH89XrsVqPCNT9Zw11gms5iVPwvoeu8
a4xXhLBOb+ehq2t6j8P42JMPbhsWZk30UbEUrMiuaMzgbNqnfNUPhdWdKzHB61NAGIT12tR1r60t
TFcnySVTU41xnNlmQZvhlC8eNrLwLi3P64n8BOJXUxtSf4B+ihrAgkzZOoaB5tOH3mswkBbyadZi
87Y0tg3ERBU0Cn9jRQMY5JKz6kmcASKcvOlOTlPCFZW9z5vE3Dbc8m+AOfLUqBN7g97dFQRbl5o7
UeozlNDj28D27F5zz85WzIB2UUwBiS8GHOE/QATULLJROtT7baK5b3Z5otNNlcQcVRLEzdj6k5dH
3+bcOSdLwSarM9J9dYlmvQagd9/+tje7QY4L9mQc+EEELY4r/vl3RyM7YwAYMw8/QUT9JOSrS1pa
fNzo+U7GaT7r0Fc4XaYKkV7GVTjXCjgEKFUvPVJqgVsKHp4bbz9EJsCs3KZ+bT98hTB7O+c3lNGL
1pbPtM5872eCKMHtF8HSLKFfoqLJJ1gpkMATiep6Mkb9Bt/xt3O4EBEIVL30dC2NDw7SR1fOHzrp
9Ne6EzSDcme6irhHwGvLNzPbyC1wbH6+HTNUf2lKxn/GJn4Tk4mDaUph+nL1tS7GuzZQ0Y6KZkQd
3v6UAePbZwpXbqFlMyffCG5tNu4EdVmpZrzmHL2FTw+QNGuTLPi82XP7zTuW/EBMoqGBmGywG4r1
FPaeqEUaR6oyITmQJ9b+YGYYdyZIL+7PCui81wBijWQXfgGE21DOgShoTxkhLHRGq8O6NdCxnKbz
ncbv+UBkuqWlKh4lZiotzZ3CgS6i2YPkS1M2Ol4i69wn2Kd6Db2gVUyEyi+//lR0LubBVUou5vMU
cahDsMoiIh4aUqwRgQJhmGtSSmnuB7752zngAYyYt0FytCpmc+El+UmBloTgRwYwJmwGf0sPEj5K
XoXwlqPRW+5zez0SyL6wSjKLnd+bHbs1Oxssl6KcaCbkK8i6sP8x9p4zUHi50CjSBwvZ630cAN5J
+uw09eUB0HHoiJieloTw1uTUJQRniFBvLzEL1v3n49pDXHcjo7ACy7p+GkeYQHWNmDpS+fIliRLl
0+OzDWmalsOokhL3IqZnHEregRcLEU+GtuV2wMbPJs8NN+lbWS4NuNbsRc34pWwVY67vL6lNT8Z0
PEbW0zgJCOgY0BcSRt7TCiFCVCfuxIPnDatnJqKBnWGl7GyEC+Jign/q/fPbZFt6/Owh9vOQpGlQ
XtQRndQnqWrKRzT+801RJAk06cDKaCRDqjtdjTS+iaRNSGkynlSYs2bNu6s0TNnH1y0RSa/REOWd
ahDxFAnpSruFucvJdJLKuDLjvJQZyDeaak9LvAyTleQV/z5hzvwKwdbZ/crU+WT5x3f5Epn154yp
DaAHV1uWP1WCxlfEiJ2+i3tfRcy+X7JCQy7CabFI9DLfsVBz9wB7J3QgjvwFbXlR6xVC3cPvJMW2
Qv+byRsxzWQCgdbD/aCt71kStrvJLNGil6KEvaJwhPDmMWGX2OIfyHGDfJtONzeDYSanjf1+qvgN
D3ItSwnDhw7aOGZL6uXB2M71n/WNKMT+iP698itJO8PFO+pyDrRnyFD2EL/7SEIRbcQpLrjnVuJD
Dw+UKwidowjLtvq5VYRGnJxBsCOt3hupNd9scTOnrQxIBeOuEW8mmdKwclcpfqGUC39Y5FkGoRjD
jLD6V6BtA3qZuDX6HOQWWt6RKfdCBzwQIM/FMdkrHHvnwDu+U0ijgVubCtMlShjLqzUB+DpwOk+E
A7/AA+p+0hXLX4CCOPSipSRBNpGx2FEA8JFbD8SZINd1usT45/H52ImnU5vzejwgtkHNXYTdE0+S
rmgM0eCj8YXy6TmTHO23qIZrIaqM89gQh8A0x9d46jjpGOXI/4oePpxsp90J+U3AlxDURabZLnMW
xgE2ObTvlY5VMaq+iT/USh9o+dIUvwDdcb7WHV44QDH79ostHVnuJsvKsvD48SArKC4suQue/uIg
/I78F1dPq10aAWfOGw1XW1SLuQQfQXM8EgxLo8zNRwvMCmFMZSfQYQl4P5dnFEQsqbXQ2scr7xA8
pH0KRsURtJf055d5YUl1uTlNy9aHqrIomPC6dg4EdwN1gNU7Dkina9NZpY5/imN1E2JW5upIThzS
YoXesLjOet1UZsKrh9v4HLTRJ5p4MDfL2QBknjcAgfgqC4JEzuGe7NaBsihiex5RaZ5zkHJ11CkM
NzhPcIIGnMhCk77nlsqhzPAFsiLd3DrVCTLMv8HfB1ZkQDv4uRLrNcwXWlq3uFeDi3IEVQb+cagN
TOS03HfqOtDsOXc4oC8ysAgrgCjBsV2DYiSEFO1TwhHbHedXURERbo2AjCWDEOkgithNd2MGeckm
8yG9EyDYIsbyd4NIA4dmC/lrFnZOekgHbgUHXtLoxAabmGKOW1nFU0rhWz6yi2MeT63CObydYTwO
+nO8iE5dnmin7KVxMKZISOLfiKyyrEurK1lfzom6TX9tWBcaAm/kzaRYDcW2/dp9YORDGLtmr/Ws
LPJc9LUd9b615xVirXQ+bLU1XggzmGT2RBEmdHqW4sAHWQumYfZmnmbP9pIA4YyDmGIV+Ohfum5D
XJmgPjFqwDOE/mDDX9XHLhwRKzeYztZNmUGs6srxgcGuRSJIre2AviVZ2RJhviNSBIBFiMl729iM
oc2LI+/v2epIsdRzaYNdmj7rg5gNnRO9FEIwcWp0LCRwe5xRb3xjzAwgfazO8xWgl/ubPAkkyISg
ejpkMpxjDnJC4Pkj9DbU/vTT7sEP7kq+Ikh4JpwtxnJg4WPduxqa+vAWQZbBephZv2hyaDeHQfh0
kRwCw0DtyKXymGshTAmLBB3Qscn8Hrw8Ba3HXyMwdWyFcgvp7vUZtQfx6jl4PckfgL+ZbMEHws9U
9Ow2CIGh9Gcp4WvQMwiFKLiB+LA32RXCQDylr/fzLLK9fxCgke4gDeAoE9DGlocIor/4H792Vw4C
EsSSFFLOtmuxPMceQm3WoDCmEUFsoF7Kc0MbFZW2o0/A8Q3li7GDbT+7w3KQvocKHfDDIf89qRoA
fdtvMS1W2MwEF7NfKaZQ8zaxRn2hUOju12GsBt7GEqWe2UiT11R5RIY7z7xrvbs96c6U5ln285BQ
kA0cnIKoYHlaUnG2fcsdmwOmsbqMm53i42oMNWT7pv4pBEhFFMAGzDEcUu3AYPfWQ1FGPj8j7Z2t
WT8jyzS7edk4IFxThDUyKtk7dBhM9V6xqNu05Rfx9lgCvzdaJuWuPv/PQerv5q92pW8zZMd3H7iW
BcWlRGUtT7e3y8l76UXMtiGv4XBlHnSQ5yTDgFjpbG3ys8Qi61BpXpbqsaLR3SRBP2unxnKwH33g
SQe7TfVJyjwXQV4DmdqD03Pwp8Oh13RjcWbhsJ1yeu/ykPe/UueFvuu8lCFKCkMhCs0otJ0yCUqN
lDRxDsysvqutJCD+jok/Mgohqvf5zetkdl0DQ4Hzim5fmeJjOkj3gGAHtcqCJtw3cjBuGZVK4yWg
YMSh5sYpHY/4lt5CPmxRIsJrLcU/2+q/QkGFIjGt/6T95J45Pxt4CmtpkTM5fdwYyYjjA76UUbNa
qHsaAaE88heWoZbO9V7hYTh81csbb/hp80oUt9y3UXaoYtd2Fx+xwyGSuixoUyYULjf1ZPoAmWnN
ufUPuFo8I+l+JMeQMVpIWt1/V8GsuP3jTJ1380mUBJcpCMGqbrj3B2gyYmVkN4RsWuZ2HMNA0ZFH
8dtpsSeifF+kdqRGQlzW5GK066z41IDIXDS5nGxvjmgB6etmQJG9rS3XovWzD3hH2xUtiTECZVrE
2KSK2T0wqw2p0UV3UFSUeHJDEF/VdwRlViydB+76Bo7C9PExkJ95WBXy5fRwnVOrHwOZSNGgQxHK
j4oG3mb7GcGpPcJjvVl7qhAvyCDj19Fj/FeW7Ld4/5EKLQPi0eafjkbxU+Q/Fve9KQyRRYQ2S4Ik
CDltNHjTkkkKHlFsSmhyy4JdHtZl5MXf0GfKh80HP5dT/yPWsKBQ5sudfnXcm2+J3LYwCjxdkSRY
/HfRNtgB5fvMSet+tgCATYh+QkTbQ13sBwIoUosIkdEcOa8XZ7bUjWB3Oom/rZJ8V0GZ/FZbb2nK
KLT1ecxY/y5UEBHZFBSHzpeQMz7iuw0QUHQNjzYYt3kpyRjSNuvEOvwmq7Bfze0x0osAXV2qDc4t
0w0yWVi7B/9uyOck7jQRwDqmAAejLVl9D0DidzdLO+VMnv2tEMQyCAaVscNIRJlDxdW/TiLMnwFQ
WXPNjXyow3YFPURNrjGiistXFjt0I6L1aeR3v93qZIhNpF2eZEpBommrfjR5v1E7dQ1BWzLLSQM+
QlxL/4Mm46el9DlNjW5WkD6PoytHAhKIfWL7IVN5sPgOlJTsZjCLFqxNhATfbSw3CsyoYAXBVg8n
Pg8MjlXNTIx7MGJO6S+8wxXJ72Jg4I0h0i1zxNOHIC/ABQdGuObMdlXzCZPk1QnIJfnYh8JQvTj5
R1fwhOnN8pAspTDJE7sZSVQvosLWWNsvMdFuBx9k17Cyk8K8iobTSDC4lA4KadD3MUHbsX1Moo40
cTTV9aBnxSFZH2yIb/fM/Mnpr1ChzT0FKDhzTnW3BRoCRiCrMfAM3RLxRsHrT7JVyeg49KD2JH8x
tyZnq05J6F8oARdDZEgSvEAsSTVUxAgZsIckectCdgEJKCsHduoOh9BEVciB4FpofuCgwIpKMsT6
HclN5lELp7baAT3MqoZoNJFKAyudjs4u3muslRu32B3OR04GbiwQSwHiiuYm/dYJdAGQvjCTHxnf
pA8TrjfwOrNK8SzaaAhhuk56qXK9HMggxninRJJTHLIciPP56Xenxceclb3p8jHn85BRhe5x8Qz3
BRkGcvwj9OdfsmDGbdKjJlPkXxIEtfX1n5IeiBTNdmGm+nLhpb9wDCmNhHETpGk7qX8XVvXWefeo
ln+agf/PShnqqYwh2Lq9vB2SQeGFFAPjd++JzziPljITqYpjBdS2m6RXC3DFiCuf27X9SHT7Qmxw
iOUsdv/Z7tZtdv15vTPYef+rC58vBGLE+/MwfSfHvgrh2xyrachU9j7YNa/U7fyd/pIiIRQar/5s
DEDalnBCKR94iy81WXNjeAlIyQBa0Mdc1+aZUgHftCHX9U0l+cZ49p7IjLwJPvetB/BYmU9f6qM3
tyYDX1mfHKtBzQUWaY3Q+yus6NRbayE2QUYh1h20NSljXmXSZnB6JpJNI3nTGTbZS3jD0RWCPEdj
KZ4envvysnHqx9Cj8/GmzxmjewEa5w1O2zsv4TQXRQxtwDwCVWy4pS7r3ihOdz//Hxotq73qSGAI
WOf+DklS6y26nWUgKmY+gT/6HX2LmIfBPTIGSqqQ/1zF2lbeoX0RWgj3NLb1jMVU4bp4RBrDwKvG
bF03hYKO10XEc0vdvhHPcAgvyv+Z82djqpwlCU1v1VEVQC6wI7LVeTM1DsMzG/byIIzA8qHpGJ1E
2Ngm2hrztHPz1WexeXPRgFKgXVddCmdO36AsnqiGLLmELZBQTqZUV8s8We3h+BTqGu9EmoCOwkNY
n0BYrH/Z4NRK7JjE1LG8Pm6reWzW9IOh7A5B79Qb8XLhpm1D4/+eyIPHVnThRrp7njJAQL+IjUdZ
Hi+ei5PA1wS0ppMbvzWKqBTPMxufS3Ydl1Lmw0/73UfkmEkOf8nmrPW3atw3iUrr2DKjTgO7qCJa
ZS4m2ToN1IQkW4LuNn5pD7eTbHOQKfNbhbYeMe3v7Wl+8dRnP28s1Gsh14rikXPClp2htvW3mcIK
5GjlUnPtvvTr8vOR1x97dGfFJUdGKkscX2DsonX9fMDMn9vGQA/gvgF0I5yeEsFmU8juZvsyFlBh
mw7b7oEyPCZd4fLouQvN15TkLSnHPJ9S+nk3dZJUdgqTOCIL273KJNMJRjKLUiiMZfWsCu9HjSDx
uPvn5pC6BrORUUs7wnNtC8aX8tPFuy2yNK8v66uSa/XtJGeNLUblmmWk8A9R6EW7UIJsc9zDsTpV
4OViE0QBw5dwo5wthAd0WnrDNkEjhiSzA6B0Of9B4w165Oa9yZmTz92c/6ssykMQHRX21VSYrCub
kD9dz/+5sXluB43pr2+uhF1k1il7ZoqX8x6yJnVNRHPNghyFoxpKtmgyNUvBq1egtDjyhTyLZWZz
tkGmcxPr1/ETdR4svft8j5ZroPE0lMuzHVtbMq1HIdH5PfEYYaymEaOfxpqVLxnPw/0L15+ZUZIP
asBNhL9m8GgKGZqe4O1QnqcjV8a8pw3tOLtqjZBLXmjBjtklt2LuIY70bpRpmAAKO2IFf7oG26DL
G3Uxoh1qo6rzZygzWT639pKe38cT1HTAg+vtH78SCRQxjVCz3SSFQ/STPERz091EXiHV/7B5rLfh
Yajhp1Nx2h8bmRmJqxjoo30HcTIFAQqZBMiiKI/Wihq1IvZMFSVH5TvUQaWyFAJuM76K/ZQJYge4
ql0IdYTGMpkjk+dc85Wv+u9W/osBFkNZxGIR1bTqUl6CM6UmJCWB2FHQbtdJzh0cfrWvUPv7k1uo
w0jWZSQN2hcBqRHDVnEFvXsxYVg9mNFbN++rMfXZbO3FX8NUzxEUA8f+mZl02eXbJDmkG/ie7lv8
4sO3B/eMdjyOT/ASJQ+rsvwTf/XAiuXfVMYdWY5uFBRgZKQwz7ooqj8Yp1/+JdEyKQ7zIecJCEsO
Mz9glb2SglN1PtRN/IxO2IslmNBrVjH8vs1uEgxuLHnWVMwWV1F/yUWovQlkmhl0DDPJiqkBwtVD
abVvuyJ8/u8lNdDEmX1NguhIKCzG3SXDEcsXs0JfionuE9h4bAIq6V0gwc8jK1NpOVmZ6bNYOajt
byngv65iI5XzOuOLRHGxT5n4jndPMNk5RZ6UIViHbq/+a1Yyvome56QeG7HAOTp9fkCG+/yzgjWs
wzPhwkcPwt5YfEv5VukkL3sEa/CtrfAUQjXaySvZergRNiNl622dsAWXE1O6asvx4RqTQVQ7ykiv
mbunwzs1uNbjLcM2fmGwVcWDa9jzK/3ux8vNdQQlkL37UvEFELD6P+KTMx/FAe4waS5e+hp9s5JW
3UR1H57kCSrSWGJjTxDSdbfBB6Zg/G61LO6TQOOTQOhi0HQe3VAquefKaR/9Xpg+Ozmx7bi1eTpC
j6MfieHEfx9nfUnq/Xlt3UppeQD5ZdBzTXEEYG5PDTosBuIhtIGVoKAUle8B6BZ8j3vZUHz99Feo
c3Yl1JqMGCWRGYMne78/gLt1+gFGQKEQXH1boZkeMnGonsmp+QtV34pfLNclUnsQQpKNoElhx8MX
3ug9ryUY9RcJHqX9/yi/nCWOtLN8kbUqAQL7VAwXpHdSRhsSgYFyO9BN34dIVVdnojyqTO84MOBM
6DMx79Mn4lCsxmOJ1BpYXvPvSs8ebJTFGbmaAHx+hMXHNLT/OCuU/zk6TKgFhmWftpyyjiJMKZ8F
e94OhESgXQ0fVPx5Sx7GQjnfYne17Eha43fFh9qAuswdHKC9mMH2ObvvZ4jelJsajTMu2O8hyqwd
qS8yYeiF2TbVIICDCVfWRcH5AGRhhq6aa4sacy/qrq76fR+1AJGc7nMFAU/WvpDzSpeQBnPt5v2Y
FHeRjT4yIvXrYKU7mzduynpRIKWc+J8buZbU8i93vyIzmnYYAMaN6HqmzwovJ4QRfXUBqRCNuzjR
byavx9OQcqCY1g/5DROwzCFmkXytw09wBmIjWk5EqBonS68o7RriZzDGPs6tpeiOO3fyltHdvkWY
CLwoB54Q3fcJRvUlfcWAITAvr4s400e6iA9JPWXuu9INEAM3eCUIamSHJP5bKJKjHW/npi6D3mH2
gPkkDMdH4J0gag3YZ7Ra24JNIwQKhnu5O1qDxiATuNnMlxGdTCrNygqmSfFUmJxeRh3Q+Gq2Lepn
0t06hDJET5d5IZZ4yiDWTfdBC3pmxWg3XWNxoiuOoIV0AD+jI40PLV0wJi71aETMjuo0Y1muQZPU
03yLVlzDWfM434/jXAXu5qq+ND2y1WE/TVe7ox9zxc8Vz4+iH0Hlgw/uNAgiJqEh857emYtQx6d4
m0jCNAvGWaW38mKPL941OFbAX6xDBdYjuEEKUJNwE07bUemj+cAmXwSO47wBMC028zqwQHGvklcQ
0QuRmvbGoe7qOOSADYRWTCASegz4lLqWidZ0C1vepT6hsM/N79rNeNh2tCvfJN0921/lcRJKNkZj
Ou6C+CwtRkdZ6459krptoBDzdgJ1EZ/9GgRikSBbdW8vV1f6HVnFwled3rg4Qxzq9gZ6Oz93CsR+
A0YNAZV7UWW0zHYPiRKJGitCRcjGx1ObXyT9SNCLeiOFZMl2DG5e9N6h/ac3pseiRKbqF2QTBtr0
89fM90as8Ax2P0Wnvci2HQAFlWi3wY7NpTEM75c8dHT+0cRJ0FXz5ZsLOICBa2dn0DEg4SGWRLBa
lUZU7+yO5js6NQ9qlHdC/JIA3ZyGjzdJI+XkrQSLfT1qCuKdKWu3ujDteVwKWnOHfFRXqm4BxQv7
KeGryV/Ap1/TxxqqYJ9n8kvibotpyWHLLSO4UsHopcf4BNGPgLBi8iSm7S6SU7K0ziPqdB3St81j
i3p1SFpqEhc2gmaimG+KBY6XJllCVy6bLzt8pwTPb5P7paEVURXmvIBrOWr4kL/xLH+WBp2eI5aw
ft1io0fUI22vnzSkphu/92W/YcypyGoZ+4No5wu/+mWKlrw8BF37o8fYLHGgswx4jSMbjg6CeMBp
XH0ObuOXEBePCIR0cJRGeGacM9X4JbGtd6/0uhKMT11NxRVnJ87MphAzmchese24FjQRckXIWznb
oBxujmjNF/BpDMK2NheAGNxUI6J9RxwzL3N3uNeUkDbM+MH2lPOfcgJ5scpNO4qoEkD7gytC2wFR
e5doXgTj8RrxA+EgSl9JyCo+onLrPTPRVJx0kT6cTrFx/q+avSluAavcUoaJ+Om8V9GDl9TI0mYr
oXie1f+hX2oZncqQaDnIqi5En7WgphADhUw/cBj1jgAe4dHqM7mnMWE5Dl/ICBJSN9k5aDtoGnIN
u+2X7dIpm2LcJhixx2hbIPh/7ivDYy6mzJ+YL4GKGu4Ut8IfbRWOmcMl3H+gjgQFfAaYWd3P0u2a
nsf48mKfTZIoCCwVnOTVh9u/iiK4nUsM/nbG8Q7KQtjrwxNSmjev41s3i/rh1aJjkZxUEJqvicAK
Xc+96GvZncyK9L4rusrfDI9UuKAaA0KZc0xIntX32ddJ9UAXkxayIwb3jeBV/UPyk4HJrx0C+QHx
4biK/6F/MeCOCYJY0RHwUyF/QgJXo2DLAxzqrlxIIqh9aLmbjEm2jtUitDkjDOjt80gkFpKNwKdH
kIZCjXnee2HhtS/gbFNUjAkoSv39lKIViHYSwb/031ZSbgNbKMSs/u5v9sxL1boG1ePTW0ywc2dJ
jxd2tsD//5uOWTs4oFQQl2jfBEYvNgbS4V/RqWfqx5YchFtfk7lGuW8uR1l32eheMIaJE+IC/pkf
VvliJkCXBaPFJ7xNNAdqId7ElmkVvtgWr82Fw6f7Cp7IQIkH7UazdYQjEoeqC6RirXW7hPnmnavf
WSwI5waDiTfuBqXjh8+TwarFQrPDMijTYJmf3KGL/bxbqm3GqjNsyG0W7/fbat+sWunq03NES/M2
YHMIl8VMpzb0CC5nHEOjqg/p1lpmIAb0RTKSwpPIotygjuHXPYhJuo97OaSmkqHh0zqxP4WjXxCJ
pEm2mYuehp2OhV61e8eb1YXUmi1Q0CuI96EGUVMJ8wsH5bwlLa7CoppX/vWGV4WbKZUmm6uMscwb
3lSfozsbHqsFAutjDnyW3uytnDQK3sdLAeca7mVWgiwJv4F/awfKQlze0rexXPFf8D7updEnia+J
Iv0poTCcm4CBcqifWut8codchIRdvgaV0zLBu32l32GpTp2Zs+qFdxXgtdbS9QqIZBC/HLBaktIt
UM1tz8j615VB36Z1mod2pBXnpKTDaAXNe7dE+2hMr+rGS1VJPKtL5aINcBDlZRP5LNsXaE/3TMq5
Q5pxbolmWyXB77jw5JAoDbfNssDpeg3pyEJ+aE69fC7UPtE2LWRbSomD+I0QgbZORhBfCVTYiwM+
rde8L77tAqGklund/Dv+GMCs11PAkICRsa8Likn+1zalfUE8tBslrUGqyBXNMLIe5YcWWS/HDOiZ
ksQupPqsCmnR2w3iOQZ414n+X9xRzPcQOifJB8x+rstpEI/khl78lU7JK0wItvdVCDvOPQzWbnsC
fi4T5x9KR/BdhclKx769D0BQOdOViAcBilEXfR8jp+UJklAR1bjP4ufusMfTKn+MD30o4Mny4+Ik
syvsdFYdbEMT47xYrvCJwqMnbnXoNVPbDW2XuUql5FIGWS35qOYl/OK5AYkbrY7ZTDG9UtQzjNNe
9GuPg8dU6FNWBtFAh08RESE1/ZUuilE8lQy8KXlpYwL0qpv8jSRAOJI6i9jcA9quOZt9F6qHA1PT
4qhx9wIHT99IzcNnh8boI5zIysPmwkLjstqJfFNMPnFVSGHmurtiQq2Dnb7nBllZvmg6VuUtJA6n
uAzdU9Zf29J/nXH4bxxfzUABbyo7HDcmJTtY9xyyxkwhNsVMRpsYnlCRaiJHcj4DZRV2chYBFg3v
sue8QFqLelU9iks27Azmm27xOtgoUadIBhrL/nOhIdWEatr+lVygsxp8wNW867ArbbaEy+vq9tt5
YtTb1MNA6VcpjBvIsh9zrDN86ru8wG8tK+TaULNjR5NTAEy0rFq/3HW8HS76fO8VHO9vQaXHn87p
7QQW5SDqOrxFflOkmMVgL1otWxuN3MVYyQk3XE9CROQX0Gcuv6T6q5G3YcttOJY5oa25qZNwS0t5
kd6SVUdZAvLiGHe7mOhcWni5fTqYPnipXmKZNzdoNrS1FgVRP5Z7t0P0KNEb0yhvvBxQ/oSZgjVR
2xAL3RnvGduQJQG1wGNjaHaoBgVr+MRNTtw2QoAGwGtnXD6FJ2KBjKo9621rnTQDI+vi80SiTAm1
WgV0lTkvkvLaMle8Jrpi3NBnhZOCtEAsHa+xtlGLRGMvRy4TaU5FSYS8193N++Fbg3o2TaOr6LTU
HUyODWgn2x6fkr9q/R2VngX+qfobEyVo97bbY/fU4lhqNNhfVAUF1/VeAEvC7NDY8SIkPzu+gTXl
wVIaV2YbuJWstUipTPOFAeSIH+V4YOfE2cNaO+Ahrzyz2Jm9N9koT8Lp0IlNKq7kkkWaTMNiIhDD
62qele+AdmXj9kNgmqlbzqEwl/GNGTWVy91d0+ureHNJ4MTf4Nd8duB7JPlk1eycj8qqLPM4XNtV
CsKjGBnvfV+2j47KXJgeFkqvdZ8jUq1wM8B9xmjR6tasGj4NH2ev6CD+rskN1A3mVpjfuAUfxl1v
lZm+leJEg1e2K0bEhPeocfWnPX3zuLZWakp4ukyGNBCCHpSmwgf+vjA9S+Cy8o0BdFvBzRVYgbAh
y8u2upgCSQHDb1VRn66Qv38QEwK0oQnssqo89n9Tts2aSaQBH8wBQ2KzHw6UeFA/n/gb33nTuH6A
Wm6iN6LmWeSemR/fKEGxlwiBCbVtJXvSRAnh8cqU2jxMVaE1Jl0vl4WD1PDhylpV/+AOYWYSLbQP
v2rAB9bWEZ2Y1OZiUuHM/3ljVWvXAEKMqLuWB3J9xBuRfx5RsDC0SIYsmpGC6UVtitkDhQhaRirB
ecBoVEOtnHtLtBxxcmIqgpktPsj+pgsHyuY7GosUyJPI7oMcnXkt7vQE6w7REaaoY+jsUoWl3MMX
RNWkUGfZ7E6x/Cgsix7xHX1jg7Gc+mIHb4A+sp0ksn7rTraZJbrtHu+n2D3LUytBuSx81ygu3lwh
/mNVfMbG9XBxv2cqm5TBIJLAmdKmodRPiN00C8kQtT4OnQQDbiBv767X/OHSGbqOPn3ppvTj5hs6
2D4liYbQn8e2ls7yv5xFWTrraju5gOH430hgnFN3lNFXCteeG2CLQdDp4TbIxriA0RMblxciQS9S
wqUcEzcI3njVZywnq3u59KuGxSkoeTH9sgs4cX1kYYRV+d/hQNKayVnXEFEfPLRqkOtBpSDTpZo1
LHjoC+eQRkHex5uBcfLJNLa38Fn2M84ahlRUKTbqXKkvfhmKa5obFOS0qw75Pfn3YojrXWQLAxW4
KT6wGMzYik7+e2hMegnjKjNAkeZ715rjO5fb1wM6MqdvUt+f5MiEnPU0yRYLkQvu4/ThCr5OMTk2
BjWmKbroj5oc4OsZHvSfSbRgk2eqnKnYvIUrk5GA16J0iUba0sJyWGtx7ZJWrSdHCHKLp7BgQfq3
fs5y1WF7a+HhxsSDMLLg7f6kockJpTHGe9E2nvxPxSCRbP1KdgPEzV9QtBuJJ5dIY9QTHbOWjdzm
sAxBZMuDZBcYTuWW5Phv/4Z8w1emfVMbbfU3XYufXeIj7vRjfNykcUsDh2KGYqQA8WJe6geJOvdU
nOXi2jaiNApNbNCWaXXw8hjKUHamCJXJstjvWoJmZja5n2MAkKx5UDhE82nRwK2QpQ2+6tRc4Y4d
dZy4bZi7hKkNnkN8Yg8+cuwERcxgLVKCwUQMJRZtFvkn9Q7rrsCVgCURv7bByzS2cOArqSXJ8P05
eotenSiKWMwTwEaHV5CbxX5TPbGTxE+eQHe4MpptYIR0zDvlnlebsNj5xTfk71auq29nW+Y3jHAN
wFno1KJMZ5Nb3SlhFw+C0mJvFf6eZ7PK8e54RT6v6waFvcD1xOo/8XK5f0J/VBkpeF0XnWZtzX2r
IPDZXahkIuwYBxTqESTvBMr/Ru8QUe3s8SenAyYACAwwI/jL3tYEUqjLQwnZMNZCMfESlQUbIJfp
slYGK6bKu/+qZ5kC65fJPu/YtbuQlOVR4I4sPooEPae7Hl6codkzUda9nPzXZRmryGRsP91ti+mQ
lGE5fK52OSPLkpBHHiFNZCkBJcP8n1iKGk8Qd0lSW9E0xodxgfKGKmYptEuJ2sFD+LqZKCMRSyUb
AKqhBf3CnmqATQ1d8jQIoIXFvOQr91SVIy3m34ZnLKVLw5pNtAD1pqvNxspzFxteuxKB8DwaWHGM
IcUeI9Z+dbaZ274W2Qm3IZ6fKo6kGeTBFMe3rvvkpLXw5y/0yRa2+1Vmjzjaozl+rG0pyGoB3UB6
6x7L91xdmMbI163a8o5rUea//oBrrWAFMJRXs3PyoNJ/VzDbVUrNDGfl4lqtMnNMnxFf+QScLXFm
t0JLPaRGPAb60WkDTlWVqHiBuWxIreB5L17rSXm6AGk2hwvJoyuTq5pura5oXF5/mLfEtkEAvQag
SZSOnUqKvSfRnHq6vX6JKu79m3APL2V0Isp8ck1mX6460Wcau1D8co4xHY5sbCkFebpJFDybnYZM
iwHX2NpCW9DcAwDRiEH1AWQlwkLWmzL5JPOcIepppb/bRox1XOc7f2kzlziMl43oCpuiEIUCcPN2
H6nbT2MQw3RuQx1M/bRLxVNMnCN+aEQjTk9DgNAiVJDJGbGmje+McXq8JKB8VB9jzbqojf5kqDad
vZMmM0uvqwdUXvEoUbqf3cdEgxLLyjk6wHhQ2aZuerG3tBM2jUh28Ju00f63HlVKn6+s6WwbqD+c
iQRugM70tdS6VhGxzo8MJGj00Eg8NZ17ZfHZ1aOkAQY8h+PzlWG74gYkKtVMuJzHIAowSXxvnl/c
0UpM9UUgu6c8vC/utjOg9XtMfFO+fVfpEdFPlRMMEup+vY9i6SwaLGK43sLAAlbxPKGLw+xV1Cov
ONur+O1YN8Ljs6YyewTXmQKgcNZkk3BMcDAMRDODhbf+1PUf0CjInyNqhkQG853HHfP4aZ0htRyS
JFY6wC4VNxmpho7AXtkjSno15OwblDZjpLH4i7J0/bauslETz39581WMe17yDjopgijh6jpJHLQk
RehD2BXi2KsBYZxS0f2063v9h59hd4os0AKyDECdT1SAax/MsOLSIx0Lr4nzIOnpj9uLqFpkdcw6
sx2IWQJ23MmgoSQVr++mjbb8NWQ+yH0ZANPSfaO/Kg/d4eMf9sgROZfFIU3powNsDT/63RvXz2V3
m1i7sNp3H/wxeS5j9qjQzN3A5Ri3MubyOWQE2mnQhtdW8otdJfyDa/qZNRNMp4rbvv+T+BzBbr7t
jH4oVT090IbId/nIdJpji54EtIKMCGT9nwl1+NTM2Gmi9r5IlqsTvFtqpv4Zee1E8HDD6KH6IHqk
lGtbLyaPdCj+EvpyncIn+A8yQBpOiYgf7WvyD4MUxaFtrmdcnMeKK+Q8wSWjs5ZRthowcQLKXvkf
ci3Cl8HFPONa4WQkGxwTaa0c7Kk7g1qF6cFkAqtB0E+yzSSVs+phaZBuw9JXXEP8FUpm7bvW+Kuc
7bISPG9PlMOyWcQaw2KvcrzvmnwzW4uWtZIBIUDFraXTRYAZBNF55nd5MQUxjdK2XYIeuKsREYNV
D5vK/pku4RPqc23Vi0+F8YNXlfZN6cb1p1h0rt58crj1B2pIdiycbnO60IXXL9OzN7FHUlhdh+kL
0z1Ju/j+9wRjY5+qrRQYPuc2f95NBCVvxg66VsSICzzIi6rQldsPHK9ss5QtDnZRKVuP4HxRX027
1NBfqKy3zLoZ7u7aCXe5N1WCz1bz4g+ACtMUM9K7AfYO/6263Ou2yAtgmKpNokuZ8yDVEzW6Xp/2
LS9skiV5i0ojfUdoNW/7lhOGZyyfd8eLz+Y79miy3tC195YQfCHbObNrRrDSF1JDvOLhJlhmMO9a
+94uFTIzUQL8I+ke8oK79TcvHR64PHF3TKa/BCx5m5YS6rN8epj5vPVX/0ZDvET9sFvPyoqMrP9A
4S+T6AAt9kYGr4nojTc3YFLuL9kuqTUXNgJJNiomxhpnMFBdXBffnQHX811MIJ83XKIfGwP45gDu
wk5jREWGeOgnFs0UHfJZCqmxnJjEyavMpDvD7tX652NgWsmefyBanvKPufVQuTV7p9qGucPO5pD1
u3FErEV+eIqU52QdLtXYEFY/rQYGn0LYqA3968on8mZi12aUKOXhQIXbEEF5Jj0G+X+s88IbVJGL
rhn3k/KrsLuD1hmf9o2S1JaOUl48Li04QpUbugfo6Ll0Z9PPj4pzvSnAybQgwrNwwM8hQyWQGMHJ
zunTcQ41+ODiq24gDYJZPI/0Tprs+g1eSTdOXqZ1zWwrIG5n5mlbJpGq3hZZ+wBJTGTJytIpXq1I
lMgb1QBp+7HgVJUsVm6n0hILEtePlfbqtaRmrZJ/a/VzX/NWtO9mzWi1zCpwRV28Wc/LTiR9CwY1
tKkbrjea2NCkDQAsiMfySyZKbaynq95I2GYgjNq+KsgDDtf0SGBfy4GXuimLe6tS6v2t0HKimpWV
meLmx6yDj8E5nv79xrfscCjkVKBpzjYrnBvDLhUwRF9eAuDSvaOm+Ng/Ij7wgiHn4inBd3obPrjO
dRjmENuDcna78I78H/jqdKYG0Djh5vVHWa4713NRfAIqNTMslwPcD121BWKEuZc69IOaRlRbBrhb
y3erye6HCJkrA/qD/BiF8tkzDV5VlhMziO7BkPLgLW2ybIqPTfgsCPdjCvbCTtbxMHUa3HdZsZ75
8ME6xcLdYxFESvXGF3wj1brGAbkuTd8Tb/UhZht8JebDsagBdTp2/DqmW/ygxFOO5WjETIe6Q6I2
IMhCcfTl51+1Pzrp24UnjDy4kZU1o994hNM2UVSyw+ZtVO8oWndT4cH8J6EHh63AvwB1KY0aFFXB
EwjKGho4RLEertvJg9CYGpTEd5Xt0kwVGYn08U5vj+NY41ib0gxL3UDAj0zpFD+Ryfy3M1JB+wI6
zqRILoKVYoRcXDXIxVGez4dPcBDuyrik4V/gH1+KPbIslBXvmbUaYiJDZKPM6t82EcOLfA2EmEkI
H9MPp56xcavekCIKiVQ4RDIlkt8FeUtVThJ9Qa/wmIsTPugLo/+uQPOvhUSXDYEXpb+2OTUzdPsX
4OTcdaH1ekXd6XoFUGFC7kQ3REjuOdzIP0LKJ1oi8FHK27YumZwBODNUELtcCfStTCZApcu0Ee7F
KJ/OVqhFxIGtjq4gG7LKFKcPtverKYZn3SprJeJM6EUGg49pIo2yr1/SOgTwyIwXJYJz7V5vBSmO
NXMbW+hAJbGQZYsWkqMAyXzxq+6p5bo9zAlP+G7c28uhy224gKPXjCM9o4I1OqKspM2t4yhMIyOl
GYPqcyh0Rjr9uteTsTVcsU4lUyul/SF1XZTjqi6mA3vNm3dfxoKd7uyI9msfdvGm64FLrIVbuVZ1
UGD7YIrik9HRBlmzbiKPBemJS8zLEOevIMuB8/ZD/meHb5GRumED21Knsmk4vg6Ez1ogm6h3tCF6
kOw0ZbirfpV2vOWnfL6z0r9qas5s5IqKzieB+WsaXrw2BTuQLtMzu1LR7+wfc7TNjVZBUKRJgUvk
z8/IAhy+D7YqAq3lMsswOFjqKBd88IwUHwzoBqFpOEZrdtRsNYNbDdnAZt0FeWZzJrodN7sMGKNE
ZxRRsQD3NYuNKwVGELN5+eWzalHd41KFHva6SjJVKyB5jV1S63rNdBAvsv56A+aA+76WMW7HS9H+
jlVgV1Zonr26r57zQPjOmGmCQt1Dtqk/DmTIvNF/LTcZq1uAP36vtKJO0Ju4PRzWN8Eq4zLCj3qo
4rv1zhnnPdbJ0JWgvoU1tV3mK9Hq6oyxK3oXWzQxEcOOINcCT3al+fRxIw+vS793m7cZCNASv0Lg
RFR22WUPb3jswFCVJH5XNHDPZX0NR9TNxhfnIecJOGjCD/FNh0epV0LzMIDEDUC38ykCsVOK0ZxO
KTu/SMykuNsVSuL/Ehr4glexznzIKqFI+5Ez2vqDSbQhzLkvkWerK7bDjubq3+U/2+czT6zdezsw
7xh0ocSDIu5o710a4HteHlq0z2jCS1V9HzNM+G9hRQ7MGhM5upNsKTjd8tJRbbT39wIU1F6EN8NK
PyoaOjuLYwIYWeSjaiUTN/CAQB0GuaYHIYpchUoGwobQ509Xx7LEpzDtwEV0NUZkp6br9ggnZ0V+
TeEWadQi3Fu1RIrHST9iLqWgzvJ3HIDuM+KUwhsQqr9/xxL4eizCHwr0++0t7sEyu9VodaCa3b1p
0kSO7EHp2EMoj5llEvZbZlgW9keNXRsXKOQyxvg2rpGCAchPXk7Wu1KTOl0+X4pQ9KDez90h+C91
aH8T9pqG/nnQ2Tm7MlnDvPts5SSY4ACgiOiJXJtAL10XqtDkcTpNyDonokWpqzT2EeSm60tJHQUI
pMPOTyNADkSTlQDDwUA++vKRVD0s9024X40nzXmqsLaYNdf4F6nsXA1SVuC32MJlSXP90pruWmXG
MQ3W6gpvr+jsVT9DO2FtcWi1Ru9uYtQNiyfqTiE3yNu8clWDBPVxJNH1NS7jPaxrP1pusJ5Z9qeb
1kQwW/9WVhrjQEkmOztr2zQbX38m+0vF84V5oYuAsXXBHTOSeMUjy6j9vZdqvdStpfV5mYy2I9Id
tJmnD7xP6Avoh/Jtk+3e90+/ZFH1VE4d4YdXqPwXA1lz/UPYu/FTpqZI2ghlys8X+K5ry9/vl+4D
gU8FQ6jqU+Nib80ZArB2OGEBSiQUEKgzDJUIP+0+mYiO/04Qq4OFa4paE1zoeVVCL5QF0HnsC5FV
FP/uuP1IrcEa9N13N5im/udSkKw125hnP0Znclla7a6OuxgeuPt2okmfFH1+dkM+EQdLMVNy68H8
UfgDanxCmRrsuFwfzjGuNWa/wHZlNSo6ERSdUosxXtOqP3LYA3AILAo5jyljjUncPZe7vcsluUf6
azwpigiQ0ywue2/1UvdA6ZRwrabuvVcR2rU7Bhh2avNJp2aIL0qkP1sbwlPRGKxacrMM/A4XHPGA
TXnsWMLTb43CZg3iNbh28ZT0vKQzvXmLrkrVEI2IQ/xVljRliOg5wpUEupY2/S9//1R/CCQUHOqA
r/Be/d+kc4H7HYbuVq7cK91jTSp0zg31JTWKBHygXRl8+L6HtPTvZ9Wv8VEp0sEZwCLVPMfeTd3f
Yx+xZgHpO0HV+Mvb2oKI0sd71kbmKhmEmethuccEOvQk7o91BDQ452u1wqhTBMFYiFKcQVAOBH9a
wUU8EsH4KQSeHCXyapvVysqSIuTTUfndO+YL98lNRu5MXN2Wh5KVVVxSxcaMUxFg56/mbqocO36B
ESuLrnq5bYzXExYEUlm1BzspRHYqFX5SCdj9Jgnvo3OfoVv3/rBq47SvvBJTSzdti/Bj2gE0ZWz0
/BwFSr4iTeqNuU+4Cp4V3dK2dSijeCKSO/lPxjZCYfcjLQ7AYh7ALoobcq0MNbDJjyxj5ApCaBmh
nBLI3gxqpM5fqaVDIO9d9LfNhrH6VY8BxfKhzpjWfBDLxtJ2XbPj4bB5XjEbkLplI6ObcQfBEQ4n
XKkExVQEUhq8z9L/xLHRaM7vDp6swXxkXxnqazebBOTLfLxwKSAUXX/lr18pbPlAQalUWoqXov8N
Urwku4MOOWOXlnDU0oEjG/16HX/NhNnIqLCwj5sPtIr2T8MpVyb5tXw+oiTBKYJrCEDyr/GS3ls/
oGjXDoiuU/qrtf5Q3X6t8NdFt3ASeGtQ+B7oU+RcXSmUrcMVyCFO5TJdQyJmIWzO2GTTg727KWkd
JekOWP32v6PB8yo2SGZIC2qF9/kHpEaUAkJzKTct7oBo07RSh3T9j/BWXnYsm8aEAx4L2vXdFjTx
A/6mjDJ8zGJ1QTuks/YZXokxnNzZihKaF+ycvXuPJKRcl8D6S5jeuiCllrwxAXk4INfaPtHGds+N
Aj9vXeR7vs6BcN9f7SN7ip//ivODj0RvUMaoVSvKP+L9nIttHsws3nfmS1mRUyd96EVuwwRcLgKc
0lVbm1GbvYJEjALm+2xxWx0JyPYzEIzl3NoIM6dRWZSYtfZtQUJiUMv+IM7A+l7ERbG12JfbTSxZ
P8U9ZD/LwluIv7kD3TgoYIS8Gfs2ZWok25djR6B06npB0aKmnN5wy4YL+kpuDNiSJSs7IBtXZ4KT
PwbkPS4ty+33Jlvy1AXjskI80DFlrGqWpXTqN/QypKtZU8OKie/S7LkneO0V7A+PQ3Bvmd10KMni
6xr+CyKYcbEtmLGZJXmyZVfybNxTT0p+6snmAE396pbBIt1vDDaaKAbVKww5pxWSiRgXglfjzyTc
01+k7IGDyh7xJdG+WORoVcyYsGJBsT4EpzWuQBDIs3E/PqUs/+hhhj/4OZws1kmsC5bslB2uFddF
CaYerp8L3UiEixsJn6nLq+i9gBpabOcRAu+zi2/oToSCI0jr9hkgU8fd78oNwR9c+hx8XJGXkZoF
PCLCFulBCdAQDfoSyRLHJNQnXHzzhYsYuPwswVBUbGZQQg347EMIVjJNeE7HjF+30Adhw2ejSRbK
ZJqjDVNGZaoz1WYTw3Ep9aZMJ9P37F7Xszimlhp5y4ZWTc4UEEI7u/I9XzukeTL69V0Gxe/N91yk
x6ZYSVC0ug4jYu2BRY5yddSRecbGUKje5PtoMqojviaHbX21nXw+Hh+rOdA6q86+Qn3BCDJSdlUg
/gjE/HnG8Glatdc+QOVQzOYw1v3PCXmD22J5KyAjsgIBrvOlMMkoU7U7ktzTEIXLyDH3jlxaLTnD
1lzey31c7H58iLWSkfZM+2EIsQ87lfXhXzjhxlzWz66eGp2Ks7Y8mbLCjgJRgjMm9Ji/fQyQ/aI+
c+2ZQNV9gY/+5P3/BLY2c0qw1VBQEdTgNQltidFzJmi/zZGgn2ss9tLOdlFn+9uMoEnLN7XusE3z
fm5kSIn27yRcLuZT6twB4otOOVOFgHsnBr4LwjdZxdp14EX7GrW21dgDMBONaaBvksjghz/w+fby
YzzkNd+vW7K75rS61etMkQMS9vFOBPDdMECD6dUn398h79DpaLXcTAjIKbsR4wXJjYFtjG3KwnGR
OH11TWdfuvWqfLNeBlCq7OkbRw4n4NsiSbAZSiMeFcPYzxTvvZT3BwpbtKm7h0oIJDhI7Lt+FAfP
2bxncWl4PO7idl2j7mvPv1wX5+5pBsOeD2fh74dSU2EtRXwSIM+dHELC8sqOFP8rw9OCRPQdCUym
SKWt2+Xm9qkyjW4RTpiDGo+8wUABLcxg/SkMivHysEFej6XmwqNS/pk0W0SWFfvzgg1qn5+Wn+Xi
tQON8T9SCxtee3PnffRRCl5j1JTXWuLHY5MMKq+PGrCKd9wcTRZSnS3eHrdqEKzPj54SPUYfkEsY
8BUhrJb2YdunqUBjuylg1hZW71gO+uwBhRwdB9uR+ouP55ur2KoT9Br+yaW4yHXYHhw9WsXdkWgz
KOLQxUyJBDh7AUIP1/atKnkuZYkOkjZmdQmA9tx0gaC+MrgsvpbBjq/l2Z65yeO98AjQk3o/Syg0
IKi8IRbf7L2WFX4+fLIyuxjmL5qGqm87wPHIP2bxy2yvMY2bCeKC0OrzFQgTnhbcXhc5FgJ3CrNj
ckSMa2rNSzP0ziudRIy9yJdciOjj3CdMrHNtaVsc+nNNIc5VZ0y+LkRsqzKYMryvWX+mqTPPeo1O
nTKyiWTnlAESHWxJWM7D3pClCNtSizLqEZCHFEcpJ+t+OuHJqHv4AcOkS55lHKC0KJopiq9w8XW+
RpG4UGVGJYUm/vEWC40m4UFbXqEckR3vHBIGnMh/U4ZHaRBbIQCl1X6tshu/Zl25YnzXbQeMzixP
IcYKTJhYBlwwPdyO77lmWzar1LG0foZV4Ff/kPB8aNbGUzpfk2KfDYyxoA9k1qfOKIkhXQH470DL
L9F+1h2eEjFy+CvNDidOlw+clQ05p8Okj5qG63qNQqJlQRHQ+Pc/cfxRBCjgjYwG2zNk33k7GtkU
tkvf1bBeCIRC1wO+1qkPyLIrq/ti6SUC6XKUdVyEdapqzH2+um+rp421BAOD/kOZz8XIFcm5vCh7
UAvWvZFRhDyoq01dNA0D0pSCa2soAT8CnZGrc9RP4OK/guqyOE/mMsKCRJIAXBQFsrr3lDTgdvpN
KNZ6ZVWMgDdIsLVQ+n9ntqeGZ5cnoSTCBZjKftvJsosga6U4/199QGGbOyDqTU9Ad7rVPDHjmTSI
S6cMSZcpd/BscXW6GyEkM5k0GRFUycB9eocqyWxgnRw49jDBE3PAFw/MhBMHu08p0DWIgorb9oA1
7hUByMtJ2S2UIzhQdRuJwXvkNWS9Fg3jvncj8c7+GviKk48RnL09pHBhNEUU4Epa+s1he6nnvlJ+
0cso8UH3IU9qPp7REyvnswao3cFUS7ymIBp/3BmVP4xJb1OKV/oV4EbDW/0CdHCjlq/BguMY1Zhz
DWt/3nDy3PmF2qqFJQ1B4CeVYqNPY8gsLwWRwY0n6IVj0ZCMQhy0k1cibVQSVFI4Wn+hmK+/eTqX
qwKkiqyicmBLPJzRWircT+HkQMP5BLNDqke/wgNQCDlYgWn5SkN7cytCQFxDYJBKkKXhu7mQiqF+
5wO7OvaPGZe/ky4cOdfALDbayGlpy1TaSk5I1AHgtgn27/3WAee30rQ49q7ME2i9fwua67kr2ANT
YXnDFFqmDFZ5d+Fg4bFQhYf3PrVFVVGs32ZrDc2hAnn9aboeofAv1AX5upgaX4aZb/Fd02jhQMZc
8BX+jMwUhHeYdizXtkGt6pYw4E/jrKybtCB7G06vnw3xaKh2WXtVZVFWfvze7evPaieQZHRxWnpA
DdryLHkvnr8yLzNnUUdpqUFwOzfqgisosR6xqrwZb5rKHnMh2g4HTRBpfNTRaZiI8YahG2stvWqX
SpktwseDP4alItkXosoF0YRp6DCN5Uzpx7o1xbdlhvLjnQQjefqaOeklGuy87+Vtd3hJTFqd0B3r
RD6jYWgcUOcIHuOCoJTddUXPBGOcrKTfmPCXUckhHQdCvHd3/11Vx38Rpq2tt4gAnGOJqAvn7H7S
ek6ocOqPjwoeCCePrrNVxeBv3g8HlkDeaaiqQzlCDHwbNgQtAs7zRMAvU3Cy0kfGNWmXDmQNJdVM
j2Q+RIDgNLa6OezHEbjN3Mhe0Obm2eO4Inf8ygPEMmL6F9blFlnW3EkeITdhNgXzU2cDz3/L193R
tWrBBprsyXA9GJFYouHIfkJCilj/EVsNOyr3R99lKZuCaXb1tBbAVdxMJ8mF19KpO0TrFn0F4IOm
sUJfNpoRC5IRWWTzTu5wxyzX+fqj6FyLHHhoULqGOQB5K+g3pFIa2VOlQtUM5uP5QJNI2Fp0eXIl
jWaMqmXWbKcBQFiMoQaAtaxEeZ/xkiOjdE4Tqk0VtrFELRqonk01MYRJ/8pUeMDWPopeu0fyl4Xw
cJYcQkRY/p+yTo8xdYZMcRoto/DoP05zGEntYDlS+4/6ohbAYZfjrLTWPFZwB/y2f/KL+VW1pHPm
8dWkNCmfBSTZ57/ISlSBJnMOv6NlPktVMvjkNzyIgzF4CO28ga7cZbx4vmyTsJsV4I8Wk9lt+3+R
PcxqkkaegCijuQcbh14wjrq7sHZRNW15aN41FlT9k/2DWMvrHKBGdYY0xxctrA+hplCMT4mj4OJ2
Q2IxNHbRD5y4iLKsHWQsDDwIoepYNNatoaExX9wFYXkgK6fWISlLQcJvLq8thEeIHdGvpXYbZyWp
M4S/9aPQ3KFZbkSL5yZDApYcGFsAeNXGmg25x2i7OAVnP/oSUenLcv26866FysRImS++ak7Ss+PS
ANHqq4TNiLwDsQN+k16tQXm/lUrIlX2YlvILGyd8N4YwLk4K0MNaxFE1UDVDBQH7t/ZggD80UJ12
csY6nun+u1TKdEkEEq0SEhPBBCUQ1c6Xs9GBh7erlQv4bMNPDQNoL3XbNt8JuOgl2hK40QHHmYND
P5Ggmmx1bWmePmtl+EQVKEKXDst2gq1vHRTmlE8pdNIuI2UlDui0d6r1nr1Wo2b3IcIBuVX7ja/u
RgBw30KQvL6PD9SdAONhBkqu6SIq5yDoPhgdh4XGCisk0OyXAV+TngOegrMhjdqoaAbhfvbWifGy
9hd0CkopuiGFs3CDQeu5UewLbaX1uWv+fmRk3Kp9IDT2CipfexPN5bUTk/KWr3P4SO9XYbkbZKzU
ZWU7eVNuRvLu1Q6m6lBAzEtOyXqNaTrX5W4wPqcWMiVtOR7k81E5Z/dbjeUgZacDQE4fGErbf4xA
jwoYVjGaHf7ZP+WVix8JjiRKWsLchHV8yQYlT04yBqGg2zHdvufx2EOrpbEtOVAnQvsFVBS4mZte
zFfmKrlU15PKJGFZcNInzp+ynDVTYWeX/Tal7osw1dh811ZqaLRu9VI1RGrAwXv+AlD2tZRA2gcE
sY7os4YQAvg9ze+ZOw1dEZzmxyUvKSly1L5YP4Irihprs/455ujIydFckzBuYP3wZHPL6V4nqUY/
tJJMi9KVsdxHb5hErkkR2YHXcoCZ6jevTnBSlu6QoC0o3pvud84v1vvIgS5b1Sg3Gd7LbWV6b3eW
AQt7v4TZHzctEWgcy9GTqMASP4r04HkMAjVarp4mEGcT1XtAAnkNYK7sIhZhK+zegEVHFebgD6yH
XyHmOmbg7On8gcr5BwknwnjcgjY93rSJAxpFGlX1PDZ9OV76k1S6UODtnxe5P6MOkltxkYXeI0IM
5iLvOpAWyEc3ktNMSZzbhNiduw0smgQ38nYq3KySSjsgwsI05MqJDfgBZF91uf+JqVHT1qK2YcNJ
J5PNlQ+oXWT3hqacRrobE2cnetWT67jteQYffytkUDfS7fS784RB5vsdpURYFINEKFRyOs8rVzoJ
aGKwEnZtnAc8hfDIiSrLhaCd+bmFKrWwTDGXstUdV5BITKocZhspNIBOkV+QdnG1JFqwDi2OR/s9
nkdFjS7fXnQbPFKCVPUltJ3jGwKoXrJw5I95d8r1PcjLpV4SBuT5FjauaiJXyjhc+T1g4Jc1rkGr
c+YF8JSOrjMMtN2afIL5EVLD68nL6dEsGFx7tmTRDg92U0a3SKkhUf5yU8nHffELN96uZp4uX7jU
j9hMAt5XU0Rs501XnA7zXuHs1DWxm/bsp3lMkly6nHfYWEN4DDrjYZ8G2JQGkzatGIDpVd1uaO5r
u7Gre1KnvlQ5GINiXqORT96iYyxXAMa4h8nXrC4rjwibY58epN5LSd6xRyYfYpG5pNALJqG9V4DU
FcXjNXttrs3JL5LC9uq63Tz8ZIrCeWxF7lnHA4F4pF/1pkMivdjLX1RQoeevdyDXPVcl5hPGJ7En
d1khioVnBPZo3goTt0ar3zTqdGY+toLaYUtiWxsyLdALv24yw8CK/tmEhKmJDxhivfCDhnvAym3I
iudk35RwfI7wsTw4yK1csYfj+5FjniggWCSloQSsHP3Pt/O5XSYgHwIuOPmFAHe7zimL9FfVzgs+
jZBAB36AqBdK6lwm8hMvupW1L4oLDO/4Vm6V03bpHfZ117hocWypmoNAuVXlAOe9IXHGzYbbbD2b
1x5kDdkVCP/43LHfd0MO24EZIPnlFa9km41mdQj4Id071DMEiNPYjic/4+N7W2u4ftDAvN8ijRa1
gYxaRq3S292rfMkHsH5eDHNhO1XqdJEVpmqH6jFKWW5D1DVdFOi3vWSs28QaJQd88zagmUXH83cF
giPFDobZ3bAB3AsFgOyHF1oNO/4bV/rT8p/QDwj4PAfXuDIeX0ZekirlqMbM8ACORraKd/xSACBi
fRHX8CNr27ISRz8gmxKQT7e4UAKW3tPNK0eJsmWJBEJCD6Y5OIDObPu//E2fddqzDeNwi0IV4jc5
0T6WsJpGGqFSi7UMXL6y5ILD16kA5LRQvzCy56z9bK+2iYH5bD5cVQ9kGOSXnRskxsEJkXyDKu2f
O97hr7jhS6yFKNO/eNTWcIFETWTB7GRgE32VrVi8n1uLY5WVvklJDR1nJ+xf3MV8tDDNzp4aRM/r
0HzVn4I0brP/16HJpAQc00wqxsUgbv8SEtM9f/085LDo/S6TxIiDXn4cx4ygQR9AbMEJ/tx0qfVw
2rr+yQxVZRuWEWIx1qrIcUSIe+m0CehlWP5kpsHmWjpp0fQAXWf8nPmtk2Tbq0Jzg0Zn1Ze8PjtB
rZOdc7jHuq1VlNoN9A4LxTAm33Fot8qS+OaM3v84Deup/J5dJI+kPf1sBPDz+xAxVSX2pAr54oWq
EQbo5TvbRU+QRaEyq0szhOMvFVVabTMGmJ9zPXWfxNH9Xy79ME6rxeBKB1f6xHX9zKOwmIrntfaf
UwzVuBD9b/eCXa0ldne9yUu02YxYbAArOU/svnoP8XXJcWwJA6T2p6wfFOWLcsz0rPl8Te5FxAvS
l2rp6LZ4Y0M9TnXWE7lpOZ+GztQ/LoYd9ZTIs3ZvKOeMWC7fhk/yQhZ3qQ1VNU2lPac3lXDO90JE
aFKdSiTzUBT6H79AJsyTjYKEXXLz9IUHwhWDeM/zjIuXPPvSFEPoW9E+8jYeJ9VyalYWJcbw/5O8
XKSC944PANPQXwOS6P3S1DAzQ4rqL7iFOH6GrqCafzhaXqIoZWc4+05AePfZIX58BhbBCsVGuu82
3GLuJUCuqg73wsPCEvARnqsZEwllrKMOtZh12dXNYrGQJ1lGxdFbJ7NKkvNdYVHbYMb+ktB+30E/
xD9mFgOwwZeDBX7CsW4WUXFKjhEsG+Xty0Pl7RivGWVsiEBZt8DxNSB+oChidOWLHDcsPF/jDoFs
NY4EGZAW3qbAR4PZN7t5MASQ+UP6yvfLsHuhpw2EhHoYQSeC00xr4P8pABN9f/Q4yFeJPVctIGzf
F3WQGPGzGIZ0hBM+gf5R9YaPnpUXa93jDH9uj+Jw6mXXotF4v2RJhQdPufiNtGMP6NS6MIl45eLX
XOxzqfhatDbVAFuNBbdRLN77f3H9UwLVqGbHYVH82FupY+31f16RMSZkVYKq9dVcVk9hMzaK0kpI
4EczbaRHscnX9cyPls0kpGwS0lFJ3FLcXhMWjAHUg1V6LHhT/KFqROMeK2tfsyjRHM3YP/t1GGxm
cTW0u841ot7yNpIFn6O+0sq/FvWFc/mvglp2d81rhmKJ+lQ6lo4lDOIeAEsvK4eYdmflcBz7vIDf
dc8iO1GTaz0pIBRO3j8KbAEoh3JiIcrM0lkx1hA/jG3eu6OSvxQUpxlBfoH1JfK62I4p8hIqyFgN
ph64IHKpXNb3cil4n6g/xariiLlTYwno83J79a5XNfp5EkhCZS6TrYLOkPjpeOazjc59N/ImVdHD
PtnGw+i9Ayja6D31QsscXEvUsCLQYMRn7ysxIvx9QlACoSVNkfGrDqY9XpwI0mLptxBBntts4L98
Malj+sT5t78pW4QZ4te1oRHWsJjHYMCs2CXgDSNZLfj91Qg04Xd5exoad5sBiydFYMbwbBIXCE6B
9t807WxZT9pp/Ocu0gJ1yCaI4r3jHuXYeaRfKFK66l9VPksbUlCqVoniyWctIEwgtcqrNnWuCp6h
/ZNLAziRhTQqQKgz+4DCjXXZ0sxPuYylaT5WLDwAbZv24OqnLska+CR4CWJY7XWsWV604YQwO/nL
qTzhTpDOWSUbNUqZ6b7CsmyJJCs8mI8ewPYwP2EN4b4ruuUKPG4O2ggtrvhPgXU0YOHWn7Qf/MrM
2ZayM3oX8KQlMzBYDNvukAKxIhqmK4D3lsdP/l7Q+T8pY+ymql0i8+9rzC9TTm0AE/NBOL/qhAxA
kwirxqf/66oNaN46sv8wSBzMKTD/0XoCzcoKJl9akAkNPsnKaCIWInLzJJPClZIy/QOC484rDK5i
EVtGUTh8lM/C/UG3kq0axwX6JENj7E3g8kB9VBXlSAYF3Ds9wF5g1UjMwXjsFaathSQhcapCOl8D
Fh+85QF7xTtcMfLLNSIB+qc1II/dIhu+eSm9dv63rZfqPjiP1i/QNKXHYjhJDWrSTE88DRiTj+Ux
BmL18nUmOLKbVRkBLFm61ISNf/D61oLL68KhARnINacYsnUZGXfDbkRHegLVee3EMqlb2yaX083N
4msE352ooF+p8rI8Bwe0y8FbMPR4LZ7xhTwj12UCQFBA9aPGSLVgDY+b5gn+joCQJjttYMqtUNV6
LFW4frIcHnnUVW/pVIFv7tVeVk+zpHBM79g5n+KTQM66D7kkvzYPCfm5RxLSFD9XpvmEi3xm0WQQ
VWFgO5X+cUIltHVwNklpNeCJKHd7OB7xm8+NUKelUi9glpoaU+rNQh5SKYnWja8lOTXclBYaCwZG
3uip6JoIbixBr4W0JmOEUEgSWo1Ppdty/pVNsUUoDn2MIy/fONS5vxM0Mh1G2lypNHFx4nTVaraJ
p6vr8w4aY9PDpmdFTTn291Cjz0sOPp60KOOkmB2qV0Q0BTQwci172BjerUpKHk0G/+g1sYBR4nzQ
d/LN5TnFhamU8Ry4ggwaZ8AkaEsj5SHjWu/Zh9U4FTENUWU3R7J3tabaMnAJGe5quJ/tnuwNFBM6
MKW9W2iWmKo+sDCwBOJpwriNbuFsDrksWzo6jHd18aIsKMgm8HkBu/NJtJkpNcetTEsRrQ4d+bHG
TKZ0Qmt5FXnV1y7O5eQ3N/4PYZgWadX2iJgeCUJaSPx+MtjSNopBsYubeJ5ZwGYLPodfpPPqaE0S
B6yn9bQWADok75XNwZsbnjzRR3vw5IcQnaIeCEWIfQw3xbE9HH2TXBoHHPI7vz5SqcI55FoP/jpI
kzvSxp+xln6xYScV73SRqbNWoqoMpgCIjxknoGmFDdScG8wtiMSloN6Gvw8kN3SK51F/a41Dr8eH
umWZULHXB7QY5692lP41A4921UQp+KHjwI3c4w6MHe4hFfPjXDCD4QVZAFxKV56m9V1RRirvRQHz
GK7yFzqOloYy+OdSCCID9dhsAIDwH//uIDDGQ7v/13vPhKxY1fkydKusyumlN6XLCfh+pSzuesSd
WM+gBV74PDwV2Ng5qshvJ7vSeeSoTwK5fs46viXxHLJkR7Uxz2SWMWtm+Sc+j9QIkRbzigw+nEJK
mnJkDLDhaEYopwEIxzSu/Xb5GQgt5S1PeyQ6lr0Jsx/vitk6WsJqn5WwDT5utzfJRM+MVUadk8bL
ajUQt+/B0jemt+WOuXubdnjfrxgMmuug4FW7X4iGWZs7eQuObAtMohcbhPCoZSiMowX6Mz0irEbA
Rcy7pjOqQ+zc9PVxsPNcpQk/VUxPlGZPmBd8L4V7BYGutXdhDeZHD/ZqeqYSn7jpfYoJeNGuRGcl
7XyV8rWeS2s4R0sH/4UsYrlchXieFAdjodjOBKB/mKkRdXexQv70EEQWvRe7djX7fT0okMdf4vNR
zcQFahUPYGd/yM3PFJItNCRLACl7XFS0nIKftXFBvgrtargTdHvoHLcW8Mst7UaLZGHG8c0b+IrL
gEc7MFp7EBc8mzS2alBTmx872WCRfdzRUSRhmHYkYZVQcmBdOlByDCW1MTlUBgKFq3NJjzFVBme3
mjNJNUZF/bIyV41kB9TzhfngGXlM9rpu/a9fkiPGpFuQ5ofMbECDu7C33pktPkL50LoeT29Pbtvf
xXh2T5YWYOtr4kemAuYeWXkFmkra1iT5O8SHUeS3dGr52nsqeUjOanfWDNcOsqurO9DOwkEB/xmN
8V6pEn/A+jgh7RG8I3JgaXTY+fizlVWyDc3gsuoPAHk7XrCydLILXqF+5XpFc4+akQaQMb/Bgtkl
DnL6wyRl6ySB8oWWTKIJG59FWEwZi/lJeOpdR2mUaervbxRsVWAMCrn+FqpwiVnCkVOMbuq8jLf8
o85lJXeclnpGuv+1xA/2AprNgT92we5KittJ2csQrIgbef/6tOPAWhyILGWPcXWUWuGD71jwdM1n
KTwJAANEq2TIk5POOS1wJeRv9H1F55MV41Cl9tsxpAzp87cbAzBLpVoElVJRQT/NjJHkEK8i87Zx
R9uFY5VeOj+DSmhd9JAQR7mtCcnBmoiqq5LD3T9gXMi6WD4Bwn5LlBe+IBdIrOondBx+r0aNhryI
7YnH+/AYJrVJSMWGmnAWLx2olnwoJ7JNzhQkL1mQNjSH0mfKZHgWXKaqM8Vkk7cbGIfYHuQ+pHbT
yr8bLeHyotf2LmyhKfgwMi6zdfYkaY2ljYNkLnoh93n2gDgXWbtne7ZuS8TqcwGwW7zdrdkrerhP
HQpn7ta2oQzaUosywi9WvZE0ahs2Z3CQISR2KZY9J+YkeN0i1v266lRT6gl1CPo+oT0QhVc1FS6Q
TJGxkz5fVId6XiZVlxoToj5XTw0xb1+aIH4mkJUGiMq5sat0afM0vgb1HofUe6PgHjrAaNYyomV4
638s7r3S/TnicZdKInsjkbt4q7pvBgDPk+igCz4pSr9dsb5Ik9YdFsolVklcA1+xbqaAJWmBiuDD
mOgb8aTTJLAou0NUJ5SJbHtSFQx4XyXeOTTHLIwfrY/SWCl017VDL2M4B7qLPcEE7slH8uaqCMdO
QKQa5m0+kCGe94TgxDJ9gwb+kMIxejevGG6eHaqbhfYJrHRTsV9kOK2HyabbOBK/ipu9R2CNXdwm
0uQJVrtWLW11VpCAoFxZrIec3mUYER3igwFyrGKOkrXQd1aI11nhqSPzqjs+fJ2sSUwCVQKj/KIK
1TPIUfqRu3tQs0WxgD1S6Dawf8wUDvOWD6O7nBnf3ZJRy4eJjlviWNIntoGo0AoNRDRmJa7LKyiA
PXRGv32l/8u6ipXMdvkuvpuN8iMGwTfBdMEOnTUU7mfnxorAyGvAhsEmHgchhVpCsTS7ABqx/X7z
j5PkkmPqipOeb11lpCfqBiuBpU7p8cd/0Tul5jhLKRbg7yL5vNUaqhdDzxOhjWZ6f4hpa4S51cl+
d1aYDA9s1vP8rOJ1tHMhrmJvsjBjwrbhlSZXvU03pSmcfzgAGSfiJ4ROIAO+nYSz1Xlp+M/guY2T
DJKhzvy5rRICQlzJwF8Q7jD1zJK4DB7fI6fOb5SisUQ7p6oSQzGan5nVrsf991uTC+bguF3QRgQ2
NVNDCx/4nCkVRkKJ/kodTUAD7jvHcF2KNLsAcKvd+rmz/T0/ZIIbak9fKMjJvdJ5oynlR6RWhcym
lxsnFOsnvn71tKn47svd3QTCfjbR99t6kunOB8eT8BdOI2wYUzXjwHcEWV7Hr1uQWmImDmm64h2B
M9t1VTQt4ZikdxoF8laOgY0iCDc3KJNldl6XNkgTtPxua6xX0T3tj/tCTRYmChbnzekmo3jPlNZt
pzj9a2UsqrHXqgj1l65XjnLABs12xnNMnSSk4QQEQtCgbnIlR/pDqL/FbunCkgWEoubK9SCwGBJM
U6A68drQyYU5e7SLytMKxrrg8BfVc8HQpC1aeSIwYc9kYim2/4q90kNAQhllGxWhnvqLH0uF8tEb
6hiE2UEw5WM/sfbhU7HKDHo1w0EXaATQ7Le+n+oOT6Cg0Vr8SoLZv8zQHbkXfQG3C9uZN4qKsw3i
e3jKtG+6szHDFHPk35nfbxAYv6GDXYevbOM3ahsWQWsH8w4Z8CUt80rbEIa0QiXxM73Qoo+hNooZ
jDoOSjNYLTztFD85pItVHhdd5O8w2Sp7C9SG5nblJjxt4SZY5ADvQ4emnQsEED5OLNSyUk1Pah78
TzhAp82CdL5sA9UN+/gL4j7XSp3dx+RpJh6jAm8XbdCMuGx3NNNt6eqlLhyPn7CKc1LXM6ltWWxu
aNZBwU7yyUTCmWOSYl33hRpq7mTsGBiv3F9KhbBqx9vLnJSw1D2sboBuIjD9/+Of8VIUS2WNvx1m
VJrV4MvYGVp1QBIFE7e9ofR+XNxrnzK8Ne1PnmH/7Vy21I6hZGrFa714IjqFvymTTeCPcW+n8Pdf
UxnwvBMUVy7sA+ap+/gZevOgkhRhLfJqxhuGLsbJrvSNtV+gYcYMMrsqwuFANoHRS8T6yStweU/P
FhlG84giHH3S+0NlOWpn/0OPGjIqVKEn8pHV8W9HAFJBY98yqrbp/MR++tSlI2W6y//oFKI6W28p
36Zt/2l0uTbho8U75LOHzUAhz82DjObcezmXxr5MMavdngUyo/qKxawAp1Dvfi1Z/L8uMOcAq9iO
XTdAItDlO5TwPeQSKrxpZ6sgfDHUYhif8o8WV8vdBI3LEoWcxUSapgk1/QrH5icTNAulkV6XPSix
Hob25qafEeLe8kQx5EkfbKQtAPISoRFGDrlvLgnalZQdnJWAU/k7eEIQDbfk7fdNVpmkh6kRsNVh
xD9mpoMVq+DJQlPuNkewY7GHucEr8T/zsTHKcWl8bikdeFyXOZdcVoVedN5mZ03BssV3u0zM4mUE
mMVLJmZAmXPXjM6vEdWxYdc4dzxtGx289m/C1nMvW9wbH3w9QN6uE7hv92heqm/Xoxz1Hi4I5O6L
uFrNcGsyTxhKthemafKpe3RYDK56oQN2/bA4iojTsf1xkdxQFkdDnGHEHzqMlCIeHZ01Ax0HlaOJ
b2lba8JgupQsidm4ivljivLyEXPTZS7GIDQSyMTFDh4XqrFrQf+53tu8QpL2LuPkM9JXfLiRrqE4
CQAsdRZ3YbSfxjl3HMnG8cdaiZfFfNMgw7Y5q7JQcreOsN2qBiRfJhaRKivjCyys1E4vBUK99pC9
IUG8gZHAve5YNZU3GYCHWrybe/8u0xf0TwvFiVWp/LWz7a/xPYQkJlocIUr1BTWIQNUmeURG0XLU
IBQqn4kp91WF1MsJjPXosouOxTu2uD3H1V9HYr4xmX8JYiJ6paDrIJLrPxoRIBOOgXSDO80ufe0g
6wX0C8S8jft6CttoY5I25Rw0LsFAzxxnrSAUE9x1Sf9oCMwoOys/0OUFQDXm6edJ2cebXPNo2PlU
qBGWs5eeRvJs5vlG09UW2eDRacKjhKuktDLRpQ8Gjzfkw5rp/+uXHW1CMNlIdUmicreeO64MKWHx
KqolDc90y+ASsqUyYzrGx65plXAlCRr6jUiXRqCkN3GYjBl1XBYFFo+Mu7ISBFt0xRojolrt3LeD
eysq9exX/6hpd2AMKFUO4qEfcCu2OV8TXZfMyb8SvRwAq3iMiz9rhwGWg+Qk24vMn3nyNL/KjpOb
Jo7Imhu3ecsTfzt4iQPwNe8dPaMJkmoKr1f+O13PiPlOtVAz6t4ugEZWAMgt/8r/P21nmfwVxRDt
hKQ5iGWl1Wkfe/JNHFXtlpwGeWPTj4XV/HDNNnwUtwrEaSmI2FbS9MGOm9qWMYN8Uiy4Lk4iWVxC
AWhli4DNRFz5Q6HDGtfXnQOmPBfaXRYDw7lnykT9KkduJPk+5kepVXoahI1TwKewWdhGncNb4GHL
wN+IrexQnzcug1w3tYNcxjM5uVm7WnWE5CLH4P6mnd+6vFojt7yF+qyaOf+aNbC6wFrKqsjrRXKS
IBc/QqvJtkELgakjtf/B0LAGcTLGg2B6N23qBmBp+X2i5+P2ESu6tCBw3MiL7VQSTNO8/Udp6vTe
xkJzm49WPcYro57yS7LJxW8taopGw5Opt+LqHaoMlBAGTO2VsLHVuOJHX71UtsSJHaPrhDsjB2if
vF5LNl/is+/V4oaWekVHLQZ2wM6zLm3WXLUM2sanetdv8dYHtDprm9+y3a9GLZbGW4Va8QJ1+zVz
CWALeRox3HpRgsQCT9OJTNA7ynVNajVZ2+X1Kg6qgxdCddIyo5Do0JeLjU1MmQUWdnQooAE9B6NI
T9hbFb2Sdmb1CvbLp6isumjQVyVqs9GpsvWAPi7ePfp9dNSNJSyR0IRCtr0VJa9qlytWzXmDPbFI
dOwo6QMXAYfBfd8UW1DiC8ufptwcJ2D8x1EOPCzT1zRM+bphu9yVaLOMXGqxYFKFe3w5v0KdD3Iv
KxnXE7pHmFMLLl3RRyGXJWEHqfDVPb5ZIJPy3i7S1yW+aIpAz4Kh0RzYI+GfWxR85W1m602rrlOc
mVVNatIwUbewHsZwnQU2JkdQLqfYA9GTFLY4xeEY1jKn9L3ml1+2FHgddnBktPKwpiCdFWO5C2ds
vdypcHcw1krgHXlzcBAgop1yemqciME/5tlPIyIhpGDeQ/e/9owBrrYvIA0BGCwg6N3Tg31kXP0K
eT/FVy1vFvUsb4A90PYa5bjDkmkNdKexCdJcP3ETkMHzuMdUOqMK6FB4o/XkzUULaPVZGz9eOhGu
8bgPC+rlDgIGJPlQD8qmq0uuzP8Ve+Or+4ARzmh04UbKU7ZLQblYSyhDUYtzs+HeUZpsCIrjC8sO
3NqHG2ftx+BF05+b6M2tXhAH//wTacdmrZMMva6QjePTKFY1oFN/NlKh9flyFa8uXCCtkhuaOziA
IpcibEYkEmRjK7qfeCFegnb7VNk+0e7e+LdYz8m6qxpfC8CelufFKUjvz8dC9cmVvxAX7YhgpQl9
hBuZ//vUBLO8Rce9somHgnPCOvMxBXlT+BWcYBWfQoy4Fv6C24ntM+2tJEiuyqGmhzZLSt3o4e7C
PyZNmzY/R7DKvZhB4OKdss6C6VHdEyKhBG6k3Y3oCvTNgwRYx3VENV8XEsYou+yQ7RsEOh5ND08y
zg+rXS9JbdClDnCJ7qqqknI4vwSrMkS4gOt/L/F7dQfJtvnYMKwI/JaI2iZ4tgtrgNXCQK92D9WX
jJnnWs0XgK/wA40IJ8jloT9DuObZxV1u9w9evvjryZdssUoXChaMCiXyQSyvpAoD+NeIPgZv1zIp
7Fq3LpENA9iTseOu208CUe/diJR3OXGfDOWQeFsZzMx76QU4sVXESlIbN2cxz7FKGK40AX02+MtJ
YOYXeJaPfnuA7M3VcDFmSVPKoc6sgesR1L7hZsJYf6QOh05TP/eu/1sP029hAUsOfAXecNICg9JU
keRaBMULe0cau10W88i76EfI9Ckqzrima809toygpOH1kTeUadKYiyx8PrhDvq6BoOg0eHfNXLSM
KTKFgaySUKMWoddOcnLTH8jzfthBqNvQUWEtojZS1hYUJsfGCH9nME6KjND449pjgRSwZCULfbOI
CTduVvS9sGRvsrfWkSGvAnct40bhvAukDz50DcWU/i5fH0ZQwnjmIVPCjO6ldmeLUakmCNDasPSb
gt2DprcO8/9ECGfD8vz/RMhW6D78T/8Q6gKKk1sqfl9E/YHVpHg+BmGtDi4hlWtxWtzRCalfaB/0
BGS+jh/1L8DeCLB5YwzlkVmFmg8FNFtTwnVLmi65tLhd2WIA/hxPov5LlZ4MibGNj6sHOUmVOply
/7topotwoiU0TMsTiRo2zcsavqF/g/EaJKZuhGry/fvDU/rlr68yh7zyDTWZqnArjryWgc12RM4J
2cg/NAvLr/8YlXhgzyqVmRq6pNpTb5pJRS15fzZw9bJVNH1M1RZ44YyaK11fSi9ek9+xr9gOTIEr
eWzwUNYkXwyYeb/tiAO76uFRvzLBZxrkc9oSACWqJdKE5nJB2TuskYFp9UP8GPUxu5/s+pbK3OOy
bwRtsvfpyEaHmIQjkjeqezqev35ds+uIvZRvQJgKAmbTBbx1mCEw7dxXxlIZ1XJ0Uj7hyVZ7i5RP
SLJNzFPslDAdO5+MKNL0p3BvgRXf2WD3QJusBFUnG1Wxe6kciysLhffGJX6RpxhKSusmzZsfhIRw
Z2PwpnyAmGr3ckYi373ZWw4BMaJxMF+bh7p85Lv4gD53jgd3hTf6+Dn/Cb/KsY5WcdlXK6QHxr2t
UsQ/XQOIH/eabNiddZ43JjIJWSfkEMCazd0gAFhi0eNe0lBYvv0wuyXhKj+ylXzkG7+hOlIRBDBY
hTQ0ljqaecEqsU0fSQHP5f+WrUJIb3pN2jF39yVNbIrAiMFaP9eoEF15o7Kj4BfEa8GrFmle9wIQ
2fl4O/Kj1xSpe5OVx7bzA02CSUdokOIhQC3X2xmsp5TWiObBCMaG8hI9wAvaeKdJCxMkNRfGLZQQ
Z+e4q7j2S0WdVTjOF6f/kmF4x2XV77p4GoQl1X+fy6XaMF3nURRzNeATAB1fs1v0mbcadGcZwDPL
JNjby7zNF8/SEGoXafAN5pKyZsZoGpN8P7SobTorGB/VXoUQ+FPPyrSZXtGr1Fw7QFPM6fZp4tAH
J/E5bEnL3nxMK31U5LJO9G+R1C8MueJb2GS6/PcAeDXsTKxx6/MFOKsMEssipR+V2P6gznJ6gbiu
nl9x7oCTmYiFeQN0Q/sOaGlHPJSVlyGd0j5YFSTUbY9w/0p0Jz3TgLD98q9wRV+lJ7ehX6EAmDCa
6SI94DOqNwa8+lTj8fjqDhws+0nSnaF4240lSfj65vUNA70gJ8vrUOgzxGWalm9dNz3g347tb04S
aSbBJ5u29BYf8BnoLWrOZD0c6kjmEnPvo9GScqGjpCfEnxDvhQW5VaBhes0wbPoosFncoij1ED+G
MJoCUq3SuldN3lbj+sJydL5aNwf96PwIVConOEdwVLCvIwMmAqi8DtqBFsyFN5+e8LkETApTGY6E
T0GZnckD2kkrKl0e5C9ZrjW0WvhUXe/lxnLVuzY2RgJHHVVUAlh0yfloKbTv1Qf1ZVxPBDE1naGA
QijnwBzTu3DXoBmBuKhP4eAvxh0Wb8Xqg3JVZ0jlyGYeVZsfaVe9oxar4chxxdKe3o4k3aisVmQM
nLkgzZOEOCkGQWlovTmCLA5UsPjnYEEkVUIket8spI/Ew9X6lUgA9L/9kVnjgiiiq491hW9vjxV/
MRI8hWUXOhQ/huz90VjGMAJv3v0Q6L5iO1jXMbvhi36Tf+zsed2yTP+qZ91btNgPiCQ/zLdxxyNv
Q1L9yP2M4yZV1RDEUuU/VYXWF66bVGiC+r+ws8REc173qZGCRgrZ793n/rQOGIuxALQevbGHiUXY
3fdfB/a7omrShluA4rYNf9guYmTL/M6NCXa9uzKVM8tYdgpF7wsVDtyWBTh2FTo0TsCPaEEIVxzc
uiIqI3VBJMkHW3fwuTaqHMl1NrauItE/Ys/dr4L1hIYFauN+O+NaHUuT/varkq/VSR+ZoQ7RBLpG
M+ITlgJPgBjWo70g0uLPXoz5Ctil+SqcneePwM8utBkZsB5j0bwFZNJ6m4ChmS/8xPXG9+OHmLJh
ezhPOmwx/olTzn1WMsRkZfrVf261D1VmlaYkX8LX+2+aWISIluw9PE5twZrjxhqhtBBQSnM3Wy40
LXAayXqddYBc6LrM4Vmcou5gz4iIhTKPVqx688noAMe9Ra5EzyYtJs1TL7G61wrsZaZh9TT33ley
7EwwxdOHg/nzFPbLX0dorrkQaWxz2kEHZ5UGzzBsev+LHyP+pZqPaVw91aeWWOjd6snJNG+mBU4s
Kxgk6/k7qscTP0+KDREJapMOF4yFb4Jk2BdC0e7gTMqYWdWu6fq9nEEYuQrAIRxp+ND69apHLg/A
1JIx3a1WMIQZY73fTrsbkFmTmxI+dPwYYhhEszWipxfLMIZwvFZfYLmfVmUaNqWXN7KG9b0aPus8
kn2M+TdHReyDGVdG8Xwx+R1s+obn4WIsPlUbi74cEcCF3FoSgfxLWdLb2SCFy0p7WBLIXP7fS5iB
TuJ8ohkUtv195NTSm69klkwFtxBDfX/wRzpfNT3X1Fn3N8Ehpd6GXGh3bAPGP0lGF3kl2ARPxwfV
3MK8YtcfSTIbDNWxFzDQVykXtYcsfEV+0QV7ajeYqn4UZI4D8mOa6I9jw4ZpC2YmGAWNM4tbbWdF
9YFyusUgAN4YuBsAAijA6JSprJeUZFTngQUQIJMq4csjTduIUEp4LzIHq34+LCvT8gtLdLGkli3G
OP1UPcg06sghlo77M5tHkCxFTRETrU46wT7lNUi1/UNr3p12vB3xBeMpo7Hn5CoaD/gyZ4ycZg7e
UHR2/BhwMXkK5l5YstJ9WAu5//ZaTaCxDDdgMc0ftwE0HkbaQ8azx3Zx7ODCbCnfqD4Mq6N03d+i
z4fTg0KVqOT91Jeq93YFjXREjm0Cgf11ZczmipxonWOzawE+/78hf8gMIAJZ5qqM8pN4isd+EJIe
HFdv2IbDiDG6b8XwaAkHN72omStPenERMHRYIzbzXM5CYP1fTrF5D1Zz14QYqabsSEJ8dgQ5yavL
O6SYitKKuyDyDqW48gud+xDiSpHiw+GbikILj3S3Hadp5IkkEZzORoxxkQwN0+g1xrzeNslPGm5x
x33/XHTtcF+oPsvrLSbFnDEmLB39WtCofPc5bymXK1wqEZcXi6303x0X5lrBZ9yCzsjcA8atgF5p
kg48UzpyWSKCkn6ta01pI1YXZgn2+rtKMLpWcXYbkImzKWySUdMeiktpTs9wnnYp9uO/mkW3lRyx
2uVgYrUR1aQeo04VGoNTdRd6zkKfnhxIN4yHRFsB3lkEkgfXEQakV+owbEh4HZBA6VR4HwnQBavl
N5Erze1JQZ8aWb4Av2ZFHPSzeSkdbZgnBb1d8K/jS5hqYAupJZCD2NvqmCvIt1NXtplZZVqFpwg8
mYVLhTLnBBr2JI8obl6w9nGKBfZXqel29FSCnJlVb2ycH+Q0jYAO3upN00qQeik3OGCPEzRv/pgk
TzuXq5BhGBoASwyss8q185Aii6U2TcnjdOll/ApccbBKp3zD9hNt4DUtgKOvqyFPUHRFm7524Ixq
RoH88y3qt2bXebvirQ2laMX9+YXq78R2djXnqTh7I2AoBFL12LxC5YPvE9XKsqQ4bGGS5JFf6iCo
jGPG/zqafBJDN40Hq57+nPAgmH14CaftmZkSkgiWuG9g4w7hqYMwE/i5f3BkUW/WYG/yHlqU4gBi
hMVAFkr9ZTxqy815fsCOpDAA/2fejW+TnKgxLfcbyR6Uchb2OKG6ho+79EeQw9rikBB8p5ES5Ztv
w4NwY/4lFEV1JjL5JDmKFTVCGWjT9/lWBCCQKxZf6OLdQFwVA5taiDrhtgPlBVLt6iUdSy9r7Z1H
ymiErBxL+JLKpdG+Rjfvi0kTiWYq3Ih7pcehdZ6v4/dlDzOsUZSVWT/hUHwYxeM9aCdkCY3RPcPf
8QMOGz9O3TQq/s8w7aDkUt4rNjFB7an8qndYQt0WLey3Lx6LrIre+RnZgdU+09K4UlPiggGrc1mv
PNo5ImPUvKFFaTAGBDye9Wj9owKK3d4DMuRiEPKNPTzmXMEBiXuvUWeJca+ul0Z0awegrsvdRisV
tIfsQM+LNUqEqPWbJBaa0gdbXNwWjBSIzCQhUN93aiWS5rV0ElC10e5kT2Kpp08f4+c5ljvR+41k
9XbpvPARK9CSNmSMThpAG2PYz4xxiu4nRWVYmYbTTOKhR3ibbl1ALZWifvtziex0UVp0UNbqPyxW
/15nPa4wB0ymlUJEaQV5VdvsZRgtmlwxvWRN9TQXvLk+ZwlsFklTRrvLU8EBKqzvkUX57M/YmhJG
nCsD6n0z6hHGZf4Yrm1D+BP26FfQWepxshMXBfd/k8V2TgMsBIWbp9DOVOWASmeNrHIiHSYfVDBE
Mz3DTyT1jXH1AYee0cAJG4vqKE5UYareFwU/cEw0QvPMzAePhXG1WMMqnU+K5YuYcwVkqYHIjhvB
GoDjYb6QM1Jij/I7+J7Qf03o3mZ1gIiRNK6X5Gp2WwZ/7w2xYVHaUwtxH42GBkAYp1fsnDuTDSrm
EqkVXKtxAZj0UG37osNtRBkGy9dsDr20pLnLGYJZVNRKIBGTiitSC6UGEAgpaHo+Oz4ciM7XdDWZ
Vy35h+kzcpYq53G9fJY79zHapjTHdBaL9hNuFatSonS5+wI9wA36XHbqN+XMuHCmheZj/prU8T7P
lcTnWW6tmfCv+r2cv1A8tRhjanR78dDaDdZ5HmgJawDmaAOKgSBrCJgo+DQNYSaTwLmnRTOuGukH
Ge2vTq3EqWjrENqh7vk38sODSSi24m4wqmdYacK91YsTstZ2rLNZdC5ayTpAV9S9C4YQDeGYu7s9
yTnWwHcCzbB9wjqtCJdYCg5aNP9hYRvA7Lm+4VNeomYCzKxCPFkyLcwyWwmZXsv8Yxc7iRKoDI+x
CD5Qxo4aiGZIWucFOzfuDy2/Ff6xxmw3H4MQTgdlmNI5QJy1CVe1KU41fo+LoMmuE5F1189gYrnz
COsy+WOvsGSgkq9ZiuEuUUei2Rv09abq6dg8ZV0dDbGBPYJmbzp3oU9yj0/doj+awX80rDMIS7Qs
15D9l+n5oTnaDdXfbg50e7BI8CpV/om9YelfBg1CBzkWqrL2fMn+4ZA0ExK2UBHpVUI8NrsY1U/b
6HX6kpiezy4eEMzk2Z20TjeA+p+qp64BfQcsvrS92E/FK/6eZhjzQL7vvRCe0UQsJVd4Jv8KT6/Q
ZqsBfqI+cXN32EzuQF//C/NRoXrblt4MgA/gG34v1RojnTKHL/OkP50v4CTpvlCRsvBz+pelGRBD
00DN0qw4CGPMgPK8NHJLXV3ZjPXE2HPq8cfC0lHw1xEXlduynIE84kSwW51ot6mFLCsAhxquEPWZ
ydm4PN9vf7xD6rn8pW9CWXgnBeAPREJR+7EahCvpf+Pq1HbBV76MTIqBbFOkVDcku4bJjC+zIG4D
DDvNHZ5BhkezwoOf0QkwQbD5Cr2vMNykoMKISb/IiPY+6U4e5hXxjLJZIxRxnMJ1+SYaRMlZ+Gx7
NyAgzZ71o8bj8NPXP0gQiXiDpEERTBb2VoIwjWXCG62iZ2Z/ANGB42hKHKlZQFVi7SiV3qTT7ibE
pT2uoSBOUeWX77eB5/n3yl3urcXW++GaB8spoqoxCJS8AVcs5gh17qPuV4iFaVgZa4NBTlCGANGZ
bcatwBvKjdb3+ETygdcvBqlfBEYuCDiPao/AbBM/k4GSCN8zgcqAzBb+Pdpr7sXu+FIVhY/2bPVz
B82v9TOq1zDRpQoOOh+qLcRl353wRujwlb5ciS2bpXhJ6bx/kHYcnpoEInWuZdpCywZItFH7/4fN
lH3hDcn4zC1bSS+C2fbyEvDA1J6/Db/go7BALrfRwIr9X8m5mSZfyHULOFSlDPj3vosDN+ljvhzo
L3kM5ymx+26GKZrelylo0sQiQzbbpKff9JFl9B0eSLqEXbLNy6RYJJyu/of5Mdv0s0U6epMH6TUz
Rf3GfnqJf2IjuDIGSYrx7gSxmFPDMeZ6Fgtk6ntn71aI32v9BEAZjuDSJr1L/DMemKdFJ9N+oYa7
y7o/8c3Ogo23RHhuLB6q07RiP4xo2x/eXyRUqOAVjgsQXSzA6UHLCMbad0JdxJwCnORwLLi/h/1B
3cb0nnunYkEdYi+bbk1YeNWKADgA1M71AMM4Pp3ieUdtJVFLLRzIRnMuUQ2LOMw9thAlQXbMKfgS
yEBTcZkhoegm+QE9MR4UA9CNcKbBpOw86yQDU11/grTlfe046bBb2+54o55f8Em6JXBKNQ43iUvz
ulWvsJRpN92BKIunQweM5fDTobMIIhETjxCmwEUoiHX30g+Of+J1ysneD+A0l1g/tlijY6yr7hNx
rgnndD3JpJRh5zxi9SAplLbsLJZqXsLTFVlIP13IyuEL6YAzF6YILHL5qUWAaH4hLPi3+SG4Mmz5
u54x0Q6qvFqdOpFkSHs3k68h1E1izD2sMQc8/e5958qBNrywXXkSqtAJRnDHGJ50kaYjmbB56iiS
oouEL9ht8lnslKv995f2bBTAvi4vyS6xsBqkW1Um4gvvKE51C2Mx3BwZtGisuLzinXUgYq+LFTfP
V9SJjlAXqYtM4Ss8o0t4mwqSAqzI9eHFsAYv0HDdJqLwPVQ+1ze5vlvgkVS+O2PDXkf7OSbzL7Ba
yfsOPyLdNCLtAaFm4eeOs9wlLT3QG7ALQvEzeIzhM/vxgo1QH89/jfpy9902zjOMa8DWaJ3gwrwz
TQrGwjlh6bRwdFi7w4O1eS/seZQVY/cMJafdomSMRhHtB5uqz5qM6eo3VHRZrxK80XbpaKk3lj8t
I2rjzrW3hrncYaSH5yDCeTHExueMIbC0tmhvzFs4nhw8vwC7tIGlB2vZ+eLNMsGgclgvmObKvJfH
3Q3WTj78veqADCdcexqXV1xopDsFoAzMICt2fLPs1VdR5q/gjDKVcFzMfP7k69u/u5/FE15rcS93
BiGTANLVyMMaygDvpE25uNDJ+CcYrmrR4UQZxlkjp2iSgpOLh/XCEdJEojLikyhHLP34JAZYoRK4
MnPwc0/+YYIRYt4nXDzZPLI97VVcPzV52NQncqreD2uOdL0cC0zOoLqS4HjrUFU6ZHKnLbjGNvbW
TmHkmm1vpwUovqPwrIwLUNseDAT1isosfYr2fW6QS29P4JhX3XeEnJFmbtxaKZSLYtPpbKOBVQSs
u0XRK0hCI4OsG2db/ir33tDv8hAMGRj+/MM5tBtAv04nFqjlvwv54Jb5cSGs4R3jg74DNp4pf/E9
cRn6TA+bhEmfStpKrcGGJf5dIqFNQLFKYN4Yp+WvcsRM5+VD5jTwBuQ4HMMqaj7NnB3Hh41PVsom
r3uJhzoqUkzVW5vTNZKRoLcHPzAlA+HEEM6Hz7HUN9N5eCnusKY0pgFfdx8ZIXveg5R73iHT2lDN
COQXJAgjlT/G/XeoZhDBanLyGiLJvGaP2RCONCjy8pJhBRHtg0y/jeCbX+KZNFzhIqOZHb5seYjy
Ha1SKxMJjA5nZ5aAaV5ul+ny7nFUlBsxW0K36vtFqTgeAcBq8+M6Oww+aGXniwveJD4U8GFDeOoW
I3827SUAquY6h41D2Y0ThQPM75QsJwUFfL//RDQLaJIpC1KZsED+TJv0xBM9iNC85L65CZI/JPhh
MrtlRm/jFzkmMeTfX5Q08YdjFQ507pfUG5cq91OuKs1sBGK6PtX0/0Jvl4MxFEUhBssxlseIf/Fk
y/Nb5Sudj1Q7n4zeYL6XnMnt/p+f/EyWeY9IGpgQEh4/IfwyF+7E9GPDiOa8ujWt4+Inizgx1ASN
rDVrgWD22rLNkLljNTOnTVa+261ZfnffB4UdvyrND6sP+by9pUNm6riT72bcczikdbSjrj2+krh1
+aEZAH98nNQmWwfeulUp+ksMFsjdPHpuaTqGx6axccw+VK21rRauDOYR/y3zVLK1fMcIhoGCWTyK
PfmIcvqDZ0J7IZuc6wcy3btJ8h5vbDz0XaGbDLrH9pOJZOYf/OaZNu51+LqmOi+13JdjxniyUF8o
JKLdF8ayjhQeLTMLp4wYtcIEsq7nHkSP1LBuVeM4vXtNd/ECDc0b+lvW00hhbrnvmiCn46n/SjZp
hx4DW3QGvwslWM1Bdt+CWBuNjDwf7LyMT3rCJyGeuqMgvd/+V9kw+kNG500shDp+8ceKcqSuwz2Q
yO1YotmccWyui7D5oYBOt6OB8sIdzmjL8OkDNVfhJUaiRJbCwOeFchYkz4+giF9i/EhVtR/cD8m8
ZsVlfoybS7xFsd/DtzJavGUZ/44iw5uJE4YcRpZAEAiWEzIOvmbwNYUkQOGPkkHPGKZtdKaP6YjU
4S0foIYiGbw9MbhiXN+I9oAWLC4465bh8YvIgV4Lcextbu5gn8cY2FcUN1o1YYwc27d1pfnCi2Rm
NVdLddnfhtd02niAbfQL5Qyma+P3mwEpAFmMP1TPXR58mncBbvb59vE+A7S1COSWwGeMVbovAnyE
p7HCSRfosDt/UIBlCzyWD4KWiRoqrbxTSvC5xjJicaoxGHdRcWYC7zqyYZclmfZBmmb3fPUQEND2
Ja2SXoHqVonHGy+F27NR/k5J0RPFYzlNi8YtA+d4eYtaBAXHGNiqS0z6JyvdAaNXOplgX/tYCeeh
ua68EkCSjI/GiJVPLFs4qmV0FT2dNyjz1R1tDklavkoLjk4aeIVm8hc3w6tMd0thX3Mb+kNmti/J
PIsVDPnZgyn3ZEpr/1mLniiFRW2YVwYeRmNBbSa0aktNvrNE+OHc/N27V7V66W+uOraup0aeSYJY
3uLa0iCP8MdG/9D7F9OD8yqdJY5ZWaAgfuOOVPEjMFbVuOTKNXyajyCWxJfeUPQ+FAEN+MTwxkvv
i5omwqRjp0YYPI17R64OcbvihOm4/WAXjZNUhtkJ6+lNemyxPBm2qXVfbWfyp+hty4TAKKtlWOg9
UPBehRtLPhJxoiPLGozF3z7y83E1cZtiElkqi0IDpkki+/dPnmqdFdT4AVyTrk8oBb0WEdNLLREg
PgkvKKMRa2k9csWGhCznAll0PyG6ki5xUVn2SPsuyEEzqINIgyoL+t4Ji9zSbncgZePG/QYsZtsD
0jWnkBKRMuqE1mqDTrpUfPJP6NZDat/1lOZKXKB4RBylzHtwJy+t9LuL6spTd1KhDA6So3SJNzbm
VDPb3Hh+0d67RLA/FFQQnIeM0FWWsX4mW8IGiwD2xRcqjHme3rfqGpX8J5t/a2u+0vzQv9dFhltI
GL9lru+vjGTR40xZ38ZiIisSrMz26WM7KPoUPBQuTuWYE28k28AgF/19moQ0zuf2qg5dHTDxeIpJ
L+9Sb3Y/A1QCynF9GHeu85zs9tt0KnxqZhd4qczrnUhNCehOuvO39WoEpxANJdALJ0trkQdmGuAF
K1lRVoPQ+1eWgqIwJrZtsm20Jr66fSQU7xA1kbL94cDJOJUiuYtPgMMX+F20HlvP1c+ZywCDab9n
yqsdLn2DsmHqIOYClGS9NXljWClrqnlOCKm0pcQIwJbdwrB8QFhNkocs8uniQ4mJXCxPSOOfBy9X
13WsoTus0PEyjx0t9vI1My5ehnusfyNumd4UeiBisFhcK94EQdhz09gpUK3S/YhrIiLAwrXXD65o
DKCs5Duc59l5C/nFJwSE++pi7/HB0/Nb2jcIGZ7PIEVNJN2nC7RILu+cR3GORlTswxtGeM6mFsxg
0hemvJ+fVV5+qfCBGjemumtaSA++aCODk/GYewZJaZu1KU1+mBJbeD8uOFLnUy9HTahF7maCg6QQ
M4lcLJVjERKzidOT1BebaXK07hXdAqLox8dIYwsFOcAjkRHjVCD5CJudxIBmrFeTA0X5C+Yi9Ysj
NLunhWEMEnuNUYFEMAkuAvqDugQf01Np6IwoB9DaUMn1TaYSPPg1fR1JIWnMh9PdtYcdf+jFA8O5
FBD7KzdXek2ZOtEmDxNAQWvWJ2ScujvSAZd+SgHZMVbcNQShDnjvgigtMbq1unc4zLrY+J/EjGK6
EfJerkEXStpjaoW/HCZAHd6r8+rncwqPYHJaBTLmlqqZexXulaco7MiuzFIO5KA/nWqdykxvGpls
YKdjbfHApK5ZEo9nCYMjymST2EpjmuI3KDmEAhPK7FKIFujYMjtUXezPVveyRxQBXFTkVmCUBkBQ
V6tjh3D37cJLZdrFmS0ivmULI2QI4MOxpgm6bMu8T9wzeFe6G/XSRW0dcYyx5qG2l8FjcbN1JxuO
G3/lbvMNZPwaAKKS2vFYG8h1zoFklFXtH8opA9IMkMYZpVIkTJRpNXlOZs+k6aB7U05m6OuHS44O
YJZMl4diq8iyfwhLVeSQ7yjQQAkXVOCxXnC8UIrb2IOEOHwA682Z4eV4BEVhTOERBMRwRtDsypAH
qrW5PmZYHT/Qb8Nx4YCvmWnQfksO7Z4KcGtH12kBQM95BgcXvTNhT+dJAaZlfGZFFghHzGSjo1WG
U8SP7pN00zDyeqyG+9Tl3V7HO2+KfUFK/LZjOCedCrO1372bK00Kdx+e3ZPuufre8qE4uvIlb/Vd
WPzK2SUgc2xBiYYmXoaBz57TrdreGK5tMoTg0phuD/rjkYs/+gnsmc8mogchGkWo8w43Ht5BNjNd
GXF4VW/CyNlf/N/oLh/32+tuDa2G7HffX/3aIHZqZ8eipRBCOoj6PSw9v0kTScIi/whPY3o4gQiI
pBduC1gPxIvAi6pdCxnV3GUtQumE9Tswv/OtGiQ2VD6PF8M9oumIRKkWGxwjvxx5Xj8/pPPDPfHz
SrAuDXDp8IS7l2Q9pNkoPcx7pL7JBlwW6UXm9EPD9p4frp/mgwsK/zqDWpfG58vUE29u5QRKgdUV
Ql/j0iCTpOgj5kS3nSzCzxyLT/qzm6M7j+5he9OpWojRE7PQr+8x5gwHsydiOPq/HnJohkqwSn+u
U8Bg0TT5wrT5dvVcsA8w4nhUeMB2U0oLCfl53xcbd1ztI5cD93RMciWPlJKr8tB1wLLgz81EacUc
9CX4uUunIPI4Yr7g7BYwDrbNXwUCRORx1o2BMIUDp/5okhAnnjf5Tz/J+53oVP0pcVFcivgYiC0w
16ohchIaZJIhKUnCBD+COB/nxQ975hkpvMe0NKxp4IbScrVpFMMNMeMkKfrZKH2ZUiQ5efTtoP6U
4HH8nDFlo3XAq5rzvs3He9G/l9ad/a6r0gEnGPWr7v0776/lpWLS8S+S7RAzdBTlk2PthuParWeR
k8TacSuEhTY9TFaCo/tidxMbBpWt7/plK5msB9mjG9tkkl4wtuxvmRDG0VMGKYhwwSuNvDSxOLTs
/U7eOZ78FBpvHv/8nMT/iADoefDbcnlg4PHk1KNPa3h8oh0QCUzggIAxERwVQl2xr5E1Yl7VG2TF
BKukXeWHgjCWqfNVnQn8KJAgOg6JKB6QJZcCmUhpB+f7ouns1Hnbl3GXUe6a8i9NjyV/cGrhO/Ig
WIN8P6EiAsr9Ylkbofh7Dd7gKCVKjT2DshCh6n3mkOIoF9pv1XJqhhALiCFtHX5fmAtvHvYD9CNX
0b3zRXHLsbeLUwCStJWWiHMtDMyky6TL8cywuayZXNjISv6yFe8/2LZ4wBj5QpyahfjZy0Rd7Wyt
anuetthMdLCJnofd6oHQWZVLHkCJhfDcElIWGmiPBekCEML2wNw+4clN82e6WCd3Be4wtVhQgIpH
+bDSDBWzvMY27hzTruvzeEyrM3GKnjz+h7Q93FNCYZRjQYwQpjqUsSaFI7MdVJNjl5QZ/4PZc9k0
bl8JIEOhrx4NZFEDiTkrpEZhecxezAIz5Im/CeCPtD84/E5L36OXcwJqOWJo7J9cNpvHa4VLM3cG
Bscphigu4KZj7wiDHpg2YrNXG0tFN4yhnFAPkqJZ8hoT0SsaXryrKHZLLSXf7irv6UMKyjjT4TDE
gP0nkeFZtilv2A2KxJnbdFMQxz0/gQTDdo852OrM8g0qYvHWiCxEYZxUxrPVY/+2g6eWbh77qCKK
W9TN99vpdVAb0psun5kUulI4qhBydINDaTlgtbRwWXXXZXriQtZWEWlolMrvQQehY3Gb9iarckoZ
CxBjqM32gDoKCarY3odmbmGutAWRDG6YIxm50HSYUXQ2S2kHPERaV6t3fjFsKCTEe4Z9U9+UVDzJ
Pgqw62TySjMNKI87C0sb3n2rVhRcs04VVAIBVLn/MQ0ftSbhsNYM9/JG0sBAD0Ba49UsFjmm73aP
3+CAa8lqNyosiLgzCQpnltORyfjEH9vudiYfbSq9zoZlktNs20iClC5Vo7pGv2Ypb1HenOkHe4d9
Ccuujh19VjL+1uQF7Yx1gDysrXtVlcWES7SJ+YyEbdo6YQCZO0SOMN8DTAmF7rx2csp18hi1kDfO
k23V9iaacv38oNZAAG1xR/Dpfv6M0chFgrZJFdnfHAf+iDS9SK7PFUfScbvhvJu+eF+W+IPRCLzO
SySQoHyG/SUt9UDUYOFie96/pwwmZm1wxWEtbvF5tBCYOpx5rxkslVmaN3aIMWRcQmW4bg+BbhjT
SmALwRytFNnYbdWg2LsQxygt26a/dk3hY0qHhTOyn4uYth3tj86LglTEFTWi5ErBLp2Qzc2i4WL5
kZaqRlJ+kpCEvQ4uvE5r819K5lpg6z9MErpksj6rQVItkZfGspwEwrDbAvtfUDIovmdSjcn1H2QW
LbE6Fmv4B+Sq2jDVYI+37/Qc1HcVJM7o2vhUQ0VWzD4Pg9HO3JrfGVIrR+z0kbAGdULG0E1X8VOH
ao9Y/XevyROCGyn+QirPZWvsM550m+MctugspfjxiX6dyCIvWIsKcrK8yYfPsEuJ5oXbgzG3ZZBO
/3WPNd5G73AY3KQym7ZfhYtCeOeSx9poD42oVfB0coaIx4/quwVKxtgWfrGijwX3qH+f8M9sJ6NP
0kFBSMXWVerUDMXNptTJsPre9oIsbgZvazf7VJ3JT4QgysIoNXTFXdvZEK0O4++XXIhHeY9O4pB8
IzcfsIouN076zVB1hJHBSlZonBuyswOTXEB574G98zhmgOtRHANX1UqN6H3hduVfTiJ8BPS3t0BR
cpLTBNfjIgN/MDGe0JeyyNOpWhFBtDMn3wxPKXJ+SlJpQs0WeG472qeVZGCj4w2/UmBEJ8gryfC/
45O5Ssy/PH+3/HJ8P2zLGIRiu+P4Rq8zyESYFvp20r6nilB3jTR+E60mOiN4xVT17jsaLKvP/RtT
pfVQIK6BsNSlMnHb3SCQf/lOETIm9FbXR6F+waxBb8IQU3K16rLNTCfc/fkXVQ4XUsVaa5bEz5zY
q/VnsVqEx16afBTBtqQCdGyv65KSv+XJujypXScvGSlE9c3uF3nB3vdDCjnlYib7cZdxzLekhrLN
pCFf0RHznek8OWXsX0l3XZnCh4wVirx8cx6ciLKJY0K9ko9jXzbp03DV/j6rI85avSyNskhFUSZT
OZW3Yi5odGesIVsUsulhxrqcHL1Z+pPCDjMsHYJCRUHI4g2MC3JwNby7gNyz4vAhmRoehlm0Ons0
bKmFOQ0zPLuMwXbfCoHGGOQnSa74kMhf5+OKgX99FLj59UPe5WlfWieE5VWqesqYxCUumDk6oZtU
NLKIKsL153xQE3kwvKonIIaW3tBoIRUsIoxjG5trmPzD8vHUYfKOtXQqyaidwnaqFYwsjIVkAlXz
PVDMluU6kyRSF401hySwWu9TkSyiwALbpcoVGIvDgrmS7T73kQYBM4Kg6Y6IiI9nRhiz2V6LDmmb
MuJwRLk98iE8Ujjcra7rm8xG++6CvLhaAiH8EHVquCxe948/XLuUjBYaQ3BpcPWhDEDMWh6sK2SQ
rlfqJISIcfY4Zxsf6+oAIqwoMN+5bI0/cR9yCJdtLmQJFKR8pIduvsxQLVFSGEKkiQAZjODH0KlK
aJEskyKkicFBtTaX5J3PBSFLXGRh5gaGbMQ72tUpc2rxWRywgfmQE2HRkRF89Bn/zlgnEgVo3P9l
mksVaNcqATwu3lYzvhvX+a5Jf3PT84DW8CLujL8P3PQntf40LD0JguYfZSK+AnCMVLiQPR6q5Erf
8cSl3a+Y50Iy9CBH9tH5Ru1t73btUNgPYvO16iPV2Agd545aZHW0ystMQ3mesMeyc44L8Eo6n1FW
HS4T0OrdpweWe7cwoJrTGyBUxiKgkuuVznjA9HtjNKKTcw+ZczMTEta/n/CbXvgx9no1dlUUlDsE
fGEfRqFT/mXpg6UgvB5d907HWRC1lyP6BpzyuwOjORzfq0cvPEyZ4Wsneb/bSPi3rJC68yIztymo
CiMUmTCKa+bvVYAJWVml0vrWoX9gmd7jh81iC0ybOLcZMatx96r6Vu5df7KjF4ENt77ju9nsjwlv
YDkjzhouY6heemEgplFZeiEnTKp0VDPl3e40elBZl041HCvD6SCy895o2ExKcicSO/H9anhEjlNy
ClGrvOQ6gJbrRgc6sv5K7QsON2qXUUkHs7O/xVdQMXa+j4e4tO2McCIbjlbYFtmtCLsgnExwTH0o
EIFfbHbK0WscB36rR+v/f7ui7BDosJx7htI1dj3kUwmvwQCP2VOL56svS89R183v7bTa+CIOosE/
1jZxAGhMSC/MtEcE0c+3e25kaQC1Ajm5Vt/VpduuE/y1EvdDn4jil9kHyH8v8ToMAVRFrTgSWKDq
lpMHOWI7MPszjfc5kU9j34UF3zbuxcBi2SzoVC9rw4/219d0d/i8GkNy564hGHHvBN5Fj4NXsPKz
72mK4pBq13n8p3F9Hlt4C8SsO/kgSaHZI3wO3vGgZ2tGewdJ1d+ROv2MruNP5rQDORMvsBbG7Yp5
sQbY1HRu/ZwfSk3/4bZiXzk/hfMQPlfuqciCC2mkz7tuOX+E9BgGYDNu6Cqu69bmm5f3DzUHx8o/
ggZWqQvhhy69u2gYhqrP36EfE4YOkaxI5cYz333La1a1jigLTlNnXiQW/JOrvuhMIdY6AqZbHYrE
MZzdy8lzxRXqEQg+hh70oig1Xd9YP8YrgcbY96efZZ3endyQeQxdEkPrZx6X3E4e9G+5pN6BfJ5z
W4K6kZ5u4SZ3Mi5gfWu3WU4wCtHvZWGWPqmrY3j5bpdEvl0eEFcXNIwYABhLnQUg5Bh7Kf000Xyz
TGFcfjjZD2XB30gzPopFXBWRxTHv+mFlPO2wqL7/BrfnMYPZjwAMoc/2PMXdpYyM3tPZEr5tcOiR
5DHzbtJlIa/0NLiVeqA8wXc9yUObzfYBkhV7ZWS35HI65qijWygk+8c6p8VJ2ip88vSJCVcJDqN3
ufkM5Nf+qSWeoFApRhELNWyO2oR85lMXOo7COudthasMbDFGWUbDfVJ+pk18/D+Cw7Hc+Ox94ZWe
21diVx1+FQp3BMpqEV1znJhvNanxNgiHaOb3Qql/PUB+VTGAOysT88f3teSasZ0W0grQlyPL0SBa
ZbeSQVOMzgz43KDpW5Nw02ZT/egPLk7QpCB3nkgEcd/oAh8AjLQkYCadlyZbtc65Ls6xwM1dI66k
P99cY+k3KIGnPEP3AXBNiVTyG9/g82CKl9wFE3s8edFe2DajAAGqsj5TmgIDozF6xN/L9Y3VkTuF
RaH1/i9H52IcIQiOgzMttzGovZpXwd4DVFsKyRmCux61kWkStpwlpAHSVSwMSXEQDKed8pzAZCA3
kKcuSAqrk/bbNZwH/JlQ2UXD3WH/FRhrnfFdsMdPC2UVZeRzW8nTFEOWhPkOEXR1OGd9iVr+Fgnh
PVfqU+wth+9C7abEWXMj4n1yt699cZgNvctIALVsKkQ8zLszKAoa8xIR8l1enaC7cJAbJYEjf77z
K2EpVSZ12IE0ddNY2pYUmiWpaibNep2q7CHanijDZgogqw213aOM78y+Vn9VoihToNbdK0sVgANd
a10mJ3YMVwHogxR5zy9yNLhw2MTP+F9xVcRMGKzeucH2SRSYefvXoA6M2Oga1cIkrnkLhAe8QmLp
7OKUO8jSvgvuKCJh0S6rmAb0vk9fjGTlEEynUtG7vJmzHgCytnAuy72661TWti3wSV+KpGrKV8K6
TeiE1W7iAOJxKrXJKcpX0frUlv9jcBjAjIHic/MFz/l713huJryO9wUstBZ/ajisII06d4/cAzaC
EvLwa23lTA0hqhpKb6X1z0/BnienT4Yulck0ZEKCWkmZF0uqmr4aKQhrG48mQEt7+/zKoGIkblEa
oU8Vbyshy9j5E7i+ZikHXOzxnMthFwDvDkQVd5FDMRYbwrY9K6qG8Ivj89/ziXlE43CbzbvFthDy
4NV3oWkTDN/s5Ld19cGH19j3/Q61R0F3zhqxagd3DUBuQ60v1WW9xqJ0IXdsT60KUFx3RtaHFmLN
M3+uWIQyc2p4/a0cJVlpF8btgt20k8TWTzIa1QBfAEw3ZlwAnri7wxG88bXwnNic6/8lmeWvP2UX
hmHSCR0uFdhU/zvA7zO+vM982HTgqFPauOwHSH3Ltg+0rdeH8aflpDmOW0/CcnNJyI2/j1OXMSFS
0M8HX6LRHPVGgVQ33vO3TppGbmdpEzJecsS+xKUGFdWybFUhO7Z8NiC4UefHnQYui5wiuruNr7Ny
d/gcWo6QQlk+pegbwaMluTA5W7JYcGSGuJiY0gSvVIGqFJZsph9GlRTRUdL71jZxNhImEha3P/+H
d++/38kJXRy/PrtA1EN9luThWrmr8Zbng1gSI9BBLIOeWBr4N68sLyJW4SxOyMqeqHkHZMy8LU2Y
/lUm3ziAE4Rqkh4Jfko3PLjUcCYE0rNJtk+Th3L1B/16j0GMDzYkgPfXnN91uQJy3WadIbn7uNSQ
haJCx1f1TcgaK2nLTHWPnFhPHd/pUCLWm7WTb4RCNgwUKWiC/oKplKZpn1DFIQBBp5ipl8YfhI50
l7vsofDnHmJg6IRPonFQeLkoVg5HfZq2VIY31otckN5pMnWZgkOxIR5ry/4ZyERX0VgkFU7z8Wvh
f3jVUr0PCVgtfNWD3Oat+ouyjA8gw2pGpmpq8X5ifEPwvxkFlO3MRkudSk/KwD/nMMUqF1juiQdH
9SItNfX4ENf2k9J23Qmy1k1oSmiNhdNtHFRixnV/SBWHKs3qR06uTBRoUk8rXcS3Bi8n6zZnc7XX
yF2Lc1Grmnc4DP8ZSIuW1D7FAUoqVJOmNF2ks7xaziX01yH+5yEUCXp1c7W7MFQBxNrYMrRtPR50
o82wV6PQ38e8INUanbdyRniw9hAZrOMG0lF43eY1WZBssU2GOkyb2ro7RuhT+7R7FC+9aqGNjijb
wvDRcKPA9BJ3Fo7qJEVOasfij/n9JBQc/6a8vuZ3B/gY15CUMTuOipaqnBHgjXCyPzAMkX8thWw8
AKq2sKj/2+w7/1W3RF/Td5jKJp/Cey3xuqmrgpKwLVJNeYdP0NfxDLV1yaHDhmzgq4QBBOS9tcYz
8HxQOhcfyeqEL/ErQ84/ZDzlBfBFcg1EhhkJMWaNWMLC60nYEu0ngsHW6Cq5kOQURMWE5fdjKVPo
JcpSiWwpB9q5H9Z024jwxBee12uEAzOOcR5i+3Ncz96bzQ8rpe2EC6vHUl8dAioxcgYbxcboF+zH
ou03RkmzQnuElgFUkMXfYXGRBkUld3kFw0ITpjEl8iuNJbuxGKQCM+xY55KZydDb3mSwfbo2pxfx
9IwWpQI48mvCS/MWFpYwEE4CwLx9SC4azgNqkZwFR0Y5gQU/ZQZPG1kNi0/bHh+JfUeMHCR267Kl
nNXuyVNDRfV2x2EuPHl5jSR8ETgzNk1KytgWRjc0OK47bpyqsN81bTrbte5qP1fL0ZehT1FQpn1g
oOrhi9PrPKtnMmjusRzMbQ+VwEQdKH7tO5uWRdu3bkdHr5YhahU2gc6pSms/85FDZtH215oUstSw
Kk4QXU2XaYtxkth5MDhvUxHoKXnADe1Jkd2yXWkggJGBEJ0CmBZC2I6Bsee6imTKozb15NsMCwxV
VGBIm+ziGTkJ++kMTRwJJU+lXsPNQulzzKemzzgshf5Lu+ab7OxnH2WTItxk/SuMkCNBO9HQYi+R
uKav7XjeNObYdNHwr+zhQnCFbBdRD7ShXdnhFjcfYfD8fqQCBr9wJ3lsaWin/hqglZvgNyvHh4Ci
nUYRreiLeoaDVQ+CpnAazfMCZDqmtmF46bAPSrX7autk7cvoNMMUH25Nr2y0AI+Y2TUjt9nlxAfO
pQ0otqMqjI7k1WFh1KzpgWXXL8wdXxr2tYOITD3lwrcAGLghpcA+bmeZpxXVcxMSCp52Azyt5j9S
p1P6EJV+Bhd1CZ+qGgLGKouLMF7l/Z3RttbDEmlquJnIS96DBew/pJdnF1C1+lEcAg2r9c4zHsJa
nJiKk0kQJjHKQN8PELwWIdfDId4wIWE0MWAbFIrqKA99orVaevqUdYuGn3M+YyREskxf8tRZDXCB
cpvPNNxdE3/I7AhIPopJoAK1i4eLMrnzwAJrMWknAf0Ra0+dQStgkMi8UjZ4FM2qTzVqkM9Acgq7
5Mh+lEVvj4gTdCYKUTaUe8jP3bwHBOU1vuMT6iDBBzbBXrOcj0N7CCk6WyJejbfekwF8M3xneRyV
XbnydXY/xAgeS/dwmEKAx3qc149hjrs0Nl/hRQvgsdl9lyjhGbBXsy/tpmKLgSlzwLWZKvY+OGhb
6qKqgJO11Q7cs4axDraN/14BwnaGiMZAIudn2gQgT3vnGASO0GNmd7roT39pHd0yPOiJjDPO1K36
bX0n9AUxJEUqd4fXoGOdRa2HnuEgEqpxH0D/OazV1rEjA+VwIzlT9mGjNMeIDjIbFx7FY6oC8sLw
w8546i2AgedZ7sM/CwBtCOY6dX4frsyYpvwExHn6ObW/ObmUQe6HosQ/mwS1KL38GUs1UAd54cfC
7tNuTpZVhpWMmdMaGLk2q6dQLQP14SYFTGd6sojB/TeYzKZWsgHalHwaYLgNahvyR43rDa7BYJrg
Cz8mgudaA6Wdhxxp+SrnzS1yWRlerp+qHlHZ5kKZ8z68X1At12Cb+6PgJtnHAKrpG2GyFkvLl4G6
9p1b+4EB0FyWWJWW73vUyPBVaxHrsvs/QqCFzT89PdMEny9JHDW9fKpnXWCBdmeH1zK0ftoB+Kd2
lBQa5wQ1PSsfk6Dt6FU3MDBFt71xkYpqZ4JtZU7yVAZVL1NXzv5hNJWmhmY2zNxF63OB8FzdjZfo
rCJXvAwuomnBvY+Ba2kvHvelbXnnXEi5TOCoYOB4ZNqGZ2WvPZOGTnCFFo8WfGB9Olx4r0k2Abg6
8ortlHx0dcSEIFJzY2i2kqXOgl8AG/ywTNkG8tXLa58nG1GQMpWFaWKL7wG1ERxuxaLcTiWFFmYP
HlEu0javU2VAWKfE5xo3PG6hMzi2wHE63wDW52Sl6O2vpfhrN/+7YTNuTtAQ7CAzssAMKvnEDt65
H5ANuIUsjPZIK4sZPPHuqx+dC3MSnpLRSgmSOpJqFbNlNfrhIBYOW5n2u+0Rv2gHNavnHoiiJPjS
Ru9BPlzklS2T7giUndKyOAGIYQif+TGgIccElf6EGJ4IaEeB9HceGlZQL9OOe+woy7aMCugM9uSp
3YMyEpfyI+VdRizVgCPC98tox8Y3j6m4q2O72oI2lKuug+5WFkblh1xCiP7TxdWWnDGXJMwcxwf6
M5ZDm1ZChoMtQEXuqsS8svV523Yu+RcdZeZjhbDDx8RbdgudE54fwpBD8o0Qka7hcjPT9pSBFNOp
Kul90gh3mx25sxYi5iSmHUgTCMTR/SviNX8hSt0d5R1YYuF93L9N1IMaRgY0jA+Gsp4yrEPkIoV0
TBDacODAyTf3uW0h4l9zM7gapKXkjh7fWBAyRaWA7sQIBkQnSs0Z23i2jjg36QkT+Z6wVzCNI3+i
qcJTSbaPbAie5meXkrEd5ax4yTKj8bXkevIRliJzQGrc+kiItn/9+7V8MvrxPiQsDjQL3IJlmLqf
qe36/VjGdebjvygfXLym2CW4Q2z2k2tgy/wyGmr8tcHVw2BYihJ0aVLPDL4sk7xlrEnpD8ZyoGvo
NfejUy0d5Lkpmtv+ePPVOSGAfwacDolRPSU08ddF3MNh/CWXWg+ddF2pzoncAWKWNTIXoQ2n9uDh
Tewkw/VupVGLdkhtD2aWX42idsakafcpyAEejsxwHfg4HAUfDW+zCNRL0F9kl4MgChdyCIuvNzmr
GEDfuLbqrINOIrN2OFWH3i8K3/HkfY3LTyc5PAwH46llGQWDcdPOpEPRfvAkrhsfztYmxyxN45ii
M7l9cRUCq3XKvhqciXfsgZ+UW3VYlw14JpO2gB0NCzHtHQip/Bt+mMCofNxBsvJxgNcAUYD2K8/+
li0Lk58KPYlUYYzp800mNqfZA39PcUGV0mXuqqelVTCEj2y2yvkKpTI30FqfnZAoDLdJE7wpVr0f
mPOboCF0pKTNgsC1+o+a+rNhr58FqSaELimADaXvbVE95IFJcvhPAMfc+yBZDPoJetCWWvECkmxP
PmTte9UfDZtails5DHPf4rxViNxY/s43exNoXyKAuEDt4UcyHreLDgBkVPi2EAUPZbE7N9MwdaVV
4D3dieYOTwYEIqhgjCfdD3dbG0x8gs4A+liqmFAMWeqSZTxv5ZQTGWYmCLeOih28MN/MvjH1I/67
wtHwOk0lAKNpz6E9hUB2gvVcRQesRp7sJk6D3vTmZhrLb96/2I8wcOtab5e10RyF8Dq80t8US46g
e40BqsNSIkrPUqF9AC6Y/07X59pg57Qu6uMsuDrhSgcwFgHyDWmZOW73Iff38vgc69AFA2P0AvUY
xFckHIkAnzBXZo96qjFiaYcT7tmZKj0uggrO2ELu9Mk16OQotaZZob22VyRLEVVZ8c8nHfUSjpIU
hZY7sQVyh//eIlWyn9rPiDQogz+pFMrhHhdDpKIxaKf0wGuSMYKEcyOJIDBhxTxJO8Q6rF1U0RdF
PzIKxt0alM4Ya5sJoihezt09/tf4PFX+dURz4aUi7JNp3F15sKg6gs2qRJGBhP2hSwar5CwS516q
MkHwqjBJ2Rm2vEMHA8dbINv3oixo1BPEul2ffQoEZqDXHvDM8f5pzUrt/d0qdTXb2hptt2s6bwJn
kWALYcou+uL90GXlxjWdkIVeEK9jsa0eoLFIZq5TTSFNzxCqNDnG5SCCF84VszCsJDq6g8zriuht
85IdsZTBdYtF3VWe+E7cxRg/NlMooiJ1atbkR/Vb9s/lFG3K0ukEp18g/NU4hNLM/2XfVTZ6K6q1
b+eaNN/vW1JA7WVNx66q1DGuOqqRXPHULSukG8LYz6F7Lg9YB4WN0byoV6ZiXqCuSmCLUTotVT47
158yE/73TyPESNGRckn8+uWkRE45+BjansCJDO6t990Z2a1A4V4teZvXwE5HT7J9TfWgQ6hXnSUA
v04AsAoU9fcVv+jMMHlaxGh1np13Rb15SSf6mwnipiYDJi2MoS93Sk67mqnU7w9EeKv2F+66x85+
A7EwM6ugWPg4HYTR5XlX1GasqbehlxTt8c2kEGF4TGIahjYKw2qeAMp9dLmaS0pyVjoJoBs0HsR1
YrTKd5akUQ2EgUTtNkeZpz9E1oTfPoU89i9niky8YI7TOtjOxMYt0Giei9UQqTSf68uyUJWoe3vn
bVzON2ibSX9FG6sPWKU52LI2h+SQ5uApLR/Xlx0m0KDBEbhHkJUxGcGAjKJrRKmvZLEuKCYAXyZO
qccpztbSkFuKVSigKzCAvIkaf7X+bvKZ7lWStpe6H7wqT1hJzJOV8jGpR10IEB5S+Epf0SovHz+E
fzpoWhJcKmGnysmQ9/0e1oVDf68jzJ9z3ji05Ykv5Wly/P0V3+c4VaN6IPZuFQj8ZfDvlYoQduX9
9U7+VMJfeEG941IUsd4dvs2Tl0QG+FS+wuPcFTOz9I2EZ4nCYNdZSosFOWSviE1bUtl3gg3LZAwB
ltJ+me3z/+JlPaMGmE/3h0mGlrk+LrpOb6Rk1ffYUiPLAFPjyu2PhoiLH03BUV4q1YzQozSAkNJi
buGNJPDHLfQI2S46KO0S7z4y/fEwXr5tTnE9hnuRctfy7xKgotVYCogcy3nedGiTqCTAdK420w62
mhZV1tSK2POwxSYCV5W7GzD63uKXeCBAH7BWtKNxuNbOxqveyZ6DSmlAmQUAYZCHtWxluzwlWaJi
ZH+3A3V8cg+CPjR/Gu9Soc7nJBpAOIORhusVb14IL1cTGlz87dxAGFoe62PnOc8M/KcebpwT+rBB
VxI+u6OAjQFosGRPYK+5g80f3AfdfI4HngMYwTMEeReU6n8nP/EZkuUlkqnqasCG35UnmKIXpPNR
5re9xemryBJy5v4sr4bxovyqlenEJUyZGb/aOJQnhh8bm3ndjBK/VXY0Ad1BoKOeFub49Gx8evl9
u8N0V2KgKnvMPMeXX281U1g6XEGp6om5jnJZ+dTEX5qtpB2wxYNQaM3CSCLkRr8N44DMQFRZx/GB
iqNrZXpu99X/25q9IpJ3jT/Rt90ZakIQa7ECzG+DcPAme0hl48Sw/iSAiaX2wldGHEw1KMzlC1GT
u87QLCQ9PGNDDobaaMgO3NsC3GLumcxarMvJLERbWnok3BUs97lQDSxNpVEfzZYMHwCHqFVKfi/8
KmcR6fucT0wyAnWBmNBn9Va4GzWgsBjQAUUdgWA0QJ7A4LvvwrrkF79xI1WmN2eINUU45/SlUHJD
BtAx5k/k8sdsxfeH8fC2lmPdP0OJnv7AKXRnmMImzusoByxX3SfPS6VVaNTBjiF1vygtfNc+r3cD
J2hIkS3UN1LvETvKxrDCoGSsYtR/3gPsx3apvB4OtCt6iMcQeibcU2I9+QeDZqUpkcCjD4fDMbS6
uI3wqsSlFzNg5+FKlYQSJVZZtjhYyWED46KkR/7NhXtdswkD5YdqSpM9bqMyVbEkBJnBSwTwKr84
eeZluMsMRelSwrqjqfV/zp2axF0JslgtQP0uifMdpGF3gjD7oQH+Yx572ezHztTpASKn8LVpUGeh
2ttyEr7FV6JLnAqwntrAgI7zCH29ZSnXNNVUS+J+PX4Ne5P6NAQbWTuEsqVGhBqSgxTRZI4u+AGE
V4/R42ITjJsx4UItNXHxkfTrtjJr3wk81iGJ3pJ9dVX2kbqhM93WshSpdLpM3h46Z83wrnruUYwb
LT+Z9gRur1wv/w3NQ5IJOZGAlOCzt7t9Hg71mpXvxz+mmQ7pCuPpGPDtqIb8c+KiHZWQSwExuMDt
lNWtM9WhFIpmdDa0RG4LAseY/e46lBdDExKOMdhF8OAtn+7KaFLkJwkiQnKNa+XlvU5V1q+vct3n
DcJCwdp6eWhBs6dXptfDnk8FyelSiow6L5dOv+b5of8cZFhYjRt7HAd1x/FOEyP8RlJ7XpDLc8N3
q0n7VXrXQ1WQS6s3s4i9YlBfewvaJ0abQfHOY26ZrLamQhG4SmLjbDrke92Yuo42+3SrbwyANMQo
4RgH7w0oz2LOWB24cV6OfGR88hr7DkElkzjdLMsB8SDfmrjyE8HoNTj8GjnDDMhU2W6wri6bKAY6
OhFNUqGdvQLsq/KaItInf2XZe5EaU4eBnUkvDfd0uGSRK5O/jQRU4xDZJgu+uoKSSyY3BuMAPows
VRkmM3/5IlAc22YvQpVspy+rCa0wpg1J7KAwoGzTgTQ6yhe0xEauTRTIrH+34HaAlfwac/TIvdOo
5VLeMbW63ef9rSVVXqLt/SMLs72SGTTStsPR5wqjbtYioiEgV2hwIi3EiKLio3RJBvf8t3QmfjpS
YCMetuGn663vyMxYRqQyOfRRpA3Z7EdIxYMaXrThGWxDzuWpAra9C7HtPGjk7yyw0VrzWDebn1iK
+k3zHDxuFHfZBgXO8mq3Pf/AWaNPGMamqXDPV2wgGHUdLOZ+I+BiG0/xTONddRz0CGWiqFWSRZTh
PK0yXlZYw+GvV1ySDLXWSOO34+RJ5JTY05ail5aP+iuvHVerxr3JTShVYKhKcOIG/FiPOltJNqjj
YFl7dUpA1ZoH+Uq074mGcjLzOwVqkk0CGBIS6EGd+UIXrEZvaxn1olLoAZ4VW+hNONaqpPbGakAk
7l7mvhI9nRWu60x07bSES74GtnfxpJXI8BpGMIjNwQox9k4C+djGxYMUx5bfVTwpKJQzpzHXFs2U
bCkNj1C/rmmOupmIolKRsHZEaDrTGLl8dIdTcQajIEWIRc6veehVXGnONPG+4gG6LncY/Sw5WpZO
NX1L7PieoLk8lFqcXYFQ1XdQqcS717vE3CSzqEJbX68K0EsYYFGrp2wXbgTR+LWIqPIPaqhn1+VX
ujuSTK5bY9vVymSLKgJUa4UrWa6aF+hzJ7ZgEQLUV9YZSenlRSanW3n9H/E+4uXwsl2ZZ5owAumn
noF72JTjgW3R/9klSQ9AERu7RPWcHrSPCoflYUnvI2G7JZQi/rCLZGkHY7ke4G670yJOB1eOQ7Zj
SRw54Rccifo8EiRQNrO05QyD+hTlRmr7leOQeoNCImUHs5fhQD98xnVeO0f+7pQlMdnYNSly6thL
WTS+PTUyduwIVd+ydor823NINunjJrVhqPMaPirpdkeNqaC6OP8+8MnG9/Eu3MTbFEknFgG5CXu2
qDwyrcBtlKk32E8WOIEZ9XDSyIAD7h8+9eYKQHC8Y5z4W92w0aPTgTl5wG+9h6CfQiu/Xvngeyuu
/qdMsN/3RMV37U9N2lsUObl9FOTvllmgmSvmVHDFWA7SaVIZVwwW6GLss8ePYxDOxM3tGlymTef2
G/GTDq20k+8hxkFLcKqleN4bFdoUsr8xKTMupUvGePwiLb3CYhdFUoD5bjtCfgPhm1Y1OjQqdm6o
IgSG1+UBbvtVNo2LUgSQBXqmhlJCVynlA5eJpyQCZ1ixNnjsUizrWyE9pEk2TKVTqTcuW1ZpmhW9
eRZpYgj82lyRwr8N9CNdVA+rZ09EbpsgjRLfmEpDdbbm8ftvCvnd5/kPDa0IUG53eyWehKSGl7cc
HQv1IzrQcP6AQN5ovGqYngCoius0vhJ4ISh2aKQlQb6CwzN083v4yNTxYO023MLQpmwWIbt+cyVz
41iX5cLx/all3N+aRjjCBh529CpYkYccujHo56oZ6CDizNfbF6hdSIVSYVb7koIA6cfCPTJJ6LjI
vXyA+fEUGauXfInyP72ha6wcTr0a0AX3MyBPGF7h9uiBWuoHTwli/GWV+HgFSCxZY873tWQmOpg3
lKRd1WOBNCtOiTb6nqfXM0g6rtO/zMOqVcE9JFfW4BES6ccGJ6moDD7lgko7jHoJTw7mLH4Sx9IQ
JaHsxncQvWNVag11OfxLugx/GlzWa+5bVQ57ehiZafH39YdlYDvkemgvTTQjRIniomIAtht5kH/o
z7t2dKkYpLY6Py2Utcc3JFJAfIwkzEhao/Ky4kh8AAIfRncg0SzGjTV7osM3XTrJsYe3ox8Df1E8
MXRqLvvvwnACA2ttRDBzUEvBTyU87/FEDi21bzkH+RDu2ZdpasoVD5ms5yY4qpoeJIWwuuxuA3aJ
qIoTnyhcwB6hZh60jfFVwCBXxvEly+/SbjKjsYwAu2AI2lFDjPqnpBVuxMutXXZBYxSTrbGunbVm
YaCLJA8uh4uD+lr0w+LQd0gC4mFuGjDowsqsRdo1s8I3x5unEMxqkV9Y9F9VVh1yK/RAYTY12P26
+pA3rMCF9qvPJgjKpbYvnn61sVcvfHcpIBT/4xs7hC9UtlENCpdpVL7NaJd9HiTXqG2zdMDLheE5
ymx9SWBUoXOd4eQcb5OgcxMZLBf0lw6O4D5CscLbrG668oQtXYv2+uDkFqWUeIOSEgTRTeEDjUq2
R37OxEf3vLYhuywi37OS+cdD/HMdOXzfGdrqO8X+hRBJetr4tJP9FYQXn01bWRpOlOGEmPUfiLXe
R7HWFBkWczOr4Od9kcUB3vJFhD1jeZ1Cyp0z/DwfHmyXpeW5rgdSSCGmPiSkmzkl8zuE2U/dsWpU
AZ97+Bb8A30393c6MdZkJ7cSn/cDwRqHbYityWMvFWhYS/vvu9qcy52OvO4enVo4p7XsEJd20pD6
jxzRUQAEHdIOsjcO8KV5JeGPCFtJeOb1nMm2H7gvNrEVBXpBKmPm7WuEXXLIyYOe4tE93BSFNczT
alO5a6gJ+v31GrfRv5OaeNn3kswHvp/YYl1Gl3PgJ4C9BT4jJO4BKb/jdwjvapXg8+0+682V3a8Z
pjjyPAkOqpv1MqgcadNtD+OeRQy3Ojm3HzYzbVLMjZcejr43Z8laD5Z4l0euMYt+Z4XEzlLIs5Uz
giwEqjJeMBr7vifYS2juESkGXLLQcWqsHmJGjF3qCLww+imJizFwPMWuTOGL8Abka05228wx8oEq
gpmWg7YIwx0f2CHwMX6pnC29niSJcOwKPOpe9YHM5p4ZaeG4ePMwgkj+aOCXRX6tpIPlYzohsJmG
fDdH7EfpgtyhfgTSeo3xpasHVrUaipK02mHVOrdUlJIsDjE7CSr3yGsGQlOo+P92bexxWKTXQVbR
2ClrDCQsu49NiNfq6+3S3gUETMKwyQbflDrOkxdjsGN3GgVlnEDelFUz6xrS/bZBEtpzOnQTVpPS
Qo3dRfaDx8c5NEjCtEONpzOAZVBqaQnxQ50/owsY9Wm5LwYJuyIDoOb49tzn97on/Oj/Oele6c+x
k0jzqii4o9hBHFF/TORB0gbif8NoUnmRB56ezU8csKdBVwK3Geh62hiLvF59fNnnpceMTTYwydlV
QKn2Rqv5XHPx8rwInZDPIa2oBtbPtD/IeFXrZ8dLCM9iKeNk+4v5F5qOtuj1jWuMkxcIgOKcfsuA
aPAjVMH4s8JCxdJiV7Lto37aIh/nVR3j2G7FfMCR5ZVwoyxL78x9NMNC1x5d64GDKsDfio/h/1UJ
9ahkEApTLlSHJIAVcawle3j/AfsSHzdD4rIv5W2eQGYeBt63VQvfluelkfQrq3ozT8r6Nw0FXw2p
jfMTY4Adm0XvPiwi6Utz0r+DLCa6iVI654oHKFQxlRHUtyDgt0gBFJjxHGeqX2rURLzwtL+xQg2Q
eG01Ru/wKxokDize6vUhgUvSE1pVdA4nPEDhFSXzrXuZoRSVc8SoFd9BNvroUDWZYu+Sbd6n1owd
oQlVvM0sOpVuy/7T/Hp4UxFYxZGm1QSht0bRif18XtpHtKiOqjWxLU1YYlVI36B9gxlt57crSv/t
MLPLlDuz2oQPgHyS3BLr8ZUmafuMeNrugqjwaR3/sI4DlF2Ukf2JnjG/GAdGwlBcXjwEjhre9oI/
Zi3XPSsCUkVcO0XMi5GJEQ1ea5USg3vXyHad1O0qQtDV2PFOC9Tfe5ladPeOMT/kptgNnvXZd+mn
y56is70ww9LM/YUzN2S1kKZhQRodcv0sZNrxZbGTO2g2MnmOZB5Eyyz0kYTLzN77xjbKLRE1XDmy
kWJwe6rXRhaWMPKNC583o3o1XT1U5ap+ZDot2z99c1Jgbyl6amfCh43J131/8PU6npcpfpLZwEf3
4DMZOiX8x6m2haQfOi4Xpf/73Pfs5cClpwGuGezTuQqtVpNY+Z3ksB91qEtg63P+jureo27mTlg1
cK3ayWyXmSQdGUGgY9g+iiN4MVUdXzgkJq90xHdg/xilotxZ6DbbeSa8sgxg3jE2yTa+RuqWZ12B
aGeEwKr1a1z/iFx6BNK7yOeXwFzooAZLYjqg/tNbo6j2O2xiPAU+QuHwLKe6DnTC6MES0V4ykSq6
ZfOGCzb/f3IrcVVt2c6y3tO4Q7SE5WSlRTMB6Vh/vGLGl4u80jEKEeQ0MEiTfGd0k45+0TL3bPLv
g5HauWzXjiEPLmB8uQhSS2ApgDWznXvlkUakEtW9jcwvVvpgEtQLTxuqz7fcvJpwfcPmeD1ng6SY
I4hTz5yNzi4NlR1k3xk6HZXBPsiRaTDqYlXplyCbxr8cF9wWrKNGRcWdC7/dmCKHmwFVyNEGsy2b
VcMFhF0+CewmKoz6gRwWsZmv8mS7/joH23bK1xTBxtNDSWl4lbRkr1Yqjc6eBDrrLdttNhCUm/6l
q6dF972zVp3IofJemD1vGWV05p05OznHpY/z46ATw0sIilkpbQsQjq1cEpupJDva2kN3vtv1+J8S
gYN7kBH7nwofyYM3T5mMk4LKsyJkXlnQHnHnjfioZGYsvfIhDJ3h2EuBbU9BPupFhhqa8z3y9rKO
QFyEw6wuIZsjkJC0cWlf6U9BsbJb0SF3Dp09M6VGk9poDoOTEYqHC5RkJZ7dgx14Je3qRahVuayx
NO04mGnmmdP0v5kGwWWjUEvR+yKjow+1NgSW+iv75jzGhfJIq5Kao8Ly+Y9OKclG2p9EZUXLxwua
hp6DWjv45lTHvNVYv2mVF5khAMoAAsCXMl7KRSHVQMMV0vuoi3paG+rb5im5gzOFElrMZEZT+Q9/
EuiwiigkX4vjmZAqcDv+2GRNJ110gUKCgPhHHMJHxpWT6/P1yYJ/EcOF37Wx3Tl5GVfEt0PhdS72
xMdgefXmrUdPn/37YqCtKWO5PHRHM1rgyDRQIWeFd0zMlSsnwU/FXvwej4riR269qjZdWlNqVYkX
76EaJqBalfohGpHYBKvVfmsRDKdMwdReTObTi88N+mT/HVhNHkc8rpK4FqGdRlUamIWw5FLXjaJ1
iMMsla9LOVlbUnQo8RX/e6V9pHyC+hvsrSyZY5XEK9DHzeFxC4t2wxPkqBiIL/mWWTIPiRDnyfTq
hYjPPVQyTBhAuQKLX6ruaRvL50sAshlO3w9k/dqWCfRHWcf1RaNjVIl5V4gofbQacX9ejkFZpNP6
xi0uG9+qG+BYeTN42LhpqMA4lrWxNCKQ2nZ1jp+Hr6VQIDX8ns13jsTz4VDtGUmnwaxPQ2DgpoJl
FfKOl3udEf8glNg1QHUbB8sxnf05B3x5ScxIoCoZ/SMG59mq9HsHVDTQKgju/eIMhIVWQVHr/pWH
KBLRrOcMsbuDbEt2MwS9W3hsLy/r6qGa4X3p9cUubgG16JZkiT9Nkrkx6HXnwt2cr0czdaqnYO+s
2JEtp0S9mJ1+gQE85G+gQB6Deh7gv/d6QbvyCvTnT2ranXNubZQIU3Opdzga4PeBR/sMrhfKTZVX
HCk3iC8KLRz5V1dhzVyycQ+8j66gYmTma8O0PCiFhTlGH2Xqn8+vm0lsSv46XOFEswJSchmnqw9a
cJ+O8sM6482O9hI5XxXYljgF8li0Jz0kfoMDpfZk9LXYhDVihOBbvuDWN5vr4W2zFIzRISdRrVTF
1J5YqGhO3UigghVhMP42Ja3iihlvHvR489Nqc/66RBtTXhftTtIPF0hVk9pCVOUeYtMlL7L3y3nB
04+AGBkAGaZ4gvyp42z5ad8IAZkOCqzbSsqiNvBTI/R3KBx9EPhYzLhvV/nt5kbZSWlN7BxsowDP
X3axHx2hT7g/O6X/MfoAeVHVghM+VNzQfN8Ay21vo28WGle7+ts9ygQ6llIzU+ktH8vXg/wglzx1
LqS0mjJYCN1pbAfQgGykNtr2GNCxtLAxlOS9ydwu1CWtWpNRkkAAbeCkaDt1h4yVkJUCFYphfLae
WWGWwj0B2sh0crO9HH1irO2VzQPTHOtMtAJ4tLS3vm1tiRuBx9ymJ1Awja++8rS/Xrk1yFE1Fcq9
BEK+VQIEzxIrkGY8ShulP3Vcvn7kcxIYyjt7qC+OIXmYBZcGgi5yt3IzgTO9ngxb85qs3y9ZJqgZ
ElBIMx3NJtELOWiSxzviCOcU7jbNs2dDSaaJqzDUtZcLuP9Hw3z65woN8sV/6nKblB9P1WNpLH7F
6cSlpkfpsSS5hGpGWpvmqq6EC3gleCGyVEJAticY9XWFJjuX6Leqd5D+1C7SPzJv6ogKgg4pSjpM
hQBvcTLQ0thsuaUEiC3DsVF3ppSoJ6AdJmnwlmILx81xknUb9+Qh7r7ZSJsERH85yHK6kSk1wVnB
P8hv4bLCSHPfRsGzPwxpcqNZF/bzbQcg8RLydj0yNFU2HYnO5zEShHzPX27JJitWnmxKmhwps6tB
rtBO5Yu36dWNKEUl3g7e/SK3QWOzs4x7WZ5mvI1yxFNP63KTZpu8Ix16oRTkI+pwNFV2R9l2GqXR
SskOzJPIMasevalL5mcoLYkp0zFuGv7tEwnXrnKrplvPicVO3zgUuAlHStHhxYPTY4ZvfL0nuRUa
+s+vp6yL1qYsa7FUCubFcUtKY3Hm5b2V7VdEYX3uN+gE8tL1rR635Q1x6pcTrudtxBC+b/85yNMM
v4ax2PPMMGXDdVaysjw1P1JGHmIdBADniybApX0XSwPE4E8V67fbHp5PRzQt3LP0Wn9Nq1PyYXqR
JA0kQpy4wVN4h+fPCFh9KDgniwfM+4l1sgVnlOfMoAy4dW61qNS8ZYbuE7wICZqe10tA5YA7E4ML
gtgOrbP+s0M3qUI1ccb/ynfOgDsaaa/GbX4QVDGwZ4wkOzlOBczaBSh2NkNlXCB6LbBww4vFdWJB
f5hn6GWOTpsvtMuc7BljpQ1s9i6nqcTR2Qjjmhey9hrBMcSeTeKYMp0eJgyeISGKlYcXEsn5J1sl
znOcwGkAqkyXFRXwCCqaxZKrsqmbjZZD0H7jkHnqnu+ltXdXizKineyBrl8mlXk9ct+b9uQGGOD5
A78cm7MidBts2CEN92EVIav+gy1WhXixb0qKi18akk3N5d2/gi/pxdBRh3EBfBw4Ln4i8e9vQFeL
CIpBPQZvn9dTtlzAOyGZj6vTB45z0Yzc9kIDPrHR2Wusv/UXnNV/W0aZHvNBxEMuPrte9r3vLzBh
xAPXrl3dAGgEXgmYmJKVU3+oSFQP631gpkWMfvHQ1v1IbCZk1yz5ubEVD57Rw/SIqQOMF3qwp7BY
6LtFV+7Q96YM2UTOMdwc0FSTJK+xUKsA2R0M20pL05MBxvymlevpNcmQjReGVlPeq039EWpDNj6n
ALK7zXv9J0Egcoeu8NXaLhmAyQb8tIIGhg1NGKH278ou1PDswOChZisJjKX5aS6ow6p9l7pHrq3a
FzDpSATpGwaH61hblTPDe41bvGQJtB+EQyuVKx7J6eohEu1yLXGUOqXDejHUUMdpb0H5MbwciX+1
rah356nc6VcGDYNTi3Vy6LhT/yMuCQSCsrxwOa7W31IxsEnkvbCfDLrHlcYEVYEZIR8HoqBbAFWB
jzVaZhAp4YCee2D4fcafUz3F2pMb2/TvaxqC7COleGzOQ0duw7mfK+d/rQijR1FlJ03wAzDNYgDx
G/fdBz7/geBaXFalNacKMZpbCATDLBhu73Peh58dzmMjo9GabTmbVJvLkUXFPKTOPdJyzpvcCpWN
epYNZNZuOrS0k4YTSIhmGlPhEFt5+e8RtoAzTN5ja8UExzJ2PiGrI0lSvRcC6sqsFw3tmtFCKf+8
v/r/letKSv99otGWixEmv1d8ckfjT/BNnqHEApwaczyenNn7UaS+bJT8ZsR4ED8r9SiFODedkBSV
t+aHq9g2E2E6WhqvPD7a2LEr01IKBrTZ0KnRAmjQErXnx/RtNgkxvrn2f9bXP2AldTbG1f0ohVhd
RvqgcMH3M/jvQ4owngnqCKC5wFiHUk/sXPPtOhemX+S03HeI9oN++lAacb+dRm2EKTDG8fwu/3vn
CNCdUmm8dH0diB4/vST8w5GhTdg63+DDifmXZWaL3ao16t6OKnrGzanUzrQNPfpLPoe3yTDYwNn2
UOf0s+7KJ83DR856+C0TewP5jdFHrgx67vhNBL6eKc9wfUe42YKjwTZoqEftjLb5Vaz3viE2rz4U
HlAGKPXZraK0KI3fcxxBacPqqhmUT5T9Y7vDppGSHxPlAHiIdSkqg4sWIYVxBeCjH5V/G6TAmHIq
ZRzfG5TpoHTQ56PiHoS6wdDakOid/K0wYxK2HfCd4zAiO5e1VeGfZMBgB9mN+6ugyILx4QEAEMkU
RXdZ0rB3g745vDAbb3PtbmDidwblHamxW5zTOHx5op7HBrdsozcBZFV6hL5KJQulmUjv1QZrTW6R
t3l07r+UQPWtE6fAS3eJ/yCl2lwwHdBmr0/fvpjJI4EMEmxCiuyFGWA7D7akbNZ4BjFZ2yL9GQBN
C9LihbnyvqYAxrclK4CWWterQZv83sNjpaZBSZU7VWAFV+fYI6FzNvzMgD63KveBXW47GNxN1FL6
4wzBivTaICZ1ubXcY0mRSfcPLO6yAPuNllEgAWyaxhgZGuktohoG3CQtcs2Rk2X0bIHCPwz1RM2o
FJuK+ANOlaYWAVGljrjRF4domb2k2s0rjAMC6DvYsvZycHsimDXYQLK1LE5l74IhFGIUIBJ6rXnF
p3hBjYVJVIf9fB8lXB0foZFi1sQgvRyOjfuD92OyiiYfUjBaLqPzNOYjydtvefDuJNaPe2GNLGve
2Jj2LdRdFtXvCo2pR37BayDHkGNhG4oIi55iU1BQwh1qSbEQTEoUeoYvSXxMKaWg0yX5DSfim9zJ
uf2qRh5vDtg2B+1+6qqtwY79sKcNNep6GQ9CJsWqvcRO3k9Pur/G6laH6UQB7xCHilbmG34WliSN
39kyP0bx/Ji2AsQzNBDWrVTOOtKDvLX1gtA+0xr1ububDsMS6tzv7GqmQu0QvrHnTYjGZ0vDh87F
g3ALPW+ewC1cfKppfMZUFnWzERZ4vLpcFAZei+dMIoo5/NsWy8w6qi+DdUlYZoPIOuFziZS+ES/w
VkoUVCvj5/iNyh48Lk5ZwDEJJIDO8cJYrei+36U2+hou6+Q2qNJ9iLkxeJDe2gCSkdUgjkGENRpO
+NbCDitI7V82r6u1ayYRxXspgIIDmEo9copnb7pybMsrdKD3q5k8LVXPTPSGIrS/19Yr2b0csSrc
rT3JVQn1Y16HhIlrzkzEDg+odvVUGc8fJkrK/FvweawoVp+TNbHmQPWfb4kr5A7ao+KADWATF6Kz
MuzBEkiQOiDm5B3ovRRUlnKUv0Gwo3I/p4zdwzRXTtgZs9WNQCBKm+FrKhrqtFTsMe+QAAcauzwr
xOMRY0XC0T7xDkTrDm4BV9SXD4HEBGnHCF/k0ReoSi9JiYWBwwM/6bS4lFK3JlW6qRK+IoCDkWdO
pF1LgODL7G+Z1t/DMSV4N9UtenxsvfTVnjmyvumBKNjYnHW+ph5fdiz1PXg1XUt44QGJVQ3QEeDD
Bb5zHOV9W2BjZw+zz5+M7U8slnWhTw+awSmfLoQyHOhO1e0g8V4qUOTJ0n09bbsvuMAdwj3wM0Ie
sT72I8E5nEq/tkZ79jL2JdOZZnNIzYLOJwDzLRdpKn/tW7Txo1RuwpFYAK5Vieqh13nkDDbJdaAB
KWzcZkGoeTKXgVEXmm2/NUa6ZqgyBwwfZMxpJQDkjqa6fTRj6JT02xTCpo53RXfUPKEb1HSbP/A0
FfBNbz4WGzZuM39lVQpGpFzkNbQE9gG0oxAgVHWES7CJDTFnVxqy/aqDK0IZeRkubk30Zr5XdJoo
WgheP3GkKviotElRnKu4WXHnHZeRMu+R7Qvw3KUTgVoUsE7FvxJF4owGx8+15RXZyg0x/Gr5i9AU
V26GR2npWFUs6ErvuRLqSjSqN96pVjsOM7v+0udh1Hg5fmxGz1XtYv+FVoSshrcL+8XJIF402+eH
wLIjcZNQIq2E3fBR+guAxdvZo9awcXWN5+BQHOzthjv7t942IJAwfT74bTijwdcglXgLxHG5w1Uq
NsokuJCokjKrhF4eNrxNTt8M4n+Gd6sIRLqrx1m+pCTJCXrAzNNEbFSXj1Kxj22TS+G3Kjuu/At9
Xug1cqkML9CwGbt+FRpmvKtrcOFa+mVc9SHLYH51uBW/1Bpryhl4mAzUuWKuCVSI4FE34nNWR0sH
2QDX50oZxEB13epxT5/FNZfO1sYRdLSwKwXltomy2CAiJ5PAfILPwWrQrdq59YXPZDfEDQFbmwuc
60Oi+H99zX3Axk6nZiTB56aU7orw5RkJLruinG/HFv67FLfDDumBd7ZHLxrfKODfmXOAa66GnAys
gCFTGZV+XB+defQfn7Dt0jLfXrvgup259rFR9xuQDy+TE7/AY7rv7gFHf8V6Xc8xSo1Jdp/UsB2G
emAkayvySt66DVHDjCNehxm0h6PB7PhDtEvGb8SGfz6i2kkp0SNgC8nZQ2XEfGzsubNLfpw0Bbw+
1vcW9jt2iN/IvwjtUPC/Vc6DNwF2DIvuQr/QKLxukGqPnciCEZPp9YE2VIHS8DpIMAcfrf6QZ6m2
/P/Lh272lnROe95Q4eYXR9doA/FLsIFmJZY8sXy1M8rCx1ZFp06Jq5ScY3JrYJIXWNWcqcSS/D2E
PUB+N5S9LsD/m32GXMUqS2ExiplN+Np2Qu85Wd0kDL+Z7imZzC9iOAPucrO+K3ltTc1WiP3k8Fy6
VR/goJQPmvqn/MdalNNzLYbS34sYm8u7h3ciLbdK4kcG6awB9MLuiieGTMCGxuzl/fmAKYvRVb79
EhQ6INwKGCE9ajkLf5G2PnteQ5AIdQGqi+JYU+yTjbrk2oGMv173zUIeiONjMs2iuXf4qvoun4Vk
+DZkb+nbLjpgyWySnopxyOVw7Nz3tZ0CoZ9vH5X+hjSlryex3HgKeukOFpflI7ygH+xnuNRlFz4w
bPEcbgmlCdhs6R4OyQmEVjI4JfCVANjda3KOqR5jE5qcxs1hrZNJNkKLRAwdC6hlZ3RfoFI7DXO0
bNGlTpqGq4iWUPMQCAV2MzOfKoAIzCZiAUO86ReJ43JG4u9Up33kARDPG5s596jiskjWAbba0Svb
s/Oh0tT+9X5kMbKkX5CM/rrFlRrA4dBctfW8M06VaMEdNUVoEySuf8B+VzAR1T6yb9AKaw0FW+ik
XmglLaExggq9H3y3vicFy6hH+0jx2Dmb3uBkH+NNULP8bqcUGA/EglNDlaGT+fLkVFhCZuMpDtZ3
11mZeevtbmagPUL/+ajq7JCeshtnw780r2JOEojAKeUVVNNk1pSl28VCtef1OYAwIFRLqpfbEFtu
8/gLOpo2x072w8ThzR8VrTX91XtJ0iQPndr7xRFSixV7Sdh/s/8sFRbDhk6YMnnNWxJBvxCGgE+N
PSr7vOQtHbg7fkYOFl2tJ3yUQ6jjrtb+YlMvnHuDEvngX4cOI3xKWzo+0jInqvK/E2ZI+1ZF6OAh
kadq0lF5H5f6PVD2uNxFIcZOHh2KZMCQbb0SfL0rOKFp+Lk7jkBrUnl+VezXMWw8bTABzq+/8fV/
WG5zsjq/eytc+SHudkK4DIBypdqyqbZXElPZBZkNIS09gswOs5gdhzGOoLqncWBqNYSNyNsCTqIz
4qoYonm3cO1aHAcpl86dGT1Uh8e3ZF2eiImxezAYkuzxCWSvSqVRfN5dzVMplbOUPL974h1/MMwt
v/MgRDv+KMAm59qIqTgCwELWIQrwg8fiNOiiX5jJtIlVDgUtEWXRPu+NEfmXqHtqs8jyZLWTLnhu
AMpH4osvDlvIlBV3BisdVcq8R1f7idMDMsZ6v9AHQswN/i08pv2ys953sCA/O1rdWjivDczdq/xC
EKtsXAEtbUhjpRnWzjzYft0MZ4E85j5DDq3JxgSEtyC3zXmNGXq3d+/riHBILpNCmlgmJdwML1Qk
zUzOwiOmW+IgGgJlndisUiicQYBMgPYsbsTVz8nSgr7SDjjcG+8HX+dtOCSHFtPdguZMRL1I/Jm+
5Vqeb6DDJprZ778uP7Ct9XY5c4vod0l0FBOkG16Q2JPNavdQetcjaLW/4LLBn0l5uKtWRbXdyAZ7
QpHMyW15vyGrjmCx9SzBfqU9X5H62HLlMWEhcfFCxxykL/RbO7jSSmgaWNyYeRf+hIvMN034BQfl
1OHy3XXg3dKITeFwkdVmt2ZKQ0LwF00E4+TGC2ppS/8pvkmqmmESroht3gVvPsERnatxxq9WAU8X
7JNARtsJZ6aaUUIvSoO+HAsl8WdjcTiife2vETcz9ZfaEPx6QfA5fzkFcywZWuzv0CcJUFphHnt9
ohqeKaSdH3KHeB5ed+NKl2DiLsEKf7PeFmQPK6hfsY4659WCb++J6UGI7xCJUF1UdGekb4vVA6ot
FRPJYCTblL+eLDgNP9lJ3yRFpCZyzYXiRr6nUQGIbSNC4Gh+bWWI1h/klOTSqDrI+J/PGUWTSp2Y
vtjDxaOhjY+M6KUIhC4KOFTJqPLiNduUa67YuHFiOQEXO/wwsrWhyh0HCAhFXXhQGfGTRU7awBDN
pevw66cBtuMMO2qQjN4v74ouJ0bsQ5wT3KSQZR5B9YzRuU8e0j/yMwcYE0MrdURPC9b/KxbeuIx0
76Bdy5zmgLft/efZfEunEaQkIdba7rmpjBufYx2xZ9eVLml3X4P/WQzssXc6xOoHSBDr4L4dPt+s
sguPmSzcG8xG4DRRYwKimpE3/dr1gn6n9edAI7CK/4hMvy1h3dKyl3dJ6PBAas6gm0UFlPqbJNH/
XloY2vbhtEZWEBXEsoiLCg/m3K52Gaqmz9++4Twll4ksuub7cJPohUCAWwPNGcZjyxwSvX9O/lI5
B1xdBdoORYwxXNLBZVQkULGeYXw68kA1Q8FXRmtpli4JFnd5r05HmuNlCa5kwVquOCDYbIOjOwJo
v96PuF1/K1eGCXcI6d7SP4pssRgW5aVCRmQfaVsGC8bySwgK1xHrzNGKGE2TbITswj6nk/5OxdIV
rVTZWb/XQHJrI0GqYuewbWsoV0WrClNII29m8MUuJPI8AGUbcyeG5nZhOHe6msK4EpOmjIEE8aVx
DMiuS0d5tUHMH/Kb9WRPzWILKe2fyUkrQteRC3fRiZQ7iNp6+pYZnh68BA8j+QT3t7b9MiYN1EKk
LNv7vLA/ostd3KoPAUjd9xia1SbRViHKHNhdBj1xTRck+bYOlzhojGGDzz7CSp4XKtRlF3e5xz25
lnmU5qo79T3sqeWY+Hlw/tWGi6qru147KuK6WyZ4stE0b7+Z7cvXaF0V5SRTpVIKp+EIP4ZuqGG0
WhwLdEnTK+EoX+jlIaBf6jLaQFlezy3EBJpM/UOEeWgr1198udttm6yB6jgzyeScUfpnhvRtqCyc
Ymyt+zoXnOImZMJSfTzjwby28ZZWhx7udpk85n3fkWQpYZDNuih6zppmrGmX01+rNLdIVkFVM3bp
vp5GviHUic22Qnxnt7U5QOavuZ8mSe9AGJXJ/6PiZNNmLIFi3e+eHdfJC1t5nNVo04ttwexQDZSA
AC+iePbq+ifm8JEeT7Du+hlbt5lm28yCBfDffzDCYQQYfH1WxinVYp1oareIGk63Sbqm2r07V01l
rzmxjj/P3sF7cBzGdGIOpp6BcGx0IMJOK3y+dqkTL0frX4W1TxwNlpvtUdkO57GTKNtadoSf/LeQ
NsteacpNiiC7Djm7+AM1Gfd6KRr880RzwQHpQkf89DSr4GMZEu1IEN+4pMC3osqYQjrvU8MgE9ic
pf7lCUOeKd7a1qyolaGjUfVgkJ5E70VuZGXolBbHZhuub6YXRIsrqZxM9KFeOnUUyQWNTsgZZulO
dTx2vLo4j3iNH1/RpRKIJE2o+WBlpqlEpMdiVwNkpxsrLSXyDXfvTWDtUsR7b3VlkySVeo8GiEZE
h9vkJHDfc1O4M/mBpqdl1L91ag+ARVE6USJFtV3iFDre7O3YVLkC4JdmDdD3CQ2N0Qd6UbVwgmTj
hxPlUOjrD1ozGbIbsnPKNWbhlBgKeC/fNJZ6YsPe4kvZgD08pUuh+YABLXET01Gkn9awTddhFiV0
Yt7lMT0kuLHtH3Z1rDRa9KwpK/vue2gEWf9ErzjobrgjQ5HV8KuBOzaFRK6QVdIpf7+HHmUKtSk0
UP2CwZ+SP69elqu6smqUw3sFOHc70myyvmH5zpD1MMbxMTNYFkM/JjTt1e7EJBlBptYXnVvarwAq
qGZx55442+nxxb8vsejYOi5kiRBO+4as6q4urXkuSOaChIXmopXblXIjGpwBRD7L3rmC3SEiqoLW
etziM6kfjFriHbng2I6q5MNEW2+wUBpw4bgm7Hc+P2AIALdSrhj3Ucff8/RSBlAd2/DBlRBXo++I
OkLwMO0HtJMs8j7RdBXfgyGHwDf+TkvZot+2a4sw5VcJM7mcIvzGn/V1Rq/SeBAmy3Wy2MlYIrVy
GhBP05+IiC4oUzmQZi4BtPdWhTf+Xl/+fTC0d0utp6vrgecbsKiGjJf6OaBqY94z81vau8SiYVpZ
NtZATtvKR9rjkk17hi+hxXEynHG5c7nmZosjj3xxLiAyY/V4vkBf40c/4t5M2i34kKhneVPirbIv
Rqd3v9AurZTtgS1NCIZRKKjEqXASB5pM0AevREkHgaDbetO1OpqfyYQOegpGjoisJLVp1sUVuZk1
ZuLZjaimU5GhvIRryiRZw/KHYCWSy6sSJC8vFxt1GZUUyFai9o0OxG8wGcsKG4wRWoo9O0Qrxoh6
yaPLMCQowkG5r9dJRFqZCQdU08ohzntAQn998FRzPPbZOoLF2ncHWHMdjIsWJZJQvdbi1lgYd8u2
EgHcjZzfcSU0hUTOC1h+rNCBPtKUmcVVAhq/ziMhhEZ7vDf0HfAN7eRLUB/opX17kyrp1YDj3Zhw
jZJLWjWgSiRt+S8x33TPN/8Gm06tk1ng9+uj7GqxxNtZ3jkg8ilhVOkIBc/okLKLLDdXXc69Emk5
gHb1N6FBROLRIflpqIloaOlPj6t0iPCnLGdGsWj52z1K/hmzVN/iS/GVM5SDYAPnylEPFcT+fnqV
GYxy4NZOyORrOAGDBfwZfiSI2gyWUyD0zwfRtkQIYeZ0u7Auq8MIkPSSqqu0ZEQwt2M9slSvIdZ0
zKeCn/cVFBl+Cx/PXhjMx8Ag1nI5nluf2VTlvFSTz8uB5Phoo0T+ei2ksa998ZWgsJstS7vnIuAA
oxn108U1LR0Wk5aH/2gUib99m2A2AYkjSH1dPWcRelKIe8RJ6umdfAIhr+NhRu4oFsYpkXJRGlkF
LXc+jSCGAWL5A1yXc4ZjyoprGZXh5CtWiqqTRdsq1AJU1AcVbAkySKUmcd+AzHJ/7ylaJDeL6GJ7
pW3pyLO21y8QQk+QmTQOU82FDj6qfvBAlAVFiPHDYt6lPNaYRrQioVK0izBdaPdJRwiUPqObmU3n
FcemQ0I2HQFbn0/vo37d4CCMdgdDJo+mXtBSDKSxTXwYuM6iFEKDAA94qKFcXVQdba+yjmYZkIsL
Aj+sLB+IdDTXFhgBsD1QcH/w+nRPvnVUmQfSaDKrFpKlVY6Y4RlWL8Kk8UZgzjpYm542mZ8VlD8m
VlMIHNE8mgPn4u9KfZItRf1Mw7Z3Cm/ZL0IRei3s7jbSeIUs8uCILTNv6ScjUGdxV5I8r92EqAxL
zsSP9bFbdTHbOtV+qroGyByuHVzyLbdsaCgHMuZqYTeXuLb9Jn9SaFw5UZZLYUPOz5m55Syl8Rxo
wMi1QM/nfqD95zcLIoSf8q0USNPiyqjqOmEINX7SnfAzlv4rwgPwaFiGzqFTt9/adLow7wtRe1kg
O1oCs0dJblkR1S4td2lrND6M+awDDQkzyPRYMrwoFFW20O4n17C7oYfO21T7fBeOHCqGF3O/lbX3
IQZvTSxd18YoYhTlFZbMH63MCaWkyTtihSwzLurDUW37acd0qrYAowKQg8jA3gTCVCmgeykIc/jS
wS5swjvYIoX6giaWGBpKxoC74otbwn7y7q8gNmNt+UScyY100HAcOc0B01BA1pBmStWW6tnL85HZ
XdbLJKDp2hTBmDiT27VF3s5xjGu5g0Ow2/kkA3muI2nnfgXcHuDwZAAMZgcXsVYXUNTO/cYh1G7h
7jrhOICFrjcjakV6UnNsZX6qucWV93IKhHx6Y9QOh8WTx8mWp4a5ZkkWd8wkSkyPbpyc8miZEDLF
AmUmCALUxBmN0/L7dhAJvtX5cn2rHWGOu9m1wn3b+dHyR4UxL9c49ibL4sS05ot6Xdrm0Ojq++u/
aUfq7foq4yVzjP/4NwAOWxoDLDl9oUn/2g3gX5EZR6/JuOxC9yJjTpZwl8h0QqOzdZqMYnU2Jbqj
Z14TpNUtQx+Sygzu5R4aJ61grGMExZRcrQzPWmvNbtvUZ9Rcz62+hQHzdS1AzlHrXe2VnAwYFZQV
+XRx3PXPqQM7rBmIBF9H40RSQw3MfjQwieZdvoSjL2sxrStQx/R2BAeVnaIOx8P/9rETkEvtsqOf
DnxTYZBkYlYRHQNhwkfkPAykg5OmSsa2QsiClw52qCjM1D0FDRBB1H1uBbkQa4mVQU+/JPATt548
LGHLpAA2+86EFE3SnS4o+eqQ24HX4J7g5B41paUoQ6D75CEvRpBNYZGDmOGnzQBr7YDG49pJkwpL
CzmGZIOPtl9WVZEbWp6Ib6hYi0BHjkyS2KIrZE2INt8yQyfPKT6fkIL8W04PF5HMHdJ6qRJPGtq2
CJarW7t0C9UsmjEupfXXLIjf59GSQrUVzHGzRMwii6rd9D3ieSVLPF5vY70qxtftx2839m5gdLB3
ajctypW4+6YlvjlF2lyKZ6dGFP/4i58fvJKln4fFAufQ4dkrHHr+CJoI9LKqa+vt17Tyi7MOodKK
CWO6pXrSvKLNffSt73Wjr0ps9dLWEqd4X0YNYFH3//M3vV5eWti2bn2tb54zJIpbXRjElHuL5KK6
Uubj3esCKAznykMjoFgCF7HHNHvru5tfYnb9D5XUoyjRB2TpJHaUUhTWDndkG+a89c/79weJiKjY
BdF5+go7hKcdE7dgvqFYytcJiXkIMGC9h+hE2Xk+n+t3B5b8c6Ffr/lFoGwDpR88dlxqm6MV3+Km
c7zh5v6tE2Ewc3ZS8+WSMtRfROWsKqIobYmDR4FeY83zLtpTwmxf0ld3iPo+QVuz1xP5LDQQq/MZ
8kyYGbQnJBo2pGErXcHdO2pQN5ZzZuLEzGErf6jUxELKhYm5iPpJEMSL4APOLhSGeNauHpPFxcEB
2JEXV6EzKFEandlZ32Dz6YJzfg3oek8qTWudsexoa8om9jYoNl0FTC+D5VvbFyPlmLcy+nQ6iCf4
Xifzs7VkU9ES0lBpLyqI4Dr6+4HrrNCtfxyML+O1h8HwHI1Ql8d9A8YT3EBcYI4pBbjsI+gjfJUU
FFnS9jfoA50T28AWyVYnTNtDaayPDcbzgfKeLPD1P7VEXDbgtfsaoC1LZLh/n4AvsAFKf3J2C6em
OZKekrPwgg7Ztjr1XEHP5BxA0leriqvpWkjT41drP7u0fgiJ2622xIO0WeAYC7dgwPhUY2cTkdLI
86S8PtH9yWeJ188Y4sYlboRcIrDs7aYYnpjpEX4KWGbkbZ7RoDFVPC5tbnJVY1wHGBJrs+iMeXbi
+to9X5DRWIs0v7V9ftSOvzJNwHpTZsBZzzubRdsE4r3JjoAhTqpyg7ouWYTk7+pu0tjjFs1erdrT
vhFsZpd6K4jpmc4TKcS2wOdld0CsPckra1s1npDg3+WVJhduEEf8Wazlh47fJYc9EHgGfNeSmlbD
Ht3OwYz/k+3SIfI8AK685KafJ6qCpd6n/hBSMGWcSKmj3gzVddLWWIlKZ+8w1eUzHm7zMFfFJZeq
n5VoXtd+bHlBRf9TabflfyaS3WviLTSofQuywEjyV0Y2HlBwvFOztZEPt11wthgUrwGGEPptilQp
p4ouXsGvcROv07ZqSC9cBpivzbXoMa8ujfrxDPwMSrCxCWa/Y5DiYtWvsWzjxH5mM1UL+s/Xdyhr
eMrL00XUawUlvnarTiSiD+mTTPvhr1gbtRLYQSvrLWQ2GzGKApBHU1Ht9JGWr2SFYRveHmPfDMMI
sL1LZWKASPWMvE3BOKI1NB8Eq/yw+C8fDzY0BYrFiTVcvFz759OhBFBoTdsD+rujLp7KgyeMva8M
T15BFOtF268Y4RRVYfgUTNg/o1fv/0+7OxS1QQpdQUjO0BTuwKV9IxWSRES/QlFMrOiJAv9nlwqw
lzMt+pUmva8LveshhLhkWjn0vylDWPls2unmpCHHX5EyZ6Bc8r1HWLdATVaANo8gsqewe01BQxiF
97iWouEncIDr2wiwvbBOXX2FJb28Hae28UjIGWgwHrdI2yPrwJ+EgTFtAl8d78U475rXzAqCz874
pAEucNzwttoofkwu9jA9MufjuSydSs88BgCRSCJVcWTP+pbRyb9Rt6LeSuSEJH5cvOTgwEQfxXLb
dYdSDa0CjyG/hW2swuASVVmCQqk2Kd6jM6nK1wdme0P8UNmh326MOWt+k8DrxvP+AVJJfrEJO/AI
HL14X8dS1iKDiQ6dV6Y1/IwPNPnE/b5iDzjW4hwTKruvpVTtoVfiSYOku94sP7q/bA1GFjJlTZeW
D1SxzhV1XC4kdPc3mXH4qbGvHn0WyoLV6AbDgB3TXS50zwsVc6vfp3EY8c8knSz+IcfpauPJVVY8
lUM5364vps3zNqPRSg4bw8ljAZZEkXJadgo5qfKSha/7+aJV9wEbsi3Aj2x2lR0bgRiL5uu0MkN0
t7USHu9iJKPQChX3BSjCyQaatu7Rew+PInqU6DwY+RloMCNx879e2Uv/3i3OcVmXyXhcVvsMhX6s
Nne0umJ+Dyguoe/xuKXXJY4+Ivi22xbJ5h+zjlEAMYyCx4f/Jzn7yKzmbTm1ASqIKGMUXDaUnGRI
aP3qc0BoQweivDvMhL+8XrO7Zxqffnebs4T0SeMYFYpUb57j7YaqN3le33vDxVR+NjOfedcOVQEe
96wo24EM21iOqVbAaKi+VGNLc6dI/FSX5PHBYTdxd5ZJ/CycCJJhfSBpOpFo9B9z0p2q3R/n9wI7
szrx6xKJqNdekmIyyv902tweCi7v0OJq7UAHEx2LjCunoQU9az2Mio2stSSvIdnY4nnH4t9CS5Zg
cHv5jzeCciHbiEvZRP+svjHMYMEQhrFJwxMrs3KDu7H67esl1i9EYBgnPxswAfgrdRDbg3+D/u61
1rHRUdeGC7s5j/RXdonEdtD8qc1U48LjYDVvlIg1eOjX19ws/Fka0RbGZn5dRYLbZOc2NMfwJSBU
JO92R6n9Uuh7yqTepMtEmZo7cMc7UN9EC0waERlcIRvnooh5scgIlxdopsQV/z00V4rFsdCu9ZXZ
9y73UFc/tyPCb4p6qZTh61h7GvNFeS0yfaHOWu9QElrmFDQucATiQG2XlAXTi6Jbl42G1eU1cg8i
14MAn8KYGDFskHRK2BvuqIBEOzJHsf41otOpKahamrmoCaX0WjWteigxGnPaUcbQ4AaTdy5eOTl2
ogN8ZOfi4QlXqtHcXA1wlOFyeCrw3CbNnKMplnHwrd+Wud47FFr2n96KZ3I1wROZZRG9CpAFjBpO
6M53uZBjGvlnWB7IX+lXafxx17U/WKc2/TVnQGGlj62UMbG89OLU0g2ci1Bt4jHbYygEmq9rSeuR
zhGFzujungpTkZp1RGOxkRHyXUkLwBitT9ivQuBzSMHxN96pO7qxXm3o9RXbhybltoxG+2JJHoQz
A7PvLvtsQgPrZo/mKDDznknnDGuerdnZVqtuCjmQyAr/q/OxeWD/xbUfpvwb6wRxdxcY1jPgAUm3
iHPxMj1jFKcLXPEin/sfwPJK0M1MFPjPsiT41pijstukz60GCU+HE6Vc2nIwwY6JVNu2kPEUsn4F
442Bv7saC9zdLkBGgQe4xlxKIW+OnDTxA3JrURHQq+TdGLECsSu8reqLTMvfvAT1yNGkElT5O6mD
Zn9WhsUypUErnryFFCe0h2k9cyMCSsETWo4EQMnQo9QGkNx6fE7m5RsP6pX4NND4TdCbUwCyXZap
DW9bw1tZ6XEO/7IvRUxch27XeGWH8mWyoaul9pXu9a+WK9skS5OvmeIYOquP8QyRT1jI7rX1RGQo
ad+2d57u2k2LQ9MTOMrixD8Jtyp/33dB3wppicoHbBLshXBkzF+mOaUG7wZwc8/YQ7JBofc/kQMv
DLp4utJQijOTOlGoS0yvqE0i1tW9shcSUXaUMynRT7HRLrvZ286b5eF1nK0dfzOKj+D/larW34DW
8lLoqsW4Gv9kmwMnPNfUG8yIoGQAI8rJLn5VIe01t4GOKS/3e7GcGfYNwZtX+9WSjjdGTCxZhppA
rQGUVPI8BGsjrYgUoJAy6ZaJ+L/dE7LlTTFK8Nc56NAeSboXaEdGhKGbxbJyBtcnPznazO76GQ8X
cL6JICQGgzzHvXf8xdza1AWSPfOYA0n5qycOakxrZLQL8gosW94OxnBkeZnpISMR5DQgpcWP8q5h
kUCaOvPpME4RS6WZaSXqXN4RGUj7mI8AmsSn1kdjDLt14Wt21nbYJ18O2CH3bP4BJhyU6eheRTDj
Si7Qf6mssfMCtKGZ5XvjN+/K/Rxx5yW16cf53/V3ot+6VHL0dTh4sx93/tv9ooDlDE9H1hVPnj3J
Pd1pizRW9Fwo/8nO9yTem1dkjipeYe8SasCTm3LwIyVvlUjFgyQRjEh0r44J/700TMwnH7DKMJDT
s7LC3xglEyyNnxvnUw6SLPyz6HBTU1bmA5TOFSPqoapg8rz7jgYP5wJrMrFqdtmovGvoYEefxMSD
eNrzA4opCBZkjEmAWiMx+h4J0/QntsFLgRNqXx8t+B6VDr/+m7dLnjPbvJInL2tka582QKxQzgbH
IHogE4B+p+dzTAo08ef7DFr5YkVFcXXpePvdrfGpG+AS6558ZkIPJ4Q0soXy+UaDUlB/OGZ1WTWA
5o5vdeg4YS36TlxK78fiPiQasAE9J8fYUewoqaLHFr8oBIMShY4rs66qCvTctAah2pxyVK8JTLJo
QTwNPcbnK9fyILkOejggfCsXHzOLSoBaoUH+oOU3fVUCox6x9bVA/m3MoBezC4kM5jN7sa/qnen/
V77kiruVaUOaNBQAk4rgxiK75w1xH3N7RjF3H7jEvbm7b7QYTWHudddIFCPD4FZ7Eid7Ui3EQLSX
Od5lSH8nkwgMGFqZEw5uRoWKJej8jUtbn9K89Fit7kyrSS6kf6FlMqqABv8ZdzkFHEYZQ6XC7IhZ
3ZeNN6HGLQLFZk+XC+FTLSTcVOT50ruGWJYvmraOTCiVCHdtv46pvYHVse7v4uoGDTGAGhb4NUQt
oJfpeJK8BJS83kLduYFdQpm8IFQzC3GqmbNh1/Iy3ANSyC6JL/2z+kpZjkLJspjClIb6fyi4zbWY
KKyVWnIBVHoHum8pAIO2Kfu7Kgef04Y1E2azD2MpUmbMEu8h1KXq0O4Yu2AhcLdQK/CAD+SFUeEU
nxZEDnDz/kvn6+TDohG+uWQ+WbeljkAS0qyDdpUNXjydRcbCZeaNjKs8UKJfq5yZVdbjx6MvcyBe
Xmtb8yiZj5/z1aSrcwUgotX1wN4V3/Ql1Y81W13ogJsqnpKA6PvCXOuspuALKGi8Jfhia8DIC5BA
lajcnlq9nqOa1hfbNQKlm/cG5fT3UpWpJoW6CVC//jdDisiKf5L5CsUl/Y3NNu7hu5mkIXDVI5nj
KmTseviAx2irhkN3JGf3kkBhLU+OxUoPrXpRaXY+Fmovl2vsEQfCM7AYv7DA9gn/uGMG0ZusRfhN
ACFflIFzSZBGIzM7i+W13zwgxGUPDYr5P9XIbn+aOBnk+tLtmpsYjl9h/3y6zhhiwY7eX9eYleCG
WkkhCLRneMrqRK1dXAEWmVSPBIvDKUA6yy/pixeKSyoMuqE/t2jUauEG8DrjJCPilBUoT4lINXsd
+4137eZDqCMVNDMDn9NGdylMP0KK8wYvkwMkRFwu+0+qGTwTBMIwZQb8uf8EL4pjfdxMYUPe/p3S
9+IKQmkjSCLKur7Myj9md86LlcHB0N19IaVguThwhSG3QcL03sjs5IRM/6I/2LM0Gjp6o+HL2Ym+
lf4KZVd6cheV1nOgAySVRJN6snrkm3Omq+kkwB4XndzZeeqo5h7mX1dw9WFkgjvnnxDXZhx32KWd
XMtPKtH/5A5LD9MW0denNXB/sAV6WdbJORUiD7HOYfCwbdfhZ2UKWqkGeY/UEkCXpbhvike2dkuw
Y1WaZqwubu3LOkb+eKe5GftWT6fitLuSgZSTAGwyD0giyzU3w69PJT1WOXErFPToAp3DB2oQyTCC
9Zt8emngj28epqUup2VVI0n6M1sX+9M65J1lYWSZsW54CiNtr02eCqamBTLlvOk77o/JfTyEBDC0
mVeq3+6+f+GEnsj2LxFvSvqM89JlI3/AgShmmDee4mnKGTmYR8sBM9AdWTvfIA4d9yBKGsOepx1S
kG/VezEkdBRI8d0CuOpLA4GkvUUxxgjoB/mrA+5W6ygyKgbM67SsBuB+Erz/wu89dayUqz7nliru
ai05Qfice9XrhbRD/fkHDAdj+FCDtvRqyDSNq3HCP4K43lj724YB/lCh6gG5xAUtYHCjsmhztdzh
pha4rvz7AI3NEZgJQbDchxCCHU3sDGCldwu9wGoGykKfDcimXxLDFqiM+jLd5G5PV0CWbRX+GIZ0
9wacH/cl22w2L9RiAonyQ+kMfPvk3MABpP2//nxuogUcx/qpSG4hoSbjmmQ+ANnM8PGkeeJKAmA2
AsR5pIiF4wUaParQm8iO1URSEGOU9J3BvFI7gdx/AfLPMXQ4LG5/RiRzc1KPtiFTgr6NEB/rgoBl
W2kzkOlSq1jJ/1L53VMDYW1I20VKj2q4ZoIm70N+4ii96fOD+yg7i5clqjtJrnYhodoMmyWotVvv
ttRtmKFUpO4lCbgDf7UY6icbDzQqUblA2Atz0lGQl1QcP+sJY7V461V5mhwYqs0MxgJTUev9gvHG
BXeSh5uJilF3mlLleS3xJn6z72cI3RN6Ygs39icSF6f6KcjW/n2XDWqpi0j7ScFB/Q0U48jZTlP9
GDw2pxUT/NvgcgljJYaJKRN23sAGYU6qHVNqoxpz94T7aGq2f9+KvLktV0x0eUUSzWCRlqyALElH
tjfidi251NR5i11btPYgvv9dCyts3fk2JwSr06ABXIsUpKCtIEdXxngsYCwQb/YNoeMNX+gdHGsa
FkOQiWKVa6M5FqlLK1yiBu0x5QxU8eCFzG3P5n2/yNG1jkuo9jdBesGgDwrjrZ4DPytxMnWnYAgY
eSlsk2Et3qFZnZug+6n6xLoDXpf424lbREkCzMhO9sWkDW/wwBmQNIpVR4KxsedWfjEB+OwVy7bE
lh4gldgS9+sY7Vo13ID2ALWbIfZseYRpniU0F6VMl4xJ79NHpKpHzOQ0p67/1MRmxRbDLvlKcav6
XocRYOmLf+4t27mJEu+dQUbJ1tjKrVwCYGWGEcXNTTMZF9lrvhg3yeaS30O6FP9K0CV8LcTASJSf
9hAJteYEgeUe1JmQ36yebCY9azHzOx4fNCHnvyomNI+t8Bl8Toa+Z16G88tBq1q5ZFaoRSG7k6bp
H9mSdqFMAmgIIlh8U2ZkgSG5YG/IPbkxD8Q4LkpneOayukz//eZdosBmtfbNAbVx90g/jUuQwlNQ
DM2043nLR/Z05twJR0rCEEKoj0p70GBgP8Nsvp56gImcWnRzuHxpBHBCuVP3jIcXaEvecD+/hkmD
BEI1g/C4JJDb+vuCHrpfk+Jz8OJzvJijZk+1NhL4xSe+qlYo3/ctKx+9bzRu9DjAZwN/tpfLERaD
Y6QjNLxOiVndjATvNSgQZ1xnCaJzNWP6QMwgNxjKkjj4fhNwOyPzGUuWTLwan0GVZHEKWNjP1wcP
nOc7Zs8Z73DM1amVUDxoPI9ksqkEOxrDTwtHb1dF65SRO0exke5DrliT7RxjQ/hvHSK53X+T9sYz
6ALc3ipY6G5MG4ySDImBB0sfBpTyVuG/wbPCra25ce1DVhpY5Cv85cKvVJaR1YfdzvRe2/087Fpf
J0/ywH5GsxpxttZ6XBNr5u+fEp+K2er9Mi5MLvhVHq2abEYVgb9dUqBe2LWs9prmjhlpuMPVvMX6
N8Hx4iyFd9N8lgpws3tsu31ko8H4BA3IrfpV4SevbJak2klQefBMo/ndFEClDVcEREtNzk9sMv1U
5/fVrURFy3aYIc8E5teq622j0tcSceMQCM81ZRE9ajv33h5ZzpMQRtdNXtGtgcxO0F3blKMixILk
g/71Tizk/rhjWSq+zu/GqM3vTSCFJ2yLEFwLh7j6Y8GsVnwmNclaUMZSnzM+fj+7eEpW6XRAl2aS
dvhh+bm5e8RIozqYQWcECmXbIYWCKQ8eUk83KgSXapTiBwG8nDR2B558WWsULyqeT7dhBXc9fcyR
JSFbZ2cKwC2bqIWX0zbDCPMKiAeTTWmL8E5e8nH01psiDjgZkgDQ87RlUuyDlMCpqyKrO+N/cC3H
xS173buujXZzZYD1Q96IiiOAizBOGba8Y6PjDDFCSpbgujNjSmQrRhbI903KZDkO8QDNTMswoWC9
NfM+DtR+JGKDcQTXYxtAUjmNk5HPnhhRc/xA6S/+o51X8iCoGUfFF7B1pJQ2bcuwsRH4lEG7Sk22
lCCbDrS/NUD9TehjyXCuWwOdZ9H0iLakXu8j7rqmwo9nYWwnH0QQ+D9GuheWLEHvD0kliLRTLLum
g6de2wfWkqDofnBaR6fLUaEgrtVo8aAUKpWdQtuCSIpUlHU27k36Y9Y42whpke20pgyNChf4YLA4
jotFnucDvtA2sDgqUJvs2fa6vdfxPDW7aI2YVN7Ns7Y9caYoWomRNGjfXIM6wkR3NQlcBqP/Lzox
Vu/J7imkMwpvveKWQIP5EsH2pQAQGX4yKriuVPr9vRxdU+jSYb5ZFvjZTvNALuu7TAAFlCvQY5tj
TI5hOVgKXf8Fx502HupYOvM8vU8otH06As0P24MHuc4dG0c7y7YzL/gh9ziXzCZRGGip32CCkpx5
o5tyO5jW5DIDVCxvFR4MvpBUbd3Qpm4FGZTdILBPd2Gy5CcehwCwaMMFMLIelaRnU7Sy+SPN7noT
w0bmn5JSgEULiw0iGaTWZ4MME7cHAZG2WYCMMmhdnmjHY9JXSZj3L+u3yu7AR5aSe9HF9XCzjx2m
E/pl1xCWhckhfdfz0n6QjkAGmSwnSgT9VkVfTnnBin2vdSsrQY0bK1NRTj78GZtPYLHtxjvMe9uu
ELu8TFmndt9zwyA2MBLJdQBdTNlGnkeetNhdVLpKxVMQ8/HlmcUxcgRmiJw7amsNECxE7OGB4AkQ
rBCZvm92Bx+bTAbx1I/bFY4BZ6TOucv3okWDyq8TIcK5FibgtTzyukmdK7xNSybEYEPsXTKdnjta
d9QrEoDPzNAEXoymJU6owBnmY0sUNmIdouDKlqH6cHsP8+9tmMcIMPV8A3hC8j39D1KHztylhFm2
s6sBtgHyhVK3Gw00IJovZocMPFidBz/Ww7un8ekm1PvualKFn7Mv3QWpGCBIJUSqdi218kHMXJZy
Y9i9RclKRTslXKTQ41BDkQwCqr0ClAlDS0yp0EeDhEMRIUWL3kHBb3gdRkmM6JFC8FhSGP6PqRNF
XL8c8DICRK3tIZ5ApPkbil2EATOZxJ6rF+bOStjsyq6hhjmHkce1saDtPtG2xW5VcUrdh/a0YWnw
PcF1QQ9wUmBco3+stgnd/kKsKuo8z5+iRsK/zL7+nSdvaoQ2NJzmTs4JtqNZsmudKPUYimXEQ2i8
l2H6ZT3LBnIp/rFRykluw90ldXJsITuMh/L+edI6gZADxz3cBJX7RnJnzES3IWFnCXrYbA+U83tm
RRPWqRRW8HNsdYstqlAaOSqV1ANciIoEwKyDcQ7tD8myGLNYIPXJssIoxoO7H766HHuoZpfgTG42
c/hI5vYHa5fY5IdTdPL9V+N0IK/6fH7p7+LZXUmuvYSuHRUvRlUlhrMgeeGZR2HcIOSQnUwQirjy
cZ2mnsV5szJZtgD9jqK11XxJv3N0te2RLuZNB3kTD2jHdRQK07Wd25R6Znu3mszcQjhGPQUrg5Yh
1yosZsISPjYxnU67VudJyNDCxvz2vgNNIO6oTmj/7q5pelDFuqKQRy69R7cD422BPeJEUvcgrnGw
SvuHSnnONFxT/i1xNW35giOM1+anjjgGoiudgf31qxzD49uM2Vfs0EJ6OgevuYEGq1nFNIclNfuF
jRqa4WFe+RX1HLisIHPoXXtnhfbv9ZptSszsRafMR8diOy1aItStPR3I8qtDElCj6qiAqeu1wH8J
QvlRrp27jqhX7DKOaLheLX6QjjeCRpCVnljyYWiA7zcsMqRKlNHWc0x12DC7Ld4HbOM36ruNkFmi
4ITUaSWAayLebVCgS4yDpJhzn13j9PmsVZo8UyTpq2ZA7j3v2+Ui968cXU1H6ikDrgtsPJcfi9Ci
VSr5Qw2TNQBOzWqL2/lToM8HpRSruvkEAZ5BL+rsnIKNmwICJh3hb+hFHPDalvjNDVI8DZFr7WBj
R4zISQk1yE6Jb8h/W02mo42O9CBt08cq4aOlEt/dxqtv2YSW8WTbqm11VSWktZecH0Kvs3c+1DBG
DI3VceBZGlQrJKyTIXqXWfAmwo4UYHcSo6kb+fYcFiCgnvVhODNjvlzyv/L3QiYC8zOPWB6dpZc1
9y/Wq7N3UjUaNaeSC8wKVsQgwoWOQu2OfeXXg/VbvfKdgUXKwkjsjWIciWWanXuqBfo8uahWPBWv
vMhaBTu+erxJ6rtrQiTLndXGkJqz7l8ZJMnafFcxMwyKgxJpCVYBCp1zeo9Arfy6cUcxGFOVmH1J
Pj25IzTy58AtejOcnTs3ULpcmfQnfB0CdYEix8oYl0nw89p543JcFr2Fo/89CQ1kYMo0wZgH/j/H
4hM3t82dSKCG8nqkQ3ps81mwPZd5R+vSxUzXm7T84/GpIB+uN+EhSezclSm8Jd/RAyy8s3uV58kc
PTeRniOYehwhHq+2NjVBihi83nCjHo25WNWs9MVYwwouti35KR6VCFbohBBP3HzjQpd0KlX/Hc7G
G5aTDIcQUG6P1oRbU9OOKh/s6pT2jI5HJRr6itpzma7sklYh+nuZgTaRMc4IlHdPjm5JH+5ONC6/
uN3TqPDlPMv7YmOPFwn2DRJFSlHmqS9ITIaqkZWi0ADFybDtqxOe8gd3MiYzFL9YaYnq0UxqqjD4
anFu9fSQdu66v5FVScomq6gTkifWYMfEOwdFxS2EvCbKlRior/YZCE9Dahv4zzBePkYajXnJ/su8
UhUDaK5p5xNX5MxpgnYvVlrb8g3nnXNdsumgTuyJh16Mu9bHafSdPqZede5slPJ5m0esyeBy1s0c
cejzXX2D+z3ZTXsXl38ht1Iuou9XMZtjg/t5QblMRKoS+qY4T4BMZ45lV1rrAAAg1lQVNg2g5KtC
ojqBOLJJ9Y511HM/B4X/pieTNq1KZIhcbP24H6XjhVKuDtRIqFrZ5pDsc06b7aVmyW7LxS7LeqPO
erzdMlIqfUHpAhIlxvcYUaSuWgPz18XkHEvMiYd6ZOYJH1auv8WCJYbRDLvShmiI7IGIWphfW0tr
W06H6Opiw3nyTSRl17A1OkA8Mv6peqBme9qMk0bUVfcxnCbywLSmH0XFX73yxVBEP+jUK8o/sl+E
8MKnENzwL/1i6lPz3BHdg/Z6lcq80OJyDKvumVwm//W/9Xlngkxf2giRNsGQvG8GNe1MLXb4xzAb
J4b6NYaxRrhNnJ9Tg8qQGNs02LODfJxhrawsGQqnWrHc9Sfh4EgZpzljefXbt08omtN9w2i6qkmX
/zqE4bym7Cb2BjBFSpaWCyvn5f06O+GuMcm/jEm/avgmRPANuuioJNY6wCMTiRS5thF5vaix7nb3
D5GvW+gdlzA0MM5/F38D1LNmNG/fPXM3b2N4m4VLrzlicoo6y08DHBm8b9cfreD4FKc8wFhxbO5g
SIBSnT6djIo94wKaKWGXMYK6hsxFHNtk8wlXETq37hdGrUuH6k1mgbKHUoTP87izLRl6ACe4/bsr
FjZP9uNl4YQ+1zcyp6TSJFNqZtKRKcP7WW2/pVY8z/WddywCOz9JS3Nc5u4iqjoHt27xGtYU/L/Q
4XKXV+qZSKEgyqKRYeMybpv90AMVgxnFeOBNC1iI+bOYDNpr412i21fBcTZDk82TDNbsuwZeC0ZV
y/MM5TdWkx7a1xnvDTJ62rSfgMX11jEQv84tEZlOarnIRY5rRoRR6cbF8rJfKvruOEp3Pr7upNC2
RCy6vDmqdph1+G0x5yZwHc08Xy+xXeNwV+fKoxNNDK5spTTLj/2u/ovkWO1qzZyhSaHw4/TLR+25
gRaCwZ2xXCN7sKgtkWw7XuqAFOy7rACBOY2n98HJtR6DHbkh2pJ6aQZzUpY4YiuAcu+ViF5E0Gxi
Il1VV+FejRSHsBJKLBsDg14u9H7NmKg5pduDGfnq3lMcK7kI5cTk8Sui4w1ee8DF360y61bPdyig
fzFehpMY36uTeUpLLmdh6CUlkkSsqI63Cz/foGlKd3vjLJujcyQCBYNa1DC+s0R9bLVaG/sTrUaz
wngW8CSrSHpo4w0k7vCZKsHi8D4pP+0z8gCu7neX0/eZaY4fKHrr1PSsbWnJfki+APlS7ZkWJczf
WRVv7VN+eAHSpPKHVvTg2yf0T7+57neL7lEFXraEjDN0vwUwxJSzeAK88WVgwvmx4qVhfCYimh7/
8+O2XhnPFactegLY7KJYtgWc/LAB8VoWB1R3P0tSxZwccOw6MLi3omDIVkPNkgjzWRKmZ5HqJtxs
VdTm0RpybzqzTUaH9M24v1k3ocTEi3pPru9POKyxJSlViK8DvWa10q2fOpdw3hSOp6B2iwIWAtdg
UJNsTkOIVDvOj46QorWtdon+PBhKY/xeFuT87XsdT9/LFp2s7ENH008BM/SqDs2rExt56bEpZOV5
HY45ts9wihLMQTAbAmYdQjY/tV9mFtoJ+z/Pfqpx29jc+5JtndLPks8TvbiG6xKsn9FKpP09SzzI
aqLsBl9z0bckFcvrNsJRTMg4IW9FkywNYj2MShtQZ4QzqnHTTwqOzFj431SitVRyxxCj9k3UvkhE
O9V8Q51VQ/tYA07LazeZ3fEoObwpzaYjvjvQDWELTlKzkDKJr0hQ78t/8zRmgqegqDxzWNyibE71
3W6dbfKlfaTVf4YNhndtkUSLmFR/IuYB5Pr/p8JtVdutU8bSw8lblB7jxrwdwqMr1miEj6+01kJV
hQVyqQrM5z1JChPvtv1QtiUQPVpc18CHo0XX00Uyv/yalT5ICyNgKIrHoOgPdvUENONiwz0tLL/a
DyTRXIHEoBCeTR9KMBS9ld5XZvxvJnDI7OmR71cxrNK8iNaP2jqO+VMaYJexgB3iH2Ep2zJcKoEG
myi+VsYnBVLHcE8XOe6W7QLlqslQ84zVW31vJiCiy3cczAJ0pMBDvxJ2N5lrFUDdiJYiC0b2JuhI
eZUgZ57NeW2MX5Riyy+iKw7y69jipMdtw3gz0kEuafiTgzqMc29DiYU47daJv4Shj+pSVFrsjZlU
9EESqajGjkZ+OxaRItwKH/xmrMI1IKpTPtZvw299SX27GLF+NEPwqdbBb12A4i7ag8IYhuvz6nl+
EgM+ZzF/JU6oaC8vCULbU5WxOtWDhH9aYkrVrGPtq+lfChEsukTpirQaYwTXCs8HrZSbrAWqMDec
jTco4VkK8KxosLAiFk7D1j9Lc4LPfL4ClPAxvQi50BXXfJGBogTdEHlUU+u4+FP5BAxiK2vI5mnq
N6lLwzZSNBng5pMtbubGX+JSp7IWkc4bYrevKEAlWKFRKN2s2Si46aMA+aJKqdJOEFho9253FJM7
Qro0AE8o2iZYRGxyPaU87XqeiMMAqM+lj/Y1Xnn80TXu4lGX+sc8Wi/4wqh4Ft2DQwNCmmNYbTwb
Qwfy4RarNcoc9FpLvP659NCXAJiJwfexS2rw/kLYmH2I9v1FST+G5yOo/i5G3X9k81vjtsH74AsG
Z5DUOPAV2dcwHmmQeD+7wJVeKkBcLcKcwfWG2rgaxjsyTmILVcacPhWMKzLL/WjWwLhjFQbcudCT
z8Pm2MwYRHtMdpkUVECQ1ZyjxXJvPMECVb5iNwLMPfWfjYOReySHfh8KkhiEUbWgUwN/tkxftOgj
yDvGnDS9wIonTBuzto2WLJ6ABpFcbPqStGmU0mJQswS6VniGEKb1cnpXUnjMXAj6Lo1ZtUc6fIlT
gLaolK0d17WqE7zI36IbWzMdbIgdMfa1XIOzByyma2uDsrzml6qIOJHeBqZHkBOTLCbdLOVwboqL
xmC74qyQK3qVt5i5k25njBYN0DMQt0wlvAXiqax/yQFs6SfOWL7meLgMpdhrkfH9U+Y7xBOZEaLi
8TbeV83LIEC4/dbp0EwBROJzrrALZTvwa0NkzC4+hKzuZzIPbvzXr3jru/NzvsGseamPzSUDwf+G
Lz7IHCFux73KFjWHL/2gXVKdfFgteNEavpxyUccgBonK0zTt5oVbRde8kubSaydc6bzUVnyjZamK
qiFop4+KThqxxMR7zmPUk8SMiGmEnLAjruw/zJFTJN481c1FXCPRsio7wLdg6soEK2m1m2WoM8Jl
92kUj+dLz2ECiJ8abj5qhmMbWaCCM7JDx4FyOkj9BTN2o4gxHllxd2LNN0+ut5as34RijKydSdBz
lDteQrhyILUd9nBDZStcVbUvOyg5k8nzSysitKW80l9an+VJLRk0NCm6O+sHZ0Sarsnte7BYAMvJ
qCoia7iUVVd/O3H0ZN7GPbDCQs/c5Ga5P2CgOX1J9QsTCXgjiWnAG1ZC436+ZOjd5f98woB4Dz0V
R28DdgGIm1r/DQyrEmkPS2RYGfkaXhi3u/IhZrQAlDDrSDHmyOAx3CHUNFswGFa3WGjMamaveOoM
cwnZyCSAhKWz4uw12VfPSjJpfTRLTarAz7z3RjsB3OI7uu91Sstw63HE9cL6chZWFRxmRMlgn9HF
CjIdqiTwoBWpq1U4NC2P88SGHLs7hGG3hmmjGgIFOvo2+bEAzMVCKnjZU9VXF0tQapSkptShSzVa
vOmMzbsPOMyZ/zmgfsV9SrJp6adoLvHCUYbbHRiyBWUxJEOaftom//Gzwlc1srH+8MT+bsnGfzNH
OSY+FZyp9Y0onTwpfHqI5fHqNjI/D9mzkh6B41cGEoebwgbnUiGJzD1CFJT4ipXFEYH1TRzSK++z
SfBV9ipfBYcepRQ1kJrnjAmjQFUnKQkbXnd3xZcl/X3DEThRfw1e7cK25srskxBC9rxbeL8YiQGT
3tQsK/gU9P14tchZRR00aX7hn4MJh1N1XkjSvBUNiDjp2xtsmOwEO2T9p6VC1l4TQIq3pBRm8Zqh
FDDFuv0XCSbcSkVEcPK8DZ0yLj/orBRZqR9I7xjX1dufivVBwWCvtDeOp8YrEgKofjDW7KRwZDzJ
izT7O8eZfrQubWSFc6UDpoMkYtawnR/9N9jNyfiFPS7GiILZnFwtA+Ze3Ic5p3TD3FrCG3cosK6v
K6lnWvy4GvulkjeU/+7unKyaxFFrNM/PRuexUxIXzzhjMW2E1nVZ00Y12J0+CyLkfwpARNqQAmOT
upAvaE+xviVDQASYG54u5X3yNfbPiHDxTjwBMDutHbVJz4xNdyFaxBcQFn/0TScSFXHCXbVKRcrV
XTuk4NAmLumlXbMt5sq1UvqyjA98OCqejZIvEJef4gvwyWPJT81jYkUTjxlWZxAGKXGoJMWdo6ql
x4U0nT7SyJOpybyaQPmrZwymcarep/YT3j8wqepEjY6/cUVlktxiGQX6DwgbE9znwpy90W7g4Flh
AQtVt8QRuMOqfsg3/6AVQUxSAKte/Ax+6Q+5dUcR/j/DD+z9xdcShsqGHlK5nLpUlp0QYm7TGlT6
vJnyo9HxT8Zi1j9sEjSxTxlP/NXtVzbpFkD5Wnb7wj2cDsclbCnT5X8ZQAIRNvenUiQxQPwHtFje
NoCVbtrn1QiUXnAOVkCdGDy5EvrJ4ROuoX/6Cu96aqG1qZk61SHfQRWAnpi3/7yPjpa7YKi9+6Mk
GCf2o0TRn8gON5tcjhtmNN05pd99MgQvg/AA16CdmtniRQljHb8fRlCXvmmLcLQ/inAsThp/urBK
yLBe7wySernkuRaHV9mnuQNXw6oVXldmoSprGM9qLVzWm1goGZXLNRxZbpc9hMSVjEPy+lkEJeii
WvdYveobgVLmym5auHbYh8NSgLodyduJfYkBT1vvm3nSFKJidTvimstYXzHCakX+1rjwtiJ0C8Og
2Bz0LIRGanGGQFJ0U/dDGtpq9V+kJMKgLOkJOvhv5vGG52OF6ZO6JEPAju1IGEwPhIU0ie+mUrDr
MBwwYxoNPNet9VAXu6+0T3w6PzTn1fr8+wEVr/AazTUWfceSriRu4Vrmsr3aZOQjoIUM5fojhPR7
8CIm5OOHLZ0Eg49fn77+NQa6j9QiKuvEzdzOzl1Et+PbQ6VAK6Jcr7FyhTJJMdJdzhVAIvnOTX6G
4YRB6Fi4USodF47RfaPYkO7r2DIuLtCfyQKRK0v/3iJQ/36Dl+cMMSsfHkq+zvLnU0Er4bB10Tjw
daWqbRo3o5Vwf+6zQrVaJzoBn5dIhtbhQAZ/lfQeOn1GIz5thHp8FJbR70Ujh2QzrA2v5JIHSlWQ
cjVSsLQBYTDClMUAdz9vshtePeqA6+/yVoIUlyc6T2iE+8L9Uzr57WHvmx/aFSdJbKfO3Xd/OV/F
5sTY3myDPkLmxKAS+cY2tfps8o0YOxzH2DbpsGgshmS+ePTCdtr9c31kbSWcAmNc8eqPfS7BB1dh
GakgOmoggXR95+ho92ZPcsw/JXCXwM1AdKG02KOcz53ZnRx2357yjAYi0iPCHVfaaPV65ZMKxOab
rQNMzJOMXSwk5u/fRDLfSTXGMkx7+OWr89PV8YRZ8CU+6ISV1DEmeltpaP6dfv9WETD9OWQ9bSvn
M1nXCjkOOgIIMqHx682uE0OcbVS8DoItdUjB6odt5Ij6cc2qhMdMP/fJvulibn6NBaZKLzJn+7Yr
PbGhMd7jPm+oPCgzeSPKB6a0CrRRdQUZJKXzfFRP/DObR9M3gNrLlpTtyfu2+DvXGfF7FF+D1L03
gg701L5E2DCo6sSkLSLSaGsKjUR6mvv1TKD9bxsYKd3BSb/BFoyX+gRCwhSyGQ2JN95jhTw8/1uJ
f9GWzWtUvF1oWFqk/v5DzYFgOtMxbcTulVlLldLETmMH6r7QmRd7BGy0qdZv6XgRi4BfZgrRspli
MzCYl4Cc4WwAcvk0OQ65C1N7jj5DVsRZz8+StKTUS/Ad1P/mG/5Ag6xpAB/7Aw4q8MMwTxTapNfI
gdQiHepbMQR9riigTkh68wg9H4lkpxd28WxWBNKV4QyH7NJOg4bWzgDeULpJVZ1ZapM1TatQd0Fj
8if09QYXVCq0GL1LO4w0ZNJ+EpRVTvmQj0AB/H5j/Afo73B9o10mzWt5YeQQNA0hnn/1qUVN7BS+
PcGYEEvPA5Ble/NqfnaeYismo1ddWNLvIOmaaXh3AAU5B3sMNXfVj3PHCJGmdIF4Pwk/ftcNfVZb
30ryE0WOaNDpkHhExdKhLsus4J42WvGtYQ7X9Z4RXAgbOTWWLnq0K+BCJtW3KDmhfw9GESNyUfCJ
hdMQtXl0PvMizIyOKWfu2MRaqdMJmhI9xxKKZzNeg0oSlNSUREw20GnHQjqS35e6sOXnaYjN3+Lj
6c4wYq/uboZ0b89IxrC8I7wupQoxn1Lwf/HBgEBQDyLd5NIUwcoIiraUfsq0uJFSqgS4oXCrJgpT
r76OdASdufZI+2MFf0s+WIYKvj6sKVAwK+/RvR2tUsPVVDrYJEPArcb3othEmJra2FcIuelDy/R0
TrjYNFxksVD3pETZRDa62jNPUw7qhs8sP+i+zRO3vfaIPx12A71pR7oMRH7zsgw+i6NJSIszYWn2
uRcYnSPVGWeHSrEJcpMDDN42wsef74keT1leUJncx/61v25AaacQaTbIiRn4rxCjChq8bYkIXKPJ
9uQMyCJuWRRj1o/9O9yhH9Ax0a7CUAhL9DPO1JZ3k5M8XqUlN3GQCOPeck7JKgWKkVPR2SE5U2dZ
10TT1DvsXuesuW/fZjfD9qd3d4YGrdAu1SEVJSFRe6Dh2WAUgAcHeCo/HD5Tk3LWLYJK96oF+pia
3Phf42I16cgoYjUWdjeHoRe/MitBgXedKgPcEmQcrr92JhrTf4dyzGVhX1uPtdHdTgT6BHYNqGkh
uRjowFAuGXlXl23Whx28PJRfIPVQbUNnwU1XBpVWDAO874jRcRNkuTCzW/MUcaI1IvG0QR5mhfgX
YQRVXh44SDtOK+4PFssRDgstC7OsocVMWcLUDUFF+aWqyPGmcyijw7w9nPcivt+lS5CPwS8q/7Jm
gcuoQbhRGmuzYnsA4+VBl6gNAmXzBdskAO0THFt0UTARJZlRZIb9yoaMYY8FQdEYzsZ6uJp1px93
Epx/5Q7SkvxPVsmkyDRfYAGm6/tYsDxQPLq6oXLvLZkGmAD99ZL3IKgs1hYglO2EJHcawynEyUMD
2PVi2/nUxtyapFeH+s19G8K/TQunXKDT31cctp8WqseeArsqAhWt6/o9clJg09dc9vCWypfTRPbT
o5B4UP6n4JLxSQYaoxa5w0YctJQnxPllkV2ECrNF5IkaQnGt4rnX9q0hgigYjyksty3mn1TLtu0H
WB/KyaQH2sRU2yhIzDKyBJa2LmeiH+5SDbgFkdbJx4A8sItfc4bdQLN/ItI33/IiJq1FKnIwkdFA
wOFGkxpj8C5vFFH9/FgOpYR+1kGdOMj51D/ftUkb3Gl7gnfb/DEoiJmJLJ5OG2uFFFcXdL85hMF8
ibCU/VAgxJcRg3pplWUbiIBErOcdcuf/5r+dMw4loYccoHVsaGmmwQRfqzFg0+CqPeAepDeEkuKf
Z+dQhcB/pKoWT2LXWopkkNiEnQuSlB1n2HGbJYl6erDTCylEGMG6/ZBrboN6aTc5jD4DjX9VAXxV
GwsgX+lliuULEtpwd7ssFZeanenz5vzKEHkPPQr0AY+6J2zK6vPl5lqvdD7B6a83ajaI8xyLKjy7
+eoX8WUrk399q3kEWI8+URhqrWUqU8kSG52iS3veHCqpqo0cDakSgC6B3KK5apEiyVBSY2jk6JY3
ieEqjYrNWfQJNzOw7kwEs2bdhtNugSOGM64Ir6kb11KrGOtqjrSYJLX/gj1mJDHQ3u04qUOmCzsp
rU48NC7sO4kghcDa5zFWfX9TBfuXqKBEWbLoEaLrPOpY7AJbyuH8Rd0ylX2cIBtRPKBI2ORX3JAl
7ARrWMfcQgTjOG9xDc/XWulUC0FSOTQ533KsslfWwHyvDBznRiVCp/zw0VZu21i7vJVq3bDgjHdG
lDwhTmmVD2J7wDBwhBOSe0Da4hsZEJ+JKshx4RC5ztEqgziBMACDeYVtIXsBB3Zt9UwrCTauCsH7
jfJcJV1+Y/PlPCx7xCKBEE/BOQKqwygIWeyfWiCpQRWYqRviNIdFaX5QMyoXDz/eeLic0N5ZhLKq
+8RqAfQNoB/+VdOcmG7MZ2c9YHR3I1CXjiXK9Xdtbeb9OtBFyrMW3dUirMORvhDhtcqs7wdxqzDJ
AmeKghHTyFy7fqzlqt+AnT/dsx1AQKZwjakfMiWGDVYdnS4N43DWYrdu3BSHCRYD5sY7Ogc+KsCV
vU283MxpVjxF8tJ5EAYcjnCqCEROkJQqURrzsXcvgEpkd15krJVfwPuv3cA8+FL5uVqWr/SlBqD+
mD9QzEGuqx04yj9lM7Wx2gYMNN0ohWCrUTinEYTVu0YbxqITSmkT+5sMaxDUOAyyWEs/aSSe2stk
tDF0wIssAd7I6bEhHiXoGc2Q9MNcylG7YCZYaDnJVxslfXksgSwGoAASxNXOkheh2sBGtqwCiEbc
mDsznFuUaVa6qnobEcZe8u0oO/BIC0GFTFM+Jg+BpOsCLwhHBzPpTbS6nIACox3cvX4tF5siYOKH
SvqyvS6gf55jvWGCfSHKz8QgU1E/PCb/wueqEuAGhiL38d77tF21JExpc/QfptO+o9o1Z+Qu2Htq
Vif4xVbAhwDiD0Y/FOda1stSgx3Rw4ovvIcxE5KtBYQ5bAoiMpTTxQfLDBDRFlAcs/iglHwjv60U
RWGzzO14NHwlb5LuGbdlw+UMjLPGcejr6L1RwCbE7vw328WNbKUlhk31iMCwWGn87LDz9PHOyXKh
jq/txKXH35nUBQk4kNiDbm0X+Lv4RNy3D3ITBVMw9yfGHaDc0n5Z4ggsuGI2r3d8hpC/4wBr2QvA
UJ05a+o2mXOR29gwTxH2OkS4CW2YQGUSqzTMOFZObHaA+VK5xFlqoKwRflMU5WWB8bj66w2GUiAO
KRWkjGFEvDlZZCO3bg+e+VJhtWiEfxs/ZUfIyNkc4HjCEWHdd1AbZaszT0sx00MNfnn/EpPSJQrq
crc6Khu82Uu6nWi28uxPWe3wyBoO4vdLOx05brw6NejryjSYMYFfUsfAZm04fdZIOfPpO9biw/kC
FuzbCwRdp0X6us2cCz7vbp/9FFjKNvhsSx6JWInY0sTOKQO4o42Z0hIxXj3UrBGLpe0KjojKCI0u
EwRoGSOLG92ckHc7p7prPVeRXHB012c2gy1paSHwlN/I0QVKcJayK1iPJGite+j7pxu8Fl9t1Q7c
Gn6wgKi5P3B74k/wfwGKWrUBTUcixiuytQHehiYSmnRbSTW0gWxmlgl6QUCJeRxAIeuJ1LSTLxEk
fH0tGm+eSL2kmxgYY4/9b17Ri6kJztQwaOY0RjsuKnFae4KwL5r/fnJPLjF/zJZIFDBGS8kXb6jm
nwCaV+as7ctXDhAoW2kOIjuhXtuFirDqIvum1/y9iw7W232iknL87TJytGWUubPGoUJmLATUuTO0
lwLm8TB6oIawZHcl+fTtBhUpnJZtYHzaz4TStfERe40n918azqsieiI7ONQ5eADq3WLIZnYJHhax
Si0V3ZmqPkC6IoLNyxzskp4bxFOvsyEL04ur0sch+odog95Kxvq3n9x6qdMk+Myi454TDyhjt1Ra
bjk2sUl21MgjPm0jAFBj70LtHkH++oeh9/8jgNM2lsN3tnrFPynApU95FeuGh+1Pwh62l2amKqLG
kAtDh2Gr4SX5BElwRg2wniUsn0kGWCmEHkY8Yyc3UWOFkA1gpdF4Ves5JmVqe+89aLJOcR3EN7C2
a2cFvbLh/iEc844Zb7LYjFCs1172yIoJ3ctwNcetjVth+TeabQyZqP4W9G7nW1pv/CiiiQ4lee/w
wz1QCnxMa+nUcGShbqu1GoxjldZMu62d5puOBRWZpTe/Z5VvErC2hoR5n62GkFnIM4R29+w5PebT
iiIylyJOGxFEUoJiyIyn2CsVUET3edyG3v0+38FHg3dgbOPkNcDhjfNaLBXfEdzdoxNAD5LEem9J
p/+25WyrDjKRERDRxhHa0QjBrX5J+Sa+cgBqwpaLm+GD0cXPGHFIPmWt8kfYRwtdF5L/5NCcUOpO
xSjElGUSH1/Gy7hbn5TsxTHdm9w2INbQlxetWl+LkpYUeE25tr9xX9OSwntktqRqYmmoQXBpdFBt
4sz89P+T3JMkGYhyC4cGF1xh+s29RTWj5WefxPj2TEaS04AK5H0CUgb8KBRdGaLTKxYnELuYw9+J
5/UiVp8SegOB2OpbK2qbzIs+brzPKQj7ZD532eRsaNTTmZw8HUMNxylOu2kN9QFZ7X6sr3o0wbaf
IS7bBIcVGC7YY2awa3SmdF5nYhsPERKr/MIh9VhGWlHKwnI/aU1OHpe0qJu+w3euO2hKFP0EvZ2q
grMxsTWVTacJ6IjbP+sZVjSPk4NVF6okP98Y66QA8jwl4QiOWkclxlojgA6PFzK1R+DQzhJZrek3
+5YTiTAa9D4y21d1/mnfjI6j+I/j8CTXFl976rP3ZScMZJ1g6izyyU3Z+9X7Z2bufD8IRG9uysZp
+p6SpvbVTbGTNRj1j0RweqNgMPNP9h6uwEzNd3GHQGiQRyS0WoJe5cH4ZohPpRyGLmPxhgtbf78L
3hFvrmIdnWlGsMfWemL/kYk5H8okE5dbYrh1NH8vtWuMxWtgie7hurdd9g+fygKnVv6rSm36qJFc
Tik5bF6JGBizztLQLlrba/S30BYHUtOTq3ixVPxkInVrH7Vk5RuZTN9JgZH7svgi3/AtYXmRoaal
MYKg36KcSD/IITVaIBt1uFveLBaQ+zNZxgs8jJNv4IcLmggm93XTO9Z+qb2kDsaSU/Lltw2aG/0s
XPXSA/J1TnOH//rck1y9erb3ZVFEfrxWAM1kjDwTIdU7adsfXtPgayvknjrF0pkQjz2MRpmOE6ja
uCaFetAZglpMd+UAeIKc5+DOLJYRI9YX9kxv2hFkPZ6EIRpBlP6Kw46HLwO3FGd8taiYBDNuQGtj
7Qym0dlJkzzMu6mEY6gjFrSuPIbl8tJUXS7HEZdbZJ9aLfFeBQAV0oBgpkqAmkRWcouDv8NS1AxT
mD1O9fPY4j16OWhr9723UxYjTcNEfQUztqjzTTIUS6UfR0rRcoIcIRhmKnv8If409J5dKgmgAxF0
PL+95xnZItOYN4wr32ofVNcnhsciQu/Wf/zbF2J3Pvr4ndq+PTLLl5K+OdrvCeIExYa2hRvAXAIz
XLFgOUOpUtrIKb6JgSmLoL3QOrOrpzwRt8s65ky90pD5CZ3oICKqlZniyFgKS9odbEevPXMfV3f2
zAzUsBURUzSDodSj8d2OH7dzslGuqMsNEzB/am7MOXHBdYDtGCp+kIrDn+a+xp2YEnX1uhEU7iAG
aeuSBN5xnLGlDDMuc15bs9Q0VSNXcI9g88mpWLjTrEqM6iMRLYxhFwMxlYHGFs/u8nKSp7ZB2d8Y
hyNswhAn6a/FrEWmUpHc3vG94QQyr0uPDMq4cPQg/CA3U7sb1pNgiJOvLQvtSDCKo/WO3mIgzdNC
GIwhIXTsx3PwaNslFCTXOBLhFRBBo6pBf86pLfiTZjVDJV87xkJVwflxUGvuBXE72qLC9dK6Mp3M
XtBZKV+7u0WDXRSQvKNIlQdPDsQBUykGaObK3uUJElhdlrlx8jk/aRBC4nlusAYNm4bHTYxtEm29
3RA3cvaMdgRzLeqvj1hO9/ycH2357A2ZYA1MITHCoGFIlEyNnKg44yPk6/ulRzy+kpXb7vNIKhaF
mkjKA5appH5hbnBZPQTpwkaCs0uwsfhsL6ZFXtjGZTX5Cnf9EII9hfjxasyS8SzH4c4Wi6kKZaWv
tpO2Qq5AJxp4bCuXsSHVbJihvXjb2a0yVF4A/9370svypIuIg5u0HXX4qzLAR0f4RIeqKpOCzHwY
FHKOhDaer/TPt+bJl25+wYXKNE2izBo0DFiRMi5A0sPPSkmJ2JjJPszYq4kGp1xZp65/MpCgno0S
nl1BawHu5iFIsW0YNYhQ2A+6MEpXcr/rEQ8JLhIl1hsQQkDg2SFWLV3J6koF5RH9baYVYZN+R/2U
lHgj9jLD1mibiy2y7wWiqKodZ1gT+976fuT+Qg5XXsjVwp3pPqAIUryJFTQiXe92mmorHz3YfFRk
TJW3QdSC9boUuZ/tmAyU725mc41SRiPiLhN1vRBKIeoBl9sp6eJJxv2R0i9Jc9NzwJkBXhg+zuKE
mKh+oSS++3U4OXqClZuYXf5jdfGqWEIgz+q6aNKe2Cd39P6pRyo0TrINZdt+5HrJLS0zg4pYYyx7
ucOnyNDRPdp2mSg4n7mDwqbvJM2+ObgurtuGfSBuZ+JlZkXHOMhs0+2wNEmzFoy6enGsFuaaHB0G
NoJNGNd8DMnn2mRSdPytL5UalCQdhueTksBxiNca1lofW2gzn9i1/HZTOEtNP2BmRWP+XoxTEK11
ueKUUAjdE13OrtD5eGZD0Q9BaKyU0ebFYkNdGf9G9VAcCX8TwkQlAjSYPB6qTxo9c3cpNpmNcHBy
Mop81J08euyUnywPs4bFzZhI2XKJVweZ6mwoT0/H7rYOnLlNmNFYW4Csoogu5uev25JBSRYN4PF4
XV3zX5i3qTAg2FxiXZu0L9ce4lA4zNbuOOVrtAdLVgEGBWi9f4aVWSJOS2Vqut2cBOJktrHCZfj1
oU1xPqs3wD7DivWlqdRqNISEac0FRhGxuFURqhz8rnbRpgFUb39bsJbX05h6dBL4BGMcPkJ8kVat
zIdSyB8llw2BdKHcWUsQ8eY2JYNgkk8vyEqTSqaIjkdNKoxlSugVTd33InZROeA+aC8OrsBuDIUp
ZVzIgGVNU8uTs3pCzvwpXIL8+/w7ks+9+MGAI2SvghZLulj/fSl/uuaP8EBUdW8x5RKo6F/HYHL1
5xyAMrpQjQnLVhPaLkzsqw72708s299aXR1sI/PTKHBEK8AVMxB40BHa+UXH4+5l6FUevSeWeodd
YphwWMq2hWxbXd9NDVa/7JtsW8x0JUicwPcYI7zT3DY5aF3cRPyku79+R1sL4qpg4om3jADpQwh5
bLKBnJPA0IbnpUktAVbWSWDRbBKNgtipGhOD9NlNgjYTjoQGPQXgotfSbFEgGf3q1xJROTtL2q2N
aOcztQVwqjiHg+cMJdcmQ1UE4d266+778H1SDgXpH5khwpFQrgkMM78rhptc73UMUyVatxYMSOBT
mgWquW2kI1ehGiPP64hcLRdPd6BNOKtywFgcl1IadjPrfe7TKkfFjtu1H8xur5YqaM8ai0wYHq1i
dUQhYESKFRadlYxxfxTNpK9lPitegCxnv3SWgM8MqziPRVQOJEFCg0I6gK4y2OWPtFObUWu8n9sP
kGsN6wS7pydNSyH3Jpkt7viHzVdIv9fVLRXGw/2UD59OQWcWDHl1ADyvzhxSb83jOtXulVR/82RS
1JGcXQVm+x3CG4fkCcGI3TMKAMKTFLcyoyjIdi204P9GQJ7sVV6GNJ3SxP/u1IgXsCC7Yo2ne8Vo
evp0CCqykcX9CRzVa81LbPUDOUb59zbGAR+RoWP3Vugz+TDfUUePEwLIkvsJP842ob+en67xvJjw
X9oTjYWQC/ivRUdDgK5WNiI7CZUJj3yiVZC0e/eW/W/AT0YdoFyUOnFIc+xTc0Tks4eW0TdOPBkN
P6uJkukoY5e2F8/fBp/Yuuey7er8sMG86N0Un2ebJ+/76zNQ9gVmWjK1tFhFyU2yhkelV/oo61Ol
+rDazhUeaQxr6JBPBf7djY+lYOvYb09XS+T65uiZtxD93po/zlPFye4cvxZxEI7BXvScLj10m7fw
SAfYiKyhDcctlSAMHqSWAyQmfn/5hg95vanxt2Rpmc+EX3yw31BJS7RFdz+z2Dur+tVm8ykvqxwk
9wQdDgAAjM8kc5RiXqescgogQotsmLL3DnvsHlJuJd84Ki9KxFM4g+EbyEPQ5eA1xvVw4OcPIhDE
0UupjoA1989IAg4Ob70FigbN2sbTaJ59JGyAkopyms+2P8kbHRyeBJbdj5y/RpS5znomSy4PSQmR
36b3hrxfiA1bPaO1emSe83jnPLQK2cT7hqrsD0O1JIAAaxo52wD8Hub4EVyoPM6xPgw3QuBVJU8N
8uYzb4iebWT2RhBkWb6byEyLGZyBsx8DQ9GSEOjoyI67GW9u05prkD6ub25W6eLqPwze+iT1OLWQ
yLjcOKapMRytlTKJyYvMcepYCuvp76kQzNkOzjSZtWO2+L+bBbdhRpzogdkH9UudAZDC+yNuLpzW
csjc0pNh3ut2oFYGMH8KFaKYDKaU5lzO/vPLSkpq6jmX+F01zYuewarMJzojJDSHQ7Mnv8YsJtkb
XZhs32GpeCkfmuz+GkhK8VRhA3pxoGbShh96PgqJjylrT6V7gQI1NX0moBw4eVU9LDRUFI4NLZiW
rficA55Hr6ZWdhLWwYpwdz8thecF0nxnaLiixREeZ/P7j2YLsHOopw5MnK3yAKOACi4Nv9G3QrGp
75qQAgBxXdsc2Ky3wZbfcbzO6y87ZTeJmy765FutIVI3KRku7OCG2ST96E8NoHXyVtuPu4GsQxWr
WBWdvbPrKl42YqpSS40vzU+oFCKGuYaB1oQX1O3r+GvwkM75CFFpWW+s81X8BTOHsXblHF+b1Yjo
CsRN83jkH4IAAyL59fvIcPVKyfTvKUjFjRkE3zodXk7nUTNARLZUsUYjmEewLwsb7y1X65Zz7f9h
UxqzFh0d22pq+RcfAhkMonUR01JikpbX8OZ4MDn7dOs1FhE1Nnxso+VOYFLrCcrFIii8ajdDFW8F
5KgW6tFDUn9qqqbpzm1GSc6NRYTI+Nt0miXiVY4qXsShR8pfWnTK6ARds2ZkEtKGpnPbbYg/xKu4
q3jixB9au7Sf846buyDMSHrbHfuzhgan6VJ2hTl9GRyH1BZl+zwc5NsEKb6DUP1+qbT6cDvc1US7
U/PiOcimLWM6k+zZ6HIlai89J6O+i3AjTrflqkneNTJduyyj7eKwj/JJ1H7sp9tiyIDGAzc2+VVw
8xH5Qj2j2/g3v2Y9quFjS+vrfWrfc7qQUXApUQQx0RZCD7NpjDRjh3a3RonF17rbidgTubDLAzbe
HfSR8T6B/OC7sUNualP3L3ivd85tx81NLuUvWg7f0sqkDBryqT0X0QN35wCpnzVDi9mms7fMwM2t
8t054VPfuZIGA6cDvS1h99GO9LhrZSbLg57N2zFzNSAk28Ts0rcnmdbmN7Y6zEo/LuZt/1HO60Au
bqQ/uGHjocJSo6x4WYklkAvTrU+fyGsI8pq4SJhmgUo8OFxUBdh18JSFv04BWYVbTkWl0p9rMcge
4Phbr5E3ftlIgUFjvKdekw9egS2kbUluTNSlV8sUjDYZHXmxxT47leJY91TkVjbWwO46sQlIGe26
azMOqyawYCMiSBxW9SxftakjC/WpMgFNy5ID8IT/W+TMhANxnCgQeHeZZ1/XTprgqPBeF6cScj22
PNySfbyIOPC8z9V1LLsNBdUZ4JX/X8dccLqg9gdQqzE2TeZvvm3tJ5HNvbdTbGWaMPamANpH4awJ
3KnWt6giIvuK8HBVyo1nhIezoRYUCaDCx6xPfZ2YioZ5wDAIQxniYpr6CVRuIoSeZXgqhN+7qzGw
d8+13iL0CBFBRVvDbGErd44ywPgpdl3lkXhh/Aa3w9a3XupalMBnQS+BxVlgJnMBAOFCBXzTFoqj
iICbbhzZAuPYp1PP2bOXMVhIux1WBzXzURT0BlTDDA8Jwkwa4E004FqgmKPwM+74+MAIk6mgEg6h
Acq8redsdcCMFeks/lfdggo7abuCKGXC4UKHDLIZ5cjpd0/oKxvo0m3orhR9Ud2X1rTTzajxGIwF
CVStQbVn5KX+OpDa88NTs71Rf9R0G3w7vffsMTExTVrLaKu1TP36Nwtv8i49tPMO26Umkyz7KRVH
+rAqo9HoqGorGQ6lWOgD8RUZM2fPpk5ewdneC5wC7nQvxKEY2UThqZDgIhj9tNvDBTCQIdLAQTnn
ju/61OMwQ+EqkkihKxi0apR8tds6KdLdcCY+F7tzZCFLJtlrWo/fh5PzVam5kJ3ry2+ACEKPZBg8
t4EKVGgVaxVMnW9XNb3rpYawWcUojjoHiy+7XvwuA1ZReIS5dvnZYty98SaMX2tODrYJvaDWKQNV
UeaMWQOsKGWgIwTJuBnhFJXcwq+9Up5eBsH8AuYIkBtTLUV3WpHwQ4THNdHoyLagiyqDc3g1McNL
c7L8zoDI3RvWlm3578Ebfl9hBRLk6OoSMeMvPZlvFu4H7yKTjQx8jOQYaVYdYb0OBUruMixPdsbX
d+LHIlbzMnu/BG/yqeJbZJnMGlbV0B67KKwemrFJXkMUwk2FImG6nI0QjUZp9ysAcfwGHepih/5i
dUEzL6TDWwvzjvVOactghpSDR6vTFLFw7WPvd3o2GGIk9yzwJxJLeWuYGQueQaVb0wyiVk7BgVPW
BBHQonyiRyQYI5EvlYyBACpCcyHZ4kMSayyqLKMCg7JpT3tfyeHH1CFjtTZYGnOfNMb5PcoFbscg
kJ1ta02egFknA5DIGEl40PrEkkOYOfRos2f0ljp9e/VZBW+t3+3dipY6I4ZScbBtcmxlFg6TTSoQ
UAavTKs0tpI7ejp+ec24Au0wuLMZ2attugSSjRizVmjG6MeBRqe6ozk4RgQ00oY2QZUuiV8lDZ+I
IfE5zgCi0IbWUvth8NNaZmB6iAGdhh+dYgMzFhV9ba+MvDhJr5atF048l1xwMkBp9VSgvHk9Yxyv
DXcVlsAPZGUFGB/ht8qGFTH9E4IyS9hKxb/wktAaCgUc3LYyYxcDz10CIthJT8Eo3UrqmXuko31P
OL0jyXpFkF7x/B4/kcUENUM14c0d2Sx2P8wPzT1WziLT8EcTxHl7jWknu34vnqgHbG7u/vfqTpN2
lpIKb4uUGZLNRtjDH1SFNc1VFeSmLAzSGjr/WKiVicdY2VVvYWY0FYcbLVLRa5xVYEwywiF5wgB2
dvvkCLT6jshWSCOnkb081QA2jK6Ly+BO+eiEoXvK+GQ17eOOkBvWJnp0QqY2TPLCnyenVngasyac
C10g0Kss0n2d5EVv65wrArHHDLEI3vcLdmDD4xzKTLOrpO7S6+7ZBux1z8OJO4vP3YOb6T1kU8Pv
Jq7JFIVaTqQWLWza/JkT2IKRNt7Jk0W+BnUoa9fTtUXD2IhdI4swEWycHOhpfJHiJlvo7iC1kC11
2LzN3Hjt6ToFWf5Q+v22Deqm4JnVt5TPMZQWHx8vNC49278EX/lTiYVZx37laDqGM/GDJG4Vk/cA
m307iTPvWt4N5Cbv8DPDiTiRw0cEkT2TFM3VpWcBEqT3JcLXweQoebh7xALOJlcc+ePZf+vadYlV
Iv0glUimYmkGQ5maSrd5Z3PmTZ1eBKpS97yVQWVc0BZbmD86uxmmUdlX7EUd71qkmB43AcZTX9CN
Tpds5GogMreZMsF8uRbsIiMu8Fcd+8eJZ398zFsBqF5FII2BVgHyHfk2yNnQMdlQLaQapLw1cHcz
EDIH65/yeSoADY6TE+UPftvU/M0gSihlSuP8P/AmM3GFomOjlFTqCK6yhWTU4RsBU4+HqMipBGs5
FjRx5dOPSHuKx940oTHVter1DqrTXEmQeps4Wsk7VTKofR2p9fgkVOtWhWpKmTN/O0ZgPzp1n+Gh
sW78JXFRj2ao2lUmFh/oqNiMPJRSorLtOXHyytvchunUQN2Z/kujOXDFnNWiS2FUiEiG7I8UnYF4
PkvbNBfIih2QuCFTxi1kaw+NKcWRLeyLJlf+BE4bXqOqft+2zCaESHxATFIFz3xW1j/+J3VvK6+l
opdP8H6Olr9tdElFoB6Ym8nr8g1QuI7Z83LRSG7rOgt42BVcPoRyGSYSxEDBg8/AxryyfkPLOTaS
CsXiYazl/BUgQ5+OFuP9OUZruJjj8Z93Z3DkEGyRmnFyvcxYbjNt9Hf5BxJw9CtVX01vVdb+Uxdh
jEQM3povyC87Za/R8LFGMnFKZmxwhRkmsU1J9hB4aeC67C67ARQEBuTVLwWM4p+XhVcWlqm0u0pr
3fyfF2YSUk7AsGJl1OcpljJRwfvIjzdrhAU0g7kSQAlPNXSYnNZdwhFi6mJpiSbgSD1Y6QWRrePL
szDLLOkgrj1pCLy4Cagojz9UbJIe9ww1s2r7NDrtVT9lh9FZDzz/GRlCOP7HrbvCO97IwBnoqo42
y3DaHvygSpi4vqSlTjqUauiH/yBO42tAzVxU6Hff0FAq8PK6VMUFR7o8DF8JM/esevZt4cQKQCrK
2LizxOHxEx9m/5UUhlZOmeJAkOVUt0spoiwtYtkftJjH2fyJDaT3l0WoNYNA7BQ8jyMfYAQtkiIf
lbgRyUuLq+J2IACRjLbPvU03FaTgbe3wPa9y1kp+6j7C/CIS+pb8H87/hJaUk7bXL8Jm7SLvsFOs
3r00khCnjk9cE6mXfo4aO/DyL+ws2PizYOmwdiD4oAzuIUYZWr8vw67/vXcpPXeIKzd5UYx4o3CD
Bn7EwxsU6wYjJImdjdwdY0INci8Jr7cHh/mjqnqfOGIECAW34+O582ndtYUHHdpqaTJfo6PQRFkS
D7+31lzb8HkPUlRMzwBEAt0E/HLE8f+f/sSPWfXX0xd/MrjP53S4ARtIqESGiETtNUwxpGj4XLg/
tzOR1v3gnIPPcPIXuEPYSxDsiVAMIw+0XWLOLpvuCH6w0kRTURvaR2Eh0DTz33PleKZWN3DEmGNC
38/7BVnoTldhXGzmrXNJIgGRT4Y4Tf+XSzTDz1TZPVfEeNQ3j9FL56aKrk+6P3RGnfpE4UmjWsc1
FP8rv9UerZkcZKsaDcryQcrXKt02LnQoKndPGkrCpd57neC/1eL+N84gcKQt4H2Uhq0r1ViHbUgu
g5DYPWyu+fzqt/YiIEpheF+Up768weJPvB4+XKEc3qPogTGOYqNuabRMCJ8EfNWbXocHaRexlE1d
E5dQK+C/pe7c/InkWQvZWta/ErTtfeWfMKEQsdL5qgWe+PQMx2pnKJBvvL9ZvsAFK8pdsA2dHHv5
6uw/COAd/LUdQ7hinQwBes7EQ1EK+HSbmVeTcP5X5xEOfhSAFC1bHPaCZySpoH/9GuHqqGo/PT5g
WeIA4IDD8XdjDZMYj4r5h5R20VJfiqFBbl3roZOlG0QwkVQcTlh7NYRwDCKXnm6UK0lJ356W79wu
1tiASv7phJ+n0fGqL/sXHoPf3t0r1wIsYlyj590wJEuqtU1tM1ptMdOU3BVlt1QALlxEeKdD7XRi
HEyxvoLUeu9u06OIJl6z+6rcuJUAoTWBonOcYhN0V79qg9GZS+izncpEb5lybMJbThFREXe+PZGE
GGlfUcrFo0Pio7oRTNbtB+ZHoCcXnx5sXKd3HXUoLo/hB9UXxSickOHQu6/BatLY0Nz6xNcJYmiD
M1YASP1cg28vbQ7ccK6wMmbawwlt2U/DWbc6dauC0VbeJ3vzufsYqrTNUm8azqFZ5WJ5uYkyFQoM
eiGAimJpXrCutwpQqT26NZPzBEENZxufq+/J4ZgekoPPzlK9hVgXJ09/8MkqApoGM5hOTvNkeAQ0
pxEcB61kr7PPlp+F9Be9m9II2Tq0vPGyJH4qSK/A8VdglPOo3aKQwlqKokzz+LP6YWSQJ4hRX+gT
8NMw5L6hZcDzS2x73Ngs+IbLav3+3y+Bp73WeZaJVz+ZLFGjEZN8ybxdj6w26SaN0qZ6knMNJClL
YaHuxSGBBORGM/wmb6bMEDUfUPzPPzzU1pJoAC04DBTjddYoEkeEwRqlcTL/Ud2u3JlJLslVlVSg
LwG0YBHkkFSF78/ZIgcz4NhD1yEla3oihh8GyIO7vEOEspJhep4JiK/WRh7wtzTo6MWtSBuul8hc
ZYIf6l5yrwxTP1vnCF5llUhsGLrc2pm6//9o1LO4F6W9BQNCeijPhoF8QMpiyBYKhYYRYhUp5m3L
ha3/FjzXmu1TwP4/eMgCNJrSE4Z9zP03K5aMiFmsGdvhEUTQb5UOhflBjuqWp/svjrzvfqc0IiHu
O1w0HJ6CDxbq4z6rXygy5R+M2LKRBZSwyGRGf8DQi1EU53SQ1uWRf+bR/KWAyG0/iW/pG/Nz43Qz
UajGsW8KJQ9OiNx83DVVTlhO6dyijwc11Ao5rwY0LJJq/C4ZlOpmIBDM1nXOSU8+i1wzvaP031Xa
dDPdnQ1Ti16gQpXNVCvR74n/Llt+6i9ehQW/19Fp5R5ZILjicd+qi5OBrSIW+N3kzmse91FKHMyT
HedLhEr6cXHWXBu+UuapITDszwYmyM+wNjh8STLd1wBNfJFwCWON2SF7BPrtlBL7IEXZ6UyCg2gD
ENRYPona4YTR1qNe9l9Dz7kHDPqYaCm4PgnoU3Y79Zndb52k/2xRTHhBHTWMutZwIjSc9Qg90iEO
tXRPgSC15e5gAShF3tJ281M5Tw7vRB1qOGW8jpyz4dLtlJFLO7CmcO+zAttf2kSmhfG0yaz/v5/L
lGFOhtNFdd+gB3i6fKbMBmFjqCMJ9TKleAtpNYNKUTNTU0WQv3Y/IaubYlD0OBGjhpXPJXo6sEmt
xWo3q9Fqc9uK4apbYSGy+ROy+vC8JIyk6b3/7+ecn3qy10V1rkm3Ywa9/xrTO6hvWZn/Y6bpFtnu
I5Pe1jcgnzCLNU5BTsyaMiLxGQp0WR4xjzcL3AUxx3/UTCblFQNHqYTEqsxnGfQFu/Wj6tozVVir
gYS8O3l5TdoUhCdgf9huPCPMPGXu9yelBZcMOsTI3PKoOx98kGUn17MKijgODoOxIjHz4Tf79fx7
Y8vz25a5+O1vQrdZewiL2h0k9paQuTi9vqjZXinrJxA2/M1kmo+yLEVGLLU5ZfsyCQzOadejo40k
w7J++ps2Lku4v/JOTYOtrn9TiLqgL6lUJr4wVqzdap6sFltVA7thsC42U/1859txZ/12reKhRHo+
r6QGkONobUsqu20rYdGbrW8LOpJw+O0JKpnZcYaGjAzAUIwMdGUJ7Zqjer16/+aYyVmFkVEzM2wh
OzSl8vm4oygYNUTAfd8XI0jdkzlQC++QQhp77YUHInt7mxPAhxpkyL2CIXy2ItvCPUIRYz+oppOY
Ul0CouryavwzPdD6a8S6XbljIKuO3xj+80O1lJTiRibiWafuEe26ivdoYj4RGJE6zsCiogeL+UEO
vRu0aznkAVlk4Fe8XPVRJ3ijsP2mFcLsEorxqDzbccxr5M1AfEWsM182H0ZfK1/DswnK6jR6FHWW
dt/89zVXazs+144RStNt1BUyYxBN23Ng+jVuWgIS2HtfFuNcfphpiaGP7wzBHr6bMAEgUSUvUbL9
XF7vgVxovw2YAVdZnDv+Cg6rUAOIT7NtzMfc8GipOHvKHSf3CrpfG7YMsDC7tfBVtXNzq5EYmtop
TdVvjn0/0vMXaKuhz6Ia5bQ5CmoPMjH9KaHKnW7yIOrfSlXaMiGJkrNRyIl3B6rwvjQ4pBrZttBw
+KdtkSr9hJQs/DS/0m6PpQn68bj/0aEpX6ksmUushUfg8JIyUE39jkmTCU7iD417vF2ySUyRIcSk
Urc0Bqwcx5mr0muY3PL9b+lBPlRQS39E0CjN7rI84DoP4moZ6RIhHlqv4a4LIJof6hxGTM2CTyMJ
30lDWlIB7tu5EKg7a8XG9aRo3frFBIbkS/X+oaTOCh3+dBJO69u7x0wcRXSQcbEI7qTLdSiXoC6j
LCfOZLN01fhFIa8v6IeG3fzxgp5gCCwFHjdv9A3RVBhbMC93RaPNtZVz72JrRjwTX4c4Tx7BQfkL
iC8on6cuca4zAy5mtJ8mJIvUUJVdH+fR8DUiESFV3/mrEGJKC+8OhLAImweQLlzSzieO3ReSXIKn
Qbw1H2z8drMbrb9Bd2bMMYjT6PR5I7RuUsTDVYZtzw1iUC1HZvL6h7YcTTPyOAmiqe4EdqWHLevg
CoAwe90H3D2PkhzdOmfMH1vs6ldLdxGZAti2640YgOblZN2f7QnyZBu3w88S3gHZXc9z6lziLGFs
Skrlsn0GCFYnND8IFXtS+a3sB0gUZ+L6o0LmZvg7g1bEu8Mbt2QMoQapKDNXj+tDYJPY+fNB0K07
4Fn1xYWaFGpgNlwvftUooiQMz3xdfuXfXo4o2s5JaOTpY8hrPdVaM9XS6wRx+7/ADjpH+leYMgIJ
rbtTQzLiqhp/rugB16vKRVFV3DNRmMETVBUnOC6Oi8y5lEyZ/qmbJkinkXBtnn//e90hbZ4OKCi/
dizMs24GbTlQo+m9RYbGXizci+Beqh1ogWDrs/L0VNAYFSdIZxJHXI+fRrNi7uCcZ6wTZsNiL/SI
0Y2Wro41E/Nl/FdlIqWjFVGvESXBW7CUgp+zlVXCzrmXnUr0kQ3mczIQAbY1TW8ADEW6GAS52x/n
9txaq3WNTq/zChWpKaVVQ13G84v9FTvLXp/zqT79VchVi6eFbD3jet8zLxBOXkxgWBNY2G3L83vM
6xNXpnYcJmYje35xgaI+OJx6IFgdS2NYRIu6RU4e29ThvmGN8oyf573pwjmsekcN7tTOO5p8wTLf
SQDw9frZdwGnACMANbr0oxJtiFDNtZquaekbFfbNj9sauak9MM4MvvCH+9W+/MhvrE5IuUapXqtQ
+BuCvNJ/LmuYQQUHYQ8uywcAh2TcaB4hPfEtxWeYxH83Q8Z3DjhfO/RO6JvyyHmK5zfeF0sBHInV
IsSLwpKes+WtvxSHkIOo8VP6NHwhh51JXnAZWyLkyJjSVrOZ4cdoEpizGPbiQI7X68Fzi9p9Kj1f
jI0wSckDOQ/o9q1uohs/T6Qxc93hL4Pc29BUMtppfDiMgXW6Li4XYD6+y4oywIvvbNVAbNxzUHV1
p6gTiVFM0szb+K+7ztWJf/lKdMTxRMnkXwGjfJuP5Ay1ZJmAinCVV8IIFYXcNpl2ga9oGgBa5NGw
vbovIaJrSz69y9n0LK2v8QmhDqb7Do9w/teU3nCPZL8cXzeO784S020nGdPC677Lnl//1mjX0BP2
DlZC7s9k8yHOi+1/xe2Z3MnDU67wqgTW4b6wHhDAE3NYzah0m1C0B0UhUJyyMqr6tmWCaVSffJo1
CABOtEU3hB8Kpy3qrx4LFizM/nncYLV1nKkHsv2oIY219o7rJi1SVL476ZBk2P5fgqUdypsceHMS
slS3z+t4UNyWRjvvp13s6pRInBM281wsXOQRTcSmjNCss/rIpiykr450uJwTyEWT7eDaJVx4BYBj
ZrjGTv70fxi4kOB9YZChZCwu9USn5IcJ2EG26WqXNvfjfJ+xUcrEMcTwiYCAg+aZfQFw9G+b8C36
qbFZ8QscQU4bjLoErBbvcEOHHWLAI1gZly++3izyw5V6DtwWW021MCJ6Do0YoDkEnTtaGsu8wIBw
iCBoY5fFMMWHzKs9zWR7fUnIlPJFs1NxJ0PfVB6KRik2rdEH7+eOPPUusFQp0YCT3xka/MqsLaSw
ORsER7f0GqMpq6eeGo5wbLXClZUYDTuirEeh+L91fOJs8CEpJ8vSf3s8tWkitukiBEe1pb99eMTH
fbmM+SZpdpRlaUvTyu2l/BH7vkB2OEbO9Al7QwiNsoJFM/Dq8UCiaLOEKkEbADKb8uVv8dNjVwxN
0ak5rAPcKmgIJndIaZi+ju/V0KoUw2TvDYGt064ty8HHQ8GdcEj0hGN18HpR5aoV5M86gH++0vkD
wsqdKphU5zllvvrgSiOrVxYCaKyF/RDFk5w4EYyh4RYUtRZxhUsRrMakXb6Ej6aNYfk/xroBg65y
lGCTF9RX5myow01fQ+v3h0VhMQcYTVr4oLUNrsZFuD23wFez7n7VRX3d9T3OROZO9M0OqNhrDeQL
F8bX2gyh/JZyjnFu4asaXHAMymXOt6JkvYbgfsHlHqb5f4HdSq9iJprk8eaZVTd74tVPyghRkep7
hC6LrJLG5FbSytn/e+syR1KtAP9no7l9DWpgYNWzwEXh0b+S9SeguoP3eG992y9xdr15dBygB1Bv
00coxEhDA4t/XRFGeF22b/cCJk/LqfsRVgGYRC4BdFpPM7mMYnAS22DjXFg8HxCPKHXQiWiAdlK0
seXHWlTkZQivOD91CFq+xFA+vg6reUDaypppO9sxoUlIdCI8qklOIfwEuzcxAN67lM0IiKd1PKFZ
khNZOZ7BN8aCcwa5epw3+t9lunVe1m78Nq4klQs/5/BksnutRHAbbjmDTjKCZ6Tb5SM7ngbets4k
HzezmOFoMrDG83CvraWjswRTuLddAd+gQ+hdvuj1DNPEbLD2PggebDK6+o7BXgaY1k4jM2l9wFJ3
vMqGHd1tXzFt2qEZPcaF/CJ6mUNWvObuCkFLQT3cB8G/T/92YymiPFVCd3vnmNRbAAgnbPAbAEVa
5c2EQfIHcdqAdKqdPPVzx/B+tIkVgiGAQHe+QcZbhITfwFAHuReTfa7gdlnuToHGOojFjyiAxzVn
1U10URcrHYCFI36J94MDhjctBoff/aEQoaUhlVc5KjjPFhuis3XnI2N13CN8tQW+Pomh2ITZ2lqU
UFyXRev7aXpYwIt0WD1DtvKImeOYxWeeaA+jmUWXwHbhFmlxCEpic6estC8hq4nqI4rcwTa1yBWb
g5joSDEAOzm91A4CXPKr+MvRimiXoBz4aPPSvMcz9F3Rz+8z3y0hRGfoyw9XwH+YpcssSYp0BzRj
gPQkUo0fkLre1KxZSjYWuk1BPFzGWy9RYxm6gpZpXeOmzwXesjzNX1QJUvXtPplR/13Ztav+fSoj
BxxVYqPRYh4ueElTZLXjC/yoedQnLtmOnPgK2Kw5+yMi56/0uSz1IYqnmBSrwMEFEXVBBilvY4nM
z420kXqNHnfcoXWaHWJDMxoO90ym5v0jahYA2xGmWE7l2SQS1ZNEFWlCyEzltCJNY8Eqe/7bYroV
fr9uozbpKJKIJdBbDXqrnS3Ok9rWdbN9wA1R96rtPW7Lw/pvpsQKHleB6gu0GeLUDbVCHIG2NY27
DfdqHat0W4Mg5Q/DhWvzkR9z1Fdefyeoj/2XsGsyZdMVLJOZEKXQ7pNJR98NAXbKDlpksPt5tFmo
uiXi8+Z/+R/d+PvkuydIUv9dt68Aghbr895zl5Go2CGiVSWh+SqS3wZ3ZTZoXneN6JJEdXNoG8+p
CD7Ls8vN/yNLqqJdr4Bm3DDPen/jfS98nu7LWUrS9TMhlEWl3fWilRI2CcFZas9aCJueMVVpNJ2b
HULRcdB6yANtnMhPrx4vN99dxNU5f51qU1a0zPAjSuy2z9rfnpG56J14bvGf6Thc1Cc4RCoqQbs+
T8cq0FWfTTugzSjuIn9K7W06nc12pvDdG0zRUFS5N+5dMUkwyWyVVwCMTu+kEYcA+rzMeOcxVPzf
DYo3yEocSTmS3t1k2I+de733IM48/3HO3Y3y/oOeW4BRcqQURlOuLMX1z1av0Ww4xYBEnSWCWqAo
4a5kwh6CQ0Aq4mQnPV+Bh+WYeJCIP14BXeJLpZF0YPwcoc73ynQVIxDfjKjL4NZyqSBnodgKJcZI
yiSb5cjiF0oY2FHctjFY7dTS9ZzKToOIg/6yhHEL/vu6a4lrFy9WKTN5QM4DTFETzxPXF3/LrX+5
/eEElttR1HUN2YX2IMlTBie8IzUuWkx+6+B9Z7j5IwavsxWFwHw8vu4OV9/F84+CMskMZBc5YLFw
xnVkn7qHeboNpfi00i4O9uN7TETDtXKyWcU34kas4D7V0ikwIKSUmlteDIqVmbxofGY0B8Zscy4A
D1wUk7OeCzWJ5nsNUryW6PmorA+5q00LlQ2OF5l+OOFP+tiTLnbICb3HOB3ybJaYDFnym6xaez4b
C9kVJqypOJ0yLm7ZIKfS8OG5DadZ9xmZl8RwUPTZXnYmxpOKJ3l9fbX2r53meqSeuGA3C3e/SeIO
JgH5UragJxRDLI0ukSU/ZZes9hSecSG8FpNrdR4ytNIvHI9pRAqGf1aT+E5fLf2hFZbU4L97OtVd
5Cmkrf0SeKnOMmkQeqLO/nzV5BSvYZqZvi7Afye97mFZ7OObgFc2y6sSmucEM8mZj3l/VHrYO48F
iMdexj53MR8PQtQshilorWjzw8H6JVTrHSKittA81//n3BpxlrEVoaohARrnONRRUp59Aq1A5veM
iVkcL/3aGVUXYJEZvLaWpcPuYyIuo2JBjpvKqOooLtxcQWnBUxMXt3Frqy6Wz1cCyLanHamnQItt
7InyqO27nTs0gId7XT0yMZdasSAyJg/8J6RDt6mtQ3MBG6nfY2UjRSjnBbak4IMt78bUEYdkUfl+
Mu82u5GjBTO1D2wTdCoSFhqhZ/oda3mV2mo1Rm8dmWtio+5Nsw3KJ1QEjF7iVV+dvAR3He+1GTNq
WxKD+hAIbbchse7VOhNZ9qblXJhiLuxer94RSqshsNCw2tB2UVBQTY8U2mZDQ1AqirGnHkRIht3i
WBI5Sv1PRgRspKdLjcEOCjkhdSJhObJPZuqu4gIVTcRK7puJ8NgJceRnwgoO/BnWebxZzne7ef9s
x+mTfNSPJmNvqoMOai4v6Uc3hpbyw9ZTuIM9AwdwUjQlq+0xSdt0Zc8dOPj28ZN5QS8jnhC7a7Tj
8MPsk+GlTubuB7+mO0suCOiMmN3eg9BBIsm78KDLac/ueHLQlV0WnzKdb077F4in4P82lSbxeVtD
uj7ZRxGofuEnUe4dy0g0HIF5mu/vvkqUud79QOLawayXnR8vMNreDll05/ZOjNZve+3DJXwa9m0x
1oJrjEWZNaWr72coNQ8gwB/4JXlgYIu9ACJoijLBJA2Aj8tk+bwokinuTJFBtbNxOtZhDm/Ykb+x
jP6tNI5cceShrOnCaCX6GJNz+X0w6KqM7ifa9Qrm4/W1jxDSjvDiY1AoweTtK/vCH6cru+lblGDX
FnoycnzlUL2nwLpjavQf/+0rroOwE0+uGBSUAGFl6BLy76Hapq/y8tS8rPZa+sRkyALqg8nepcqi
PaLoDye32guRGBDWsldQbl1zYVd7k+CSvSiSYidiyYqmOCvJU3pheTQ3NDOJt/Z+R8SvRLN5Wffl
7g0hjbByyD+ulnqUJKxB5u1TUYbTcbBvMD/jTSK91WG5tgIeN5qP2S1Ss8j/FiMxePuSa3YwV1wD
RecTIogY7whrnSOiyxxCXvG3XnsAoJ2k6+Huy/IXZQL/Nej/NSWGNVzDFmPsDFFqzQzPah6zmSr4
1/FNNJn46onH06N/AouExfU4DzAVOdAdsv4cqvohXatxjgQr40UFO6ikjP8EMKRr8W7DYdfAYezC
86syDOdZt+gwLe+TElje7xAukYesSblxFIqokubVDH0mN2ZvsaEBAMea/fsZSTyWZtYQnlaMSJWB
aRnXQlrYeQaEz5HoSi5Bb++2QrzXN/MjSJx6soo0IJ1VdRXw8vFqvFnkFd2M2M+SPX8YoRdTvfln
sq3e7v8zGVl/AvGUy5MM7GlO3j84Q4hzvnH9lTFnp8poFiWSdxNGGXrWt3uRnKO37tT/IstwpKUB
I0oi9AeUt9Pw7QUIa5HrF70jWKmiVfqx0TGsQnwXaZ1yVpu9roN5djpeXQNG1qSNcT8Ch6s1sGZY
s2crdanMPNT8PeGFJxT4dAFdAUeE/1OIsDtCqyPDDZWo39s/bgGoUX2ZKkJ0BB8vvEo/GsZYU5TP
7dyJXPOZWkFqTJdvrOQooUWoYmKVq/XvXesNxGe6WfMTDlMOSpnl9Yv+bWeCEocyHG2lb0aGbYw/
awayo5D19omP5Q0feDc/ktq9p+bsxhTc2DtQRRB8f4Vxz2JIXYBd4QD+0LqmsS+7wGrtngCxRPNs
S5OKYVt79AQFjEkJPvrQ7yfbz3pEQ244NcmA1X5n3x9czuA/iyblGlhD1RAql5ojK/lhPyPJKczX
Iw2RdgxW23QYgCp08ELl5n04eiTDwGwiItKzXK79RoK+ZlCn1T4NuQJNfXWRLYkRgzpc6b5GSLS6
y0SzHKKYFmMjT+URnp1HqeoMU9AqWhA4y+tnY9JrT576ONbu9bd1lLb9VzRk7JBrCcy4S+vDnJLT
1rwpse39Rks/9S3wxNQtSpdtEjXOcIatX2FSNMBBcgM5oQhP9YzqnAHX2RKPGkPmznpZQMUl7GOW
ngMLjaAJwGTDbMt4I31FWd01bkqesNhCnJIvd1aXnfOG4HgbL6/o4a4c6Xubo/Q2pfL9LgxC1GwZ
jtFIfPw/VgbAaNKbQT4+CXrlwgTmO6vihPmZBhqpH+hN/KCl7J7+AytqGY2PmytjZzC9XjIXvjNF
pnNj8U+RjJa4wzxi6UdNWE7C70bcmdHbkXRzCdzj334HwR+w/jmN+To5zDrHv7WilG/v+cSJCqJ9
Ki/ms34LFSvgEYZ1gR/H1y0oT0OhJfrch0Mv4BxIa1LfsMSpi+kyQ+4gk7ZJdii2lIhcJmAtFnSd
e7+ajrdJBQhVak3jwdPL7B09zqyJza3L01Pw43cptqDOJ3z7kFHiO2NU75e2HV/SLx3RIiNae54I
355SANuGgR+DMEf1kuCp6pRIMH2hkodjGdPN00Lm3/neQj18oS8VRqcq5yEwodagT/y24cVMFaav
mNiAz4y23pDnJWh/N7L/flB4wWFnv5Sn7n5nz6FOyUTXI8/4Qux0KhtsW/57rHbqcnlunHnyMSSx
ebxg5VRPc6KYgsYNhnNnVGT1MT8cFBJSaXIbwDMrc9lAXjp3cgTOUxbZodUdo2aUQB2b9XfTeUIu
BA6egQwb1AFBaKD94ER2gvtZXoma6jqL/JGE+i4z9Xj1dMSKdVGNXs4URjbo23PdVaimQP3yhxe4
qhhb4aD2YkWqIEF3mS+Ok0MBXHLG83WhpCnl9x5aui1KusfFCWNdOLLBawXxajX+HGDjdmjr1MP3
PD8MtQdHYDAhLmESyecMtr0F5vXT2FlFj7ROXJFhxeD0XXdobMaLzg2unC20/3MBWJJD/cGQLEFi
PEZJJw0DEz2sT1mpymbms565lcM0YTwn2ju7NFoK6TCwdG0m5ZK0wPHR84n3zVPueb4niHIMVpob
IMWesm697eyrz/MjDhUk2Nrl0C3B+ZDngXmLAc1Kj33RniVrILTJkMxo5Ag1C+Qlj7W5QOkKhGr7
2qHAXKDL8fCC32e2KoR/1gmAhlPvqMaNSyx1aBrZBYfvuaw1u1Se1FdyB9R34nb19ywwTWi7oXop
PXeNY3v5rQfxn3VZNgBS/pVW+QgKyhCqva9/K4rscLMEhgnKLWwJx/eiXAI+/9A9M/Nx9oAhXE9O
6EwSlRjmHd/GmzpuyWzy6bR0qZZ1RKjvYRH2/Cx2ZveqIwe7YrNWnnehcbFTtGeYJDzjc0Ge+jrn
dAsHSPOW4ba53R3q6yfivVLDAYVcjzwwrD8n7VxSbOT17Arz75wJ+55k/1ks9K/rtV1nx+zPHIeE
pD556RHqSL9A6AYi7ISwvtsQx2DZgVLHZxdKkowrIxSYiGM1KPOA9l+0I+yF52u73PBN9ZByKGoO
HljVI0CcDz20mQqRJReWrPtUmNKYXwY+S6o5sqmZzwmBdIOM8x2Xj6IvCxz4QqAvJUB8Lu4YYZIP
4rcnthYE2eDjIy5QreOf+JaVnGPhOv4TbPbrp0CQ8JDWf+AMhRIyz3wzm1thw2Aa4OVSOdJ6w8U+
xdzAqc21Prr9B2tOsfPG50Qzt3gIcF+cmnqUHlNJ5ew0OVmp4ydOvSqdytBzy8NvnYdP+EOw78AN
oTcgp1xAM13Qs2FFG6bAa4cKPvOxAZ3zRmjumuyU76yI5EsVqOhTuezthVpOdCaGU+ME+hZC3POO
TNcMKLKisCJOi1SmpHDoT7MLslr2ItpRGffQ4+O2BV5ghj68UQHr0gOCsP3z/OZKQGI/cbmY0thG
DvuUxlmFfMnqZd43Kf2ZVc9t08gBFpDX6Ww0Gp9cb289b46Hv7z6Npag8cCMTbznnblwr0IMGVsZ
mWUJ1DcjqMUC/hL7oy2S8KMr3wuizrg2CPt1dQIvXG0zkVzt+aXWZpMkUtjPj4/9l+QAu20MvZzk
lI+xmISwXhS9oKzpk7Im13P4UQyMl4k/dl4RjezJ/9LSz7fff/IOs33NoJNoYQrx1J4LmJUUigTt
QKQN+DeskYi7hRjeGr/zpIFI/zWH4DsgOXbdYOkgUHu3XOVlVuqe/GBQMf0PxHw7CyUnWB68hrDY
PxgHzEvAbOsItwwqRnAFV/y2eTqOmBXRcsNjgGJXkan8HTqqVCvNXPG3p0jlTisXDEZgEp1FkDAD
YZ+vOpMZ/AefpbyVcgrICjRSNINqZ7gmjHJP6BjRD+GmRMPkLUycVwrqx5JSmDDOLGAxIRmarzjP
73Gvh+9w0DHk3c0iJZCeIZ9UYMq22oCw42m/iy5XMXAxUpm+4Hrw4CIlnFKJmRUcF5cSudn/Jku5
B7TZ4whuDbQpMBwA8oupPcjrUx5hUiY8U+EhU8UIdCttD0UD6KBv1TqcS+UQkMym6Gt/mmW+VPwb
gVCIGXQD16CB8FMkQOIYEuAtT8dD5pic1XkJ5HFUGeXp/T+TAjVvME0bqd6Lm1apZbNndlIkfrEY
yoQVKxeUtNYHHQyZY1xCDBPr43td1/R48Fc8IvD4SC0UYdTPHBVQxwLjiQGUa246LpZOEjcbQzr9
wlewoI92oLmKTAr4rDdRZLkyCA6UQx/j+X/5t4nshN//ks50qfmCgoxe6hh5QNXdHpLCVkovGU1t
pdladS4x3bTl9s+CVEE+OhPF3yEuWsIZKtCWr5Lflxrq9yCB/JETzUpkYeEYC8p0sGfI0ApiLMF+
gWHZgb4mRXW2ZumfROZTLibh5HYHfsjGhl5UkZffGff7buwwiMpFbV8dUF8bNlJKDrRThxZA179o
MAnvWoh89WMN13iHgxb1A9besrqA0mMGktdyetvSZZzoY3Fe8XA2B9mmzKSnhzt0GA7sDss6QDUY
xNc3gvVsObMJpvfkwkbA+aiqP7QbY7di52br/gtDzstTWJ0qQPEygaKI9MPR6inNSY4AXZCVdx3D
F5JLOOKpulbJlTd556ntzJCVTDevgRtL5NEXXQXZeh80DBSkgbQOLiaanTiCiiglxzCf5rUKxOMF
udL52NVDFJ3VbU9n90XYwDmEEe3g9ALPbz4qc20z2mzSOBS2U+/3OFb4myhhpfTVKtkp5XIoRI4t
xHPr4uBoHprkBmMnRc6mfkJiJHvJrGX7U6UN2maR23iOd+GfMTr+dn0F1cX+rd6osQ4lDXkEO96W
QJY4oYC4Sy92dhrGQY1cA/+GQHT4je0TBIaOtzdPoxv7w/QuLXPoEG5YG1E0z2oRcwPu+RM/pjgr
6Gg1/dWUT++B8NbXPIGepa6F5bvt1Q5BkZtXcvyqVw4f8/JC1xoMOaPD++6kvjXMJ94wlGqTOVux
DoaUKr44OU6WFOI6i57W9ZYenmb8GdZsx2Ee5PMOWrPueaycc91OcrjOc4szzqBc/Wi+ClrtOvLm
N6KwmE/9csekrV/3AGo20eaptdV4+kQq55o/5j0l4xJQ1DGUgoh/aXsYsKU8aH8QwS+KBi2Hk7f/
Sei0viylMpm2ouK0pNbkv68BnzoK8gJC5ko8XxaHegCLUcvZClVcFigpwKN9iayCWqi+eXYzbTL4
02s1Ge7jnKQajcOH0PFRkk9UdqaRNtpwLzvylT8daPkhsn9Ap6NshdwHAbKnABSP6JxVL7atWY7y
fbTeaX9uSOyKv9a+umtgNbELqCr4qA/FEWc4EZ39fWHn1MHENOuxIWrX9beNJc9qVrTkSg2qjWLQ
imdx2U9uV2RKWnP03dkWCXaDuOhUowK5LUzU1XaD0Lo7+FSnlQQDZMj0rNDZZkV29wRkeP1fwmjd
IOzlKmCVW8+ZI9JoyzOrVObgNuaqm4UyT8bh7RFROPZCshU20/qGTTGWP1Cx7xa0VWxgLi/jc/4S
5rnvyyYt+4EfYEFDk2tW4FSMU8vnVK8k9Qt+Qz03OAcdnq91Jko7m4vFBDVs2bL0fWQE0D0YDZ+G
V7sZgY8F56LbwZCUyn9fQgH4SBT3ejDEIFcIs+MFyC33kQSwSN/1aiZsi7QLUSDIXi218+Wtp8fr
LO1Aj1Q539PFOOElTISeU3mwZUiihnn1rIxGx+X8uVXDWDYbPAgnkPFVp9iMwVH0RP7BL6Bsm7jx
vMUA6P4PrxC/jKxlj68Zx71gFywzUFs/pYR5XdElwFFvJiycHhcgxM+MvaUbsmtw+wSaQRrabxrH
uCU0l6SlGC8OmABApxOvjHBKS6IUQocqM0btLFZ9jIm+U4Mp39q2vKvLbwD8//z0oZ3DXHvAlNon
TGj8bQxj+HNDyAWGCbMmLC6wvYEZJi48FMiXUFAvqEKn3y0ug1k0u2SwxhzA0Nokr63WowFP0izx
HP6U06t3b2JNJScgKGuW+KK41zDE9KB4Trps5xLBI7R3jU/fvE6MrfD372LziJXJBVqXBdbLgZS6
uJcVcRLv0d2RH970L0gTh2ZseOiibtNGI6pq6rMoo3EqCrIQTnqnTDNHmKsyAC8Ic9qtBcwTRtr/
8KCRQHdkAG65Rc6SP3BjdINapH46MDcC4CvPKKqZIFtIbafIGfm5d2rfl90FDG1hHezRzJkJAXBo
7FRzP1kJFrjoHDOO2GT/RW+AsxTy8woxrNxRMQ2Sqsn/XQq9J9Yb2Khwr7Ej4ArzK7AclSBiy+bs
vuQa24U10FLBf++IvTRtp5b3j4Pv4cwdxQ+NcwCbKRqILjgPc0wlsVUZpmo2HZURZZ2dVS+jFCT0
IoZlcjTNAeuRzToBrhBjl0eFZrsnO0NuRFAK0mF42qwvSDauFIIn0QcDb+4VbZ/vIyfhVKHjZcRV
AsU7goukZeakQuLhT7z/tdrh+7ZDKyq+qOEK7G9j17xb1rQOARee6b8FdG2pUt8tIFi/+9BuHl8x
mBjP/VLEf5jD1bc+Zo5Xbq14ljJyRaibr4tAt1Ph+4KQI4ATNaonePQSrH591deSP9LbSMW1oMfL
FM1WVM9GZ8zACw7CMZu61roPEmeoFCkoZs2I4sBjn1LotYiniN9DXDKt6A/o9Q6Vhn8ZX8Vdj8o4
nJgA7tYGRpwRUMR8+aU1c6oCofMZXfO6mpZCesGsxQgIGyO559RAix2zj0H6CoA2WFfDxyR6/2Zj
Z6A7muOJ6AI6qKLc4EOV29v/u4WYETDFMzoiJr8wTiSbYqiVRzP59DZuwSZb50/oZNpHM6moVf66
BfSnOjU/JUw2uLfgQV58XpXHfHUiXgf2P1Cb0qBZsFx5JSgPKLIcV/F+lt249wEQGo6oyHw5cE3n
2si387Bkl4fTSvODT/aNxwhLylvamUMLFNUasf0IhQOO1mn5qGQyPT1ZhNuxUqbEEjn52tjMFYOj
Tbb4RbnyhUhpfk66WIiwPnSHWgmrQyUZZc7MvukjqUyE37N+ovWEU55wBTwdi2bxk2lzn5hSZFyt
ooZ7H2DrdC1wv/UjdjPO+mIj8Q5t8kCNU5yujftWlEUpbQVBI+JAV/iYP3emTBx8lGGlvZfOw7IE
Om4tJjY1s2RV7r888YgQ/JPB3uF7d9hC5IelySaiDT0ubuCWEaJBLEqMn5kSHu1Y5G7fww0wZAjq
K1iFybuMw66Fj2+Y4/QruzOYfd8bn7ICXljtxry0ZfYdme6XNG/ZQ0hzHf/N73erSvW+1QMWzUSp
CaJDKf3nbg54tPhzkj6CJejaA8ufuszDN7Q06X4/Xgup60eVJOVaANBX5VpHYHk/Y2e+t2ikShP6
mWcREiMeV/IuDhdapMISTFGGs9TKrxr6Oq2yL99eyN+vZchlaXjQy8PXv39+zUzMvPQHNvJ9oY6m
FHjoblb3F0+lhym9PP8nEPzx9MGxaX22v6d5vJ8gTz6CILneWYlom1EXyOiCP9YJNvVoVGn16S4T
PLnQHAi367wH6OM6slhzk/0g90rYZpsCVk8CK3pXokSzD3tOMWx0iV3T1s/LDEcAH3ditb+mZu2x
+5iaCxpHLB5udgr77GWwrYFoUvR8w4sbDfal5a3idMtiDxAeU4F9ZVrt2Ynt1Vqespbc8NjKd8sc
/FZZh42LllChYPETuYcETo7rgIxQHYRyBQa2E7MlJZ8LMuUzglY5Xfgfj/CgC/BHIi+gUJGAzYrG
VVUXsV4eswLrx5vFM9VpZYbX0sSkAtlzvnLy36KIhZTox7REqPDqSTbHJt/U01HbNiPpGvbBfcnw
a/EVhGaQX++KQj2IY5Cjm5PTjfZbMU4QiRHqAjWcMMlIWZWcOvRs5lMT9gu9PRonUcePVD6EYcDt
pFSKn4fKcit6MVmMkU3CDxIlwihsPd2NTWpstfIkpFgrieKy4cvNRC5Az2LVFrkAsc3XQDzJ9wzH
xu9ljDv82zVEzuTyaaECtOSFL34Z+pGE5B3WC77ybRVM+uomSykEc/8lUsbxbjX8yMxa7ELhN4fO
HcJSs1PydUaoE/odncaEyTjXZAmQmphoKzfK5WcwzFmmKjn22Hipn432vqVReDrD1OGV4vDsm8Vt
omhXeiOW9bDSlJdaP83rRxIhX7egr6a207He7yLckgMVhSmNbkZWEz5YVyw/oq+hmm5NJWJpPZXX
k1OgVIpu6FajCKzxJoc70eHlBMq9jguj9gvWaaYy6rnE+W270wr3go2AWpwFAsU50UyncphWyFHW
bGKjl4spPrmVOFxGXm9Hemwzliei7MKJ/hTgd/ZYTfUVOJDsBMrSd0qtsMnrkUKVqpE8SYuNCLXy
WyZQYsJLU1qs439CNkU714DMUKEgvQIVrJk8iFxhnGI8i2JLoK6mHhpetoHozy6NJDK3Yz8PJhLh
w0vDvR0BJDYcC3SRJ4inO2jdTf6ZB8eipugV+7jODSZIOpLWJG0fZ2LeiIPy46CnCYMZpodsRNvn
KsCCaUFAVkavDmel91vpQnyXtxoL6tzrodZ/UYL/gXjWlHKXbCvt8iXBBYti6lBxISdyMP/hnNBk
JxGu3nt+0np4E/x3wWfytht4LYj1aXw3MlDMD5NVZTbVAy+R0t1yyDEG7AgHddeHjnmjjF0h5W5t
zINjR7vuZdr1gUVYp8QvTOxP/S9WNnI6d7oI1FioWHMqmbn5nJ2ztQuz0PaWKZVoOKgs3jU2VOcH
fSmke+2gCBANElsrl0xcGcgQcdFRURojjwBMTrix6KuaNg3dvpSxGiUWSRZq03Sp+5cFLeGTcANc
054x+FPIg9yN2UVqLL6JhIa0w8p9TTddhnqu5D8iyHSUxkVYUuRc50DD8E05M7OZXop2G73e769k
mVWo3efq79p4mdvjzXkH6IKDe6aDhaEQskaa9cjWzlhCIPyby00QLzUdBfC0XkY3+Gm8aaBOR/Os
aAri35DE8UVCC6ImL32sLWF5h/9DjV2Sx8N8UbaZHXaKcoH22YAlsUopzHll3PHpX/dtWplLaimW
swZPYiNBhSGQoe2XgbbCnNuH9HkKhzDgO5EdAVZ0b1LNpai4onBe2bNJhc/p0C4J5O9lU7EpJigG
q/mIuX7VOtTiIBGQP2J2UU5vssERBoxGOrSePqbUMJ4yw9Grqer6zFbAVOBsGZVPhzwixYiCFGaP
yreNwQ5Fdfn5rybyM5pP8R0lLcMavaza46gCWGMMlA9duNiKw5AtYRohT9NmUfeaRTrE52ZS2/dS
hI8H2YUJ+Yr0PVjCA0TlXfPiSzisaZYQw/utFRKCpeLbxvA6kGU0X7jgqvQZZv3ExqC2azBKwwD9
m9HVkEhAOh4g68pvpEQ3PKRkic4vxPX6TyGBkzh5wKaRPmq2WK3gIqqIsBYvdcY/K4Re+yF6Jqc2
qZMkyiRg0lfPl7dS7URVuRJM56ewwqtaeaIiYzqrK3R20yDR7cekhT4DyNJv48mTsRL82SJc5aUp
iUDevBpdjSebqF32vt11esecHURYL0xefHsrJjcg2AYbQddf8oJTcDhLElDZkUjcMXBYpLDfNQG3
L+mYFnnZvUVOGDkNvHASaztWkuxy65B4/sJuxX/+vEWaC82OT1BTMceuC57xi4DZouvORCF4lFln
xvk/W6peFzdxSArN7hLHyzDQValVXeBK5xI7GRk2a5WTo2++2eEmFLae0QObjO1lvvgTr5/O4oZf
R4MCI5W08Jn4stLYh7Z0c2TUC+hx4PR3oW6+2BBQgJ+6A3PyZXnUcGo1Ex1z/pBkfaE5cs5+Prk5
AtaUohKjflrnlbb4XU0OvJIWUSQs5wPjmhfFbW0kVrDb0fgNZVbWeRMrD5yJeYmU2/qp/uoI1ey/
QwxusoYQMykirAcogwBFwCQRsSF90oMsyinCvXhEBuvv0nOaNxCmriztpc5c1onKYr5klAwLzl2J
hKT8T7fPnRjBCBrYWmRlta5wfvPWrh59vfpbOsc1EYMWXYpJz/H6QKLKoBiQnPv+e/acNONGvR87
viFLFNYPnZv3lER5jGkLtKFnUUUKH/a0aIx3f1cdtAwfdGBQ+NiSPeJkU5NNEIYE40hKyNjsGB6N
9BSwW2ISM1Pdf389krEo+AvLCd2zazG9QM9JPzn6feL9KmBK0Osj06rFUpUXYHNNFz2slJ+WRdIT
bBq09cWU6hXqsGATWuJb3UVy9/nEgaAqZBU+EVbsBnSoK2bnKjsRDQJ4KYiRbE4hEnm21hadWZ0L
TGkqYLSz+cJb+KssknPy5mX7NN8bZP4LEDmq7XelGm1Mh5T/CggYQDsz+xJoIsxmfLjnIBNj54IB
9uowYxtf2Jiu8owjabWV/NFyYBcgxpjbWiJ62o5Wpu+yFMsV83lUhllpcnEBbJvG9mEymLphKtqh
eN4Z15npwiCWjU3rrHvln7v+U0MYUbHs2PqLDRqGxWpPv97FjPVDo/cyWEbqYSL2NXRt+BFtBOrw
h+brSDSihXsYkRoAI/buSrq4VRgtQbmFkqA9bUpFAfREbKHIRg2nXMGhnYhgz/uS4jgWCtWbzQ8Q
mw+NDhMkBdesUwr3qzpyNmz/BLkPYxvkkbBC7q+tnLwazbLUcCSMF4IyrAP763D4TYrmasy93/y0
nfHHn2QLXbwPgB8XWlxBdRzzDsIbJYSjVniu5gSqRiEfXdKBiXrFQG3IMrY4dde8o72Sa+WhwxOm
jMhenZNjnpaVYPAcd4vm66b7/CNNlnRiT7Wy/Jnvyf3Aja0bPmIw70NUUK+zD60A+bp72Ul279Mw
VtumOIZQNUctxWgzyOGeuBjnWLvauVlB2MWdXsE3ONIG1Tb5IiB5vwhi++dbvfY0Qaze/IUTYKYj
OMQf2ENsp9MTh5cLRqoXR+JYBde+ImqOfm9ObLF0+DbX+ykXfXaKeGMC4IzjLnG3uYZN2cDsv+uY
lSaliC95PqQMJSHmIkdnZNYXGSyEM7BzTmFptWkHHb9KPzN27u0wO7CTY2jdnjwLkOFoyLOwxrxn
nvciqmJQMz9QTiFyRK/l7uCMUno0RdQtgUEpKM/f9ZAHdzKICZJANsgDuBmDaOTgTiZsa6z+Cpi+
vV4jeM3PtG1dsGAfGGrD8f8CnPWnJUd5K1Awoow4l9Pni2tgtwujeogEg6bfpLuqOzFbcrmSrAY2
cu6c/UCJ7ibHOz2LIhoRCb8wuGbLj179LpzZ9zT05T7P9+nPnfin4Vx9fyLpvWJMS5/3YUPWgCog
b+1RyME84lBod5mnD+dFEledPAnp96gf77Kw8P7mGo7shRPp6WzaKrsOC/V0RJJEwWU43CN1oSEm
D1IaDSLNtN+ZjJ1NVhaf1jEEeEuOcIjmdLHp1WoSLSl7kNlBscE5HF1P8+KyspTBWGInjTsYlVPu
6HBUVFt1QmpOGGuZLLsoBLEWN4lx9dfeNbhfzxctB1EREAGp6ubYbUGX5PRcLIO+O8sbp7Q5M7Li
OanqA6UnxGb6K2THbOpl/r7JaNIBEGJ6/OP2P0d091O5zjuksM16V8ZjYhStyyCuMwjc4oShFywI
lpxGiH3FeGqtrtFEwyMz6QLyzZbPGzYoAVgJ2S29AGr3JgDhT/z/YzNTjglMjtL/9hmCRVCD7inl
/hmrfMtgkPMTheKHnatKMo5iP266UjZ2ZGa+94wPeSwIdvkL/7bgfQKFQct4JAWbAYA3XQI/8UdN
1XyQ95BNNlt2KKW7lzFlf8DB9XzxSrXdewiy0PLSb4tEv0dqNHmmHuvQTtWgit8cePj01swToi1X
yODbda0mb+qfsn+ODPJl0JiRWVs/Dm10PxFUSPk6ZRXSEsSvs/vrtWp3AivNV+BidwYodZXNk/1I
2/0HXhgGqxqxESn1g2UoT6Wuu8P6JD3H8C80Q1FUQ19vGugC5BrDIf17WxQxPZL5bQ+JDX9oUY4P
p5tuL6IEC5za0dulimYHD5lnRd1sjAj1CrwD0Do/dxDCkIPlXPFkP5XXdpDwn+YIO1zkbvt2K2ks
G/X579I5+TjHJaLeI0D/Mm1QtKVwazWtSSm9uU/SAYveh80bhCV355BychWFaNWZ4aqAYceooxYF
p2q1yF5HsiQCmwHc3PvwBeI1mHoqnp6TUbqeSDAC9Ym+H5qsg1miZCZJi5UJBzjxk3rtiQ+IE8nD
280n8d34mhRjDw0HB666uRv6vrLwo3N1RHRzSUdf5rQjX/ol02Vc72URAP3ChiwkHXlVmz5xIm45
VpkvPwdbnAPT8tL7fMBDz5GxtfS/SL+zQo+FycJVY0p9LZ7J4zO2ME6ty32A2xaU4aA3FESf0SJK
qNba5vV+F9ltypObulOzH+uttZG+Ls4itEsjaQf2/VYy6439erUgW8NdY7nkgCxaEiV/WJvUa5jx
aQc+Tl8ORYoHimRQiwmKKTgn8X2iHjMc+O7Y8t21/B0OPH+7b9Z7WLeyXqtepVowgrcodZEFztYa
2UPkZRFRi9Mrv+F7qsKQlbIP1VKoepSeZmsI3Dbe15vluq/AOdTZRlCH0bUNcodIUkihRJP4m0cS
k3xQccZ4u17FMN1ryMLtN0AxP/heV+HscfC3zhJinRXbIZkmp0jprAfzevi66hpSQC4kZncTscHT
g421J1KErr6Bnv8LxZ93D/RX05vt+12HUFNEIM0+RrququAvnB9zm0DQdwQiLibTH3Q6digr+1It
XI/q4WOBbyU2qCZReCzefwKnbYLZOu8R39SdJlb+fQv986mRLGwX/n93dK2uvxMp9F0QkiV+DrXh
JGM0Nasa04PW6KfpzLkywE+wJMZI+bSH1QWQ1Y2wzGE+7ZpYi9+fsD87oeQUU4kSwgIVdc4daHBB
bhNOHZcTMkg6WjYv4Vh6DBtp/ShiS52q85VlJDH5w1xzXP6+15LQcx0Ies2KrHSsonfwHG0WQd7V
DrCy0s4rUZqK8FqQlgEyzhvUxLd3e3sV/4Fpeh/xgR0dh6N3/TmkkkUrSZz98ANnozX9c6C/ribW
LwQx2lLwuTypnKMj0KF+TY27WCewvttV8rcsOy5wEfOZKyL98Nu/1nCQa2SOtBPYSIJZx7YnkT/F
KObNq0Wqo3+DSjVXhgTs4gjfPRZQ9zT7aDvwrqJgpUNq9tvks8vxAPNCBMKOinBoLDVHfX3cWI9W
ph6NdUOPx/RUKXz3coByc0Z8/XXLvZhWV3ifZxowcFdZj9jfHm2vrxGlPo7eOMzf6mGDw2/xSGBt
efiCcP/BlzyCrD4AqHZRupLrkd2l58KL4yBJtdxi4upDrLG6VCwpzp1v5btIUZujEC1vr9b93T/O
8kejsIM4s1YklRkoqY6cwF9D7yWwAwFj0qK8VbOhxk/fJ6nKQ3/tb9MJfwlHRdmxwJseVQU1W/mj
1J+8o52DVxInbKPAqH5kiXddB4/hK4Te+rIwzUPXE7zQpKpz5p2qmoErjVfZFURHn1tduzyQuTkv
P5b6cr5pnNsvcowwpB3HjsJK8ZZsWEOh9wIs1oTadxqKLlGYsdPM3oNsvsCJepl7WeL2ntt8HEbp
6tVvf6FS+rZr/ArsdMOeiM+cakmuAZm/NVYRglg7tT6woRDtjHfmzBCfsTE72QeV1DeahCUH4KDd
mYym+Ti2gN/Xgo7BYQCp7kLAT0BBQr6safcxbDMduBXzR+lHYgPkAtQvNSYmXyVexUIa1AjBzyor
PPaekpCnjLTdtpq8GhescQyB/GDs7nkI4s1zMRJHwynkunBLIKkhPpN7L0/4Si/CIvfaJ+tdF7rC
agz7kBWWEIMYPH+vCh7VDN2XutIW9YPHQMUk6MjdrOOmpQKBC2WN3qMPplWDMcQ2oU/YcKDL+S70
ucoXYEZuuPxTKsiUPnvP3h4A4Cp9f2BoEaBGvc5fW7XAG8sFdQcDvf+/qMVI400B9Y0Ew/PkcWaY
WPjURR1lLOP+fjQmMQm6J0PxdTMPjUVRBBr+izGoJzSktOQT6Pr/uhMUmrYhfzquCLCkB50HPjQi
ch9cK5Ug3KbxX6AE173ADUgjxV4UQrdWUECs/LcOsBPKPqizV16fB+oTjJkjZzP4dB/MHmEMl4EC
0jJGMZ1wuktj3+U1jiMFyCefDai9WkVI99yEyZob7jIk+o5t4XCQEZhNRcaPMKxaal3HqAgdYiot
DbzL0pzKn38PREDxS2H4snLNRNtjpfwfP7+kmdIdtNtUPZZXgkIp/8sk6VSj0k+psvsrExmUWzP3
pplyC2e6DLMNG9LKwmeO0x6Uv1LYJF9KOge00DG99wzcgi86IUlgfrulRaSoIWDwhAYWhHYr98dP
vWZ+6gMSst20A5Y9h8XxRoNG/KTpr51y5oLcruCnAWxKbQesV+PjBjUp1Eqyd5X32e8wvgL6q+6n
Mek3F5J0sfbKKmW/VaKLPJ+L1Np50H7ST6jR4IQYOgxZy3yvNz0Kpud7UirHDAhQsqrxWw0chTWB
2soSBngyYQJwQ9zpzTnt9oEXZZEPphgChczweq2Il9EvA1fouUHEl+8RZmn1exHs1fqGoFOvMb2R
MqaEGpyr9opYUWMrsx6Q0eMncdrcE8Cyp9gElfLkDJOi9etFGmMSITrUfYD+aUWDuMlk/a9HvGG7
sxjChLPHH8k5lOEMhz7gpBDmqcVyCWUN3811fr+lSXJUpd4FbybndmnGeCEG1l5fM54x0nlqTyQY
dTbdS9rhBpXWEvxUcZ/CmzM/itiz0m4HXWOk5oW8X0qO7qh69AKOZuak1CoJWKiIYjQ1XxA55+0G
W4DuUqLl8oLNobcZESUmlHhfNkR4eyz0EUbmxXwiGhXaePoMz3TqKRIt+Wh5a5f3nOvye/64CWiu
/B/+VYRoF2g9aY/qml+zhv6ofK7oG5TIsIx35pl7US6aFjLIzMWu/juQlybTbTOmIXEyh0SRv61Z
2epLx0J3818Ny5swNjAAjMuirROubGGwzSAnHQo4QY8OP+2dbPoZiNln6p2Y04T4BXAMA/bv+4UK
UYuNaKcHOKAbs1sEsCD0bUAAAi4ybZQFr9LLSb2CAS7rthVbNP8/mw+sc5w1287FWwAjrgEvNek3
hh5z/V4ZPEdSTAdsUAPIEyvJ+Wo9iHbLWv6mw4dYBLDgC2RNU4lqH3IX/UhvsDpphdDRil709L1F
4l4pqITBNzTnlc0FDGvhx5nez83S8K2m95DPA1Y/PtqQQYyK5OS/8rqMqnYm0O32SiDh6+m3knSf
1ixRK2HuH030N4deU1yAvWNtPhVDH5Slpzf8CUXewjF+JvKoT9Pw4CzwZUaRm90bV9Vd59Lq8OSk
7+7hGeSFnPv7DcvCbaISFxfLVr5SYTYj2bo1Xh3ROU6hrd/ZHxlFUQ6j+fqfa9RV5tNbfN9UYPE3
JtPurqY9J/nEa/QLVYwVgseUrtMxzln5Z67GsRumcQYIoj2Ns3YrPP6XYNVrM/3yxzEmdXhBy+CF
mYSVH7xq3rJ6zI27gwAallqmu8J6vtqa3RrwpVqGZigqg6GXyGhtlGQdqcy/rwigyCmvgNp5cH4o
fAlGsXZRcLUZ4FlBHHmNCzZOob2QyyeKN7fDZRDYuNvpzF65T8DhtW6WU4nvD7oZZZs3hzY0VpQE
+HiBeD+Zf7YKDWT8HNCFQ/v4m5HXPQWH/97taa5JOINbP1Ugj3vJlcPG/Wh/AuTM0uvJBsFWOmZV
h5ToGtRsJceuvmzQq/5SvviPFMrXKGfdqjWNg/pvdLNM7wISpoO7t8E3CTXFbrFHYx0NXSXUcp7t
ViuPo5vkyOOWY+yHnd+AJJWVpIs5KhFhvinlkm5hEUcyewbaDZxd8R4/74YgH3i78rlVqIXie3Gj
kgD+iPhADCVyHvZzfKN+N6doiSs+UBlyCeySuU3sU/pzpCS+qv7M1SJMF04wYTE1APYvGp0xajvP
k/HlhFfmFEVjN6oSuQq77LNvHRn10udgLcdzyt8Xzpn8plsuhKgAnFB3xnpuA3GHdR7rkrSYCw37
bmX9F2CfrnBTNb66g8BPjF5nzCls6wD+fRnoEFatqrc/dpF4ms1MheBXsEidHqSFT37cwL83/mWW
HVzei4Y34dqDWYFmMzb+GRkNzyI0v2rhmwN3FVwCvnpib5sITL1+cX3vY3/kOOcWhfdpcpMDRET1
mLLwyqRFXvY3PlxwPhSxmz5MYhqMBfSmW+SDOLcgdZSxxc76l3+1TicTOVlfBdkO1hYxI+tdFEEt
byVNBh9YmRq4upiiaNeo6AoTj+fJlIITIa/SN3bFe2cnvP9dLUZynA5MurpuQAsuHL8d29wQoffv
FCBt7BM1kKK17JMyPLIXqaUMpAYObHRGEfB6E4PULAWO3BhYgMPqjN1YiYLDmyCXqqZvs7cdzXdJ
ugE0jktNS3PfhqXFGJnEc2aS99aJGx5UpsA4irHEjU0WbSTIWnGXhqn+JqeU21pc5nguosgpKksL
yFvPI5h48z1caQ2xDCN7NlHxcRZkK1Cnv/H9J82NQCFEniOXYUp4YYtsxGOfN28c9zEO7duTdzqD
gi6dDyglsJ090MZcbo1QpLASxhBxXvPVqDRo/6VukSbKuiN4p/PMZxiNcbW5Ti6dy4wl0rVO5Pwo
8pYcSvqwGgff0m3b8Ualw8Zw3BE27k6vATxCzMMcHwAqpkuhDB1fZZ/KiDHXzBbu/cBTZu7e/8im
twpdGRwf8IWnkky3oXuPrTd72L2hULjpEVp/LBJxrQ2trgiuDraeCy05b1ttEn4XWRvEEnv67CSO
nXC8MqWwhbiWfv1SPjk32/qCTvkuf2zIJkRnhP7qImhtkgjWFr+Mc4hXH3uK1MvIr/byqDTTKc9U
kx4xmXaqtk3R/COF4SykvbPW4txwOFcSj48ABJ9IrAFNHAI7Oa0sZhKo9dfA+peXeJDue62LZkYJ
gRssYqJJM6Zd11NAQZ/KKQcurE64AVHnFuu17RfdqZIUZ3n8ceCciqZpTEDaspfHxp/rZv5329dv
AaYKFJTzCzsUGC7+5Mb2YZiXox7uWZlFCUIRn51jUVUg1KYsYbQQQyFilqE456K3iKSqQGrftQNn
EBzhk/XT8KitvrljjlPyl40G8tshIHp2sFCcf+dlBGWQE/57btIx5peK09X09W3jK9z1TgcOjooY
SBJOTAzmAXhcHSopdexnF53ruO5C0by6mtZs1nf2qJp1uVU/R2p1hkDyJs7rc8rDVkNKCCRP7oWN
OMmjdcmf0/63kgatTQcAlxnZqRb7Hdd8wtH4j+okC/HGD0hEotsNZYwDUN49ElWLKsxDJYVKd9vR
icttkuRfBDKFRgtb6DaeDxnH9cqry8EZGXHjKpOVC1Xos8LHAdYKjzhf0kAyMovVB9aw92p0yBoJ
B7pJaOl6f49RoWn0Zha1bTjDKMhOznATy//v7ZrT9fZCxI7z2c5oh7IGhBde7hu1AVnr3PnUkuZv
vgGBoZmXNZ0AC0ThNHGTXT1M73T05I+nfqS2jn82dSViCitjTs1sG5EZguajf4B4TPz9zZznxjxi
uKgAssaYDrJ4gKpQ5XFWqgafYdMnRkZDDg0cqfbhTYpd+CLf12yyW5qMpwudgDhNM5x7WeyHqgf1
K/BD8+vK1KJ1zpT4xJThrEjTF2n8a3BUCbUEEuHlEvTjGym/LBuQqgNnln6OAaOj+g6WiIO+dViS
BUx5D2oGoriJ5lr5K73H+3llZ7o8SvJbRIcqe1H64MCwz/lyW8QEbWZu32NHn/rjve+cpO5C9wtf
EUJMXBAWKtiSI61ZS/2eU/FzhPXorgs8LRjxgefxGT4s0QNquAiJw7Z0dMx/nRorWPaohzfc/D+6
U5OcquDa8yoA1YOca1HtanIDHV2s/gkAELvAHUBKwY+o0rxyWHCcYD29dMhVfRy57oFoKiaxYB7K
BLnVW6E0WBEP1TOxuIzmO/8hLbfveYLnHZuHJef+3wGZyvfWu7XSct4xIUSzUWFb9dM4WhyfmFH8
sBCpXKhnw8wGiS4MB/97hbQ27/IvUWZobzPzOSIA0gNvqKgEQt+6DVKz06u6qx0HkldwPiOEd48o
wIVmfFEfPp7ISxAsM1fea11NGTDRDqYCGU/1V9DtDge3HmZ0aQqzs6VZITFxUlraQ19ZMQcuZQgv
uJH7bxld6yM7vfZrE4TibaKgCBMMgeJh1gHrJKOJGzZEbA/jTC59ry05xu7uzymKHHTFi2HnvhbC
2DeZ3ryGeA0z2pOeAcejOdJJ/ILvUNE1KUJfMN9GNHGsL4h03RXt9JH3La3HN/ENC4mfVBVfHMAK
KiyxHRDivprUe5jXD+dlrjSrkdhiwI1lJYch36l+DrKIBCtgN816r3LHtdO+qiuEl4s9IcBr2ZKq
B2yVrAG3c/zeyAezgm5LVC2cDszeu27KVgjm0Up+xrP7VgRu2mzfVpG7iq2VaWXBl/2zVx8R/2RM
BqQsZh1LTQeLk+YWwe3KVFzPI/WuzWnQCbdzK/Eb4GM4LR6Zf1wsoTjMwh0aeEY3PmmBmmN5o5yy
sX7Ho//au+wzHJaRBAXQQshqSkpvp4IcCV+5Us9URWF/EkWN8sBkILNHqIb6T5+bdZrzAfEQgTUq
TBTh7/RDsX8lMS+QBGtpM5RVqVCOFKhaO/0Fnw+LvKbbBz5m+xHN0g/FHSxCArhhe4+21YhZNhTs
kpmPSj8okSR6mJbJV6Xlp6ZFJ5jW1xXm1TIvmJJfnt2Y3p2OBvjHXfzlzSG02iPOi4URx+ZnwizG
6bKv71LKiuehN9QUclnXSK5meWpfAuBnEIZLLLrTkIvr9KP350pBvuBcIHCUDMFWB1iAfLPrnaeq
rjHkJNN/mpzpkiaRuvL5isJRNyAaltQQdoGM829MfSUcFG5HOmpg1XNGZtSQZ7L7Bjv1WCA+eTEC
JSv6lfePJiT/zKMSQ2ssoez98fMTzPkOb/PdyQyEgWv3Lhqp67Kt46MqWcF/2zTCprvPuGDuFV24
X6O+nuZdARJu7kvI99wMkxK/hRTlN/RqC75+249xoWnar1W4gxyJkWUcIVFxysw3GGaoas28tWcm
3xJ2wNos0AfEr9E7vNsXpezzC7TiGip6jujBt852SPNB30vHmFIFNzN2/biQ129HVjkn712kh3MX
9BCYMtHdHJsF8ZmrOiRKWzXK80swKc+w5PxXSnmmi69JUCdVktU8DZS/9lEXcsaDNXFL+NGRSMHe
nAg/9GI6qam/ha8oh/sH24eb1C5K3bP3RZKESrvVBhJ2O0hd8ZgK2CT2swXrir+wU7a8vYcrk4Ih
omRtd8xN+Ke9ukyOzuB1ryuxN9sQHXvcjfOpEpqn4xr/Wq0/G4uPTfCHU3iZ0BnQuQSCmBsoiGTo
vxh7QqmtmYk6u2dUP/oQ4ghCY6/+6h8cQBwrIHvGJaVKgcPcB1hqIyDyVdPkoYjANsLHUbzPbFzl
0G23npLiXRjNEyjwDpyWimd/+5X6Mh3vrAwTfmPXqd8YAhoaDgfXy34/9peD8zfrqEJuPnYx/58x
3GBcIIt6H0B2DASWIdGdJHDnmDd0eNM4by42LRU+P1cTh14SadNoUNbUtfC2V8NKAAbQ7+l+r6mZ
7zGiK05s4VZr5MSnpJKn7k4NT7osR6IIoHHmPpz4j0YuxmuFHT4jxoV/9v8CcwxFcqUXbajibmCz
TLSa4fXEr35Vmj7QgFcYopCfg46Im7WrAitZqLcX8JG86H3TEw8kj8/9s7D+tPnLmWZMy+bN6upv
nae543HvPZYwSoYX/yjE1sJ2+uiozcWeBEwF0XPTZRjiYCDqNDYe65Td20dK5N34+7B6A9evqRqg
tVEmyO9eFRNlKpxQO4f8on0OrJ0xv/h+RaWGzgeBYL8yhR5LpM0y91zPLAWTQIzYUztzGnUl9QKV
3tyPsXr5COfosg5CW4Vu/6ulJxutdJgJoyQbBETTed53+IggnE+BHbj0WcASsQeiIhlUhhzsrm2P
PONTpXS2aqNI6fbjC8ccGcS/f/gXM7kgrrDAMhudFgeeyIsu8BAEPRSrtZy8LwfHGfHqzStalKZH
m+6oMMhYxZBJZ5+wUie2GycAmjTmq/HFTw4zYp2U21QT9MOCmQ0d019kyPX3hzZB7ZhzTcBBLKsC
UpItoBfxDkWaybloqG8KRYMyGLC255lHKRV/IMPgNr96TdjelIXuhhNnXqfBZeL8QfiICs5Huqn2
59FT6TlWboCV0+jrUZfFVvMetNVdcRgOvKhvEBifiEngwb69Ryeqc7w00ZyuRTHl7Kzhh1Cun2pT
rWzzdGFuDVGu1Hm+FMPco/lLtDGlpB++pV+Vyok8OTgmiMwrwKESb6auBBSEDcWSOFltTQtdEkav
14P5YmiwIoqy+CrNQuHOH/V+I8jOD3RCx4yhhBpynoZtOgUuQq0zFbVblC73cPoqOlcNXWCajqq4
y7bt/RyuQaUwS2WpGTzsfUjgLYBqLUPGZQsHXNNl807PunXhNwYywT/tBnJvgxgZYovbWoPNZsUa
BCdGvA02Aovn8j5D34tBdRjWbqJHUk3Guf4+pK1QJ+3l0Jp170FYhu2EN/CZrJI8kKECmwQWNGGO
6+6rRAy1JKHkfcNFRZq8mCLZv4Wu3YyblnOhGt+O5N1XhH5XHhToiRzDbPQtXryxskxJwge1Fwsb
17MxXw1+pUb58mlmPSaaKeq9lsYnyLGDmBtxFd6whhmi72y0HSTEukld4q26NZzHrbOUobR6wyFN
oAdwfDLwT0t9mWQva4YeRwWdLR4HFDhFJyJfBqqBXg18KoB17APl5Dd4DQcXISFTyoVZWz2fJ+rC
85ouRw2q/xXmFrtPgGI6zZHO++Vi2F+gNKXRLNdZSWNsN1Gm/p/pVa3bf8Kp5Yyol07XptxiL6uU
Yk69joi4t45FIjArcwjbyym0t2j5azGHdOcLPlPSyFeI8VASp7TgIYxhIlZLfbMAYo11lriigZiQ
UG6IeJFkbxjedfiET+DTxOboGk0MPFsP63bBMpQypq738u71W6258Q4fHd1pHHY6RHkdV6JTNuMU
FYDb1Y123mBaH5KVdhI8Cyzzbw5IXiYFwWMjpzdRfku1uLOT/oRZNf3+Jh6JK1F2C2KkXJT6MbRc
U881KI4SI61/t1FW9kR14c40i1sguW7SoQQZqJ55WS984EXy7hEbv7FcYfy4Bx7El2wqCLYFgYLU
vBtRA8iukr+NfOPTWB2kKfhFE9IUIEeyGtxBuzACSzT85qlDDqE0v8RKbZnUDC42IplI4PvuVuOj
7PK28ENo+z+QpBqp8fqseVNfo33rfKpybvHrgC/o5S8THT3GufPn2kL8YqaCM5lQoGruoLEcFyHw
wgYvGCWdVACBm60fcgkUKzzT13FDIMLk74rFcEUWAkvLu0laEmyyyOSvovw3dPoD/Mmfr2XFbOOJ
eSYYprFHqobii/wuvMxGQ2r6XecDKjMkDkKMS1Ulj2OktV+fixwkd9Xf5rDmjjY+yfd8k8wgTr1t
JdqkfidkiZnetDe/jjKrIY9uGWfNz8lJFNL1B7by0gPrdsujJW8jgYee1830cGT2oWwPTFq7JGy7
1Uusg/7SdsVq/kMJOWKwHL1FVPMkv8UjfJI+g4FJnuQhwNpaWDD7U09EyMo5JfTSShjjmmuTI5tV
rbuz4gOcaWr0msnmKNhgmBMjp0OL5qcD1bHIJSLAFwBaT66XbQeJbk88b/365PZ92mBMFu15w6nr
o8fXMmj+47GcGPAfD/k/qKjcLpomrq8B+UwietHKGApleyvWqxydyh2U/GtjPN+w0kQPRQccHatX
8HhAldkzViclXTfWusWLY2ALAZpGUGDlP7fGtBL5pUKbw40a/ocN39dpE751Ipfqvcn/+dWZnSBR
NDKgEa2QVxmSh0mIbUlOFyH/aSIblCJPGAMqOqaAPDOoOxwCeIwsl5RJBvyQhvrV4j1zuCoxl8Y7
CNVVfkMPM6LvHkSR/DXP9pmom6GzzWSYlx203e6hIMvM8hJkKBBL2m0wV8RsNtHZaJ9aB/KitXNm
NFZQ0Hw32wsLiXqwbrW+kx49fLo9dTPkehaZt6G0PLYPAhnWO/PJlQtLcyjdHvqsf4GzzIcLM229
86WJeCuKp6CfA5jdPiQyqF8o7p8ffjPrcoZk6ska1rECyFM+YhWwbzb0W7uYz3zpTb1A+0JPhyIc
+6VlhoWACt8j7agYrl1NCM3gC2ebK9i3wugrq+Ay7AXb7sEWSGbMUYHlBizR6GCKLHTyfDoG2kqg
Hz16vIfZe3FlV+y/M76fVNHlK26yY3Wm+o2x1/0/yd2/B0aEc+u2YXUifEyJ4ROsmWy8Z9njqnHA
62ImdI7+o7g4EEwRSk+k/YyYJMreeABtHKPV1uvojcmFRc2VQo/B48Sh4fBa4O6cTfZZgY4kkoZ0
6ckF6Ju2nx7xxcQ4SjZpAhtboBRyW4c6G8dyqv4xWoryXyJhIdqgefBAAYdcdhmGiYBSldbxlPPt
DKfkB7j/0FH6YkKxyvm7c2cXfJ5NDNYX2CTJ9nGVjXWcgKnYF8+hGRbET6JK2B+NY7PXPqP6DYmn
Ovs+vu8O29w54VkTkdyaKucTuZqu4ryszTvRKAXzlRopwR4IAIasnA6FylabRyNeHkk2jbSwJ52g
jM90bSBhQFYYTtGfzLmjYm4ynEPO+W8qZKCcYJ2tlUUmVJoPueBhv5vny6A6ZuVK7qGLdvIQCoE1
xqyOUnWWL2aNQTmK2dPu0Pf1IeTQh0homaMW2CWEGNbUMMCQLYRdydwxFYMy+JNyc/CRPT7lSZ4u
zl52/10oRUJVRhXTCEjFllgJg1xVTVQYFE1dhCHnfZLSDafCTnf0PUpAxEgaZ59jYu00ns4wq0LQ
afyZzch81AaSPylE+gwBUvt/sYsvkI3E3GbohR+JyNP0XnD8iKlS4fkYad1mVgyH+sJhHes+tJpa
58n/YuCWL0lHTlqbpGYiEXWEH3GbwiJk3ZIzqtQPkk+qKU1V90BvUKZBexsHAUcFr8mfEUCMuWhr
QBSdsZny10z8fxjIvT2tcmesSx5JtcKRWMFHi74aAozFrYyGIo721faT/pTq4SFmN8/hAOK2839Y
Ccbj8ODGzY6uWmS2mi6WsV+tFN+nNbOt4GYNm6e6aoyWRljFugw4C/E5mNfJJQLxXkQptx0XfAdd
xCkVvBd1npmNINc1bDCM3I0e3B5NFpDJQ8YAo4nkGViILC4VzRHvmQspJE0v7KwaM23mLwaxLNAe
OaQQRbDdO0znGl44X53GO4Q/U0qOnsNo8wy4LdOFfXy/mW8MMkPF0mSrLhPGQhdhfN2nPJsnD3f3
SkS3lvC0xkodlX8o0U8w9xRzKX5wjTTAL8AzrUuyl2i91T8nr3iJf1fZ0S/3ERNnJ5ywKCzX1Ddj
joDqV3FN0BvT2PIDjXg54JU2gj7E6B7yIhcqT5Cc47f7rEpL0H1unph/XGmKDoiaqN54wTwxaiYa
BHXq8PYpobzeR1M9hmioyP6/6+8qa557iRWFB+yqqAeyBip5N+YAWFPnM9jcKPHqBvzOeaOXO8R4
lffsLcAP0QtvZ1po/x/7fLXM6qFyecshO74lenq8f6wMA6VXyPRnbzDHz1tt7lkO/0qp1DZOFC1B
aj9lmcJqFe9MP1ccdmwMLAyQFt5W7WldoPfkDZzIVuJ6+S/AYMFWr7EbsPQXTZSie+rG1NdDyl89
r06doe4ts4lWZzg0ooMgNapMkAywMM1CKwgyy0+IfUjfbylEbc5RfbNaD1nCl2cYHWSbc7/oGDVL
QRMtjY2kM4OGrRz5YfLW/xcSl5pLQAO/VlfnnEPafbv4SGR18zJoTCeEVh1z0h3NH7EsNtENf6vU
0JTqUEkrC8G55Dn3hyydgh0xni7JtL9WudlMJSrfqxqmIpHYx6alsuZiJI4PyCzmUL7d96/qB5PQ
o3PuLygUzyum2CxIOMC0zrjiKbbDScqDAeL4oC5e+jXxtoqFPbWIWv2nqnqqjHtm1GHpVjoDYbH7
V6wQL4OhsZA73mb0qREwmOPQPPINXtNz5iLQmAs/njqWFr5a2MRf42V6eewPgJLCS+0iXOlck2N7
Oz8gmHRO0YssiYAISC6x4muppJY3K55C569mOQ7m0uYRgWP5cAilCyyhay3VFaY5nFu3uHje0qmh
uHxnyUjfuEJbxbe2DxvF694tlzJgVBlBglN3KHmnwCJy4C+flZbEtQdZ8NrvOGZ76u32hluU1bf/
oWdjhOmubSeEXveDMd/nDNA94Y43uExLBYR6TvL2WnnQBLHyy9fwqyZ/rH9J1zx+4Fm9Lfgn3lWw
QTAh+/nL4K8pp96emi1i1SBOBCH/MDVWzwACvE7E0gY46vrzbXGS2kxkTB2Lc6ezVK6ttfQcjpZD
YDE+DUxlHhW8hh3yYqhCSwn7gEIcSP0P8bmL14KK/KQCRJtShRPR6tG8yT9LT+fTZoS7+vKuQ02t
ySXPGSOcVChL8qvzFpKBSxgChFxzsLGdGYwLKaY1TM+sgTsLUj3BWYmb2cs0ZJqHb/8P8K38dRSY
BtkJblr/lWUTRJBI2y0elSgAPKLI0iZgLEZ+mnA9w7RG+iL4C/pbv2t7fsnwMGqvi+DallKGlShI
jwlSLKNluliixZ8jeYWW2mo9pDFCC6h+o6UTE7rMdhM0eC2O1dtED29X6oafGcfTFbpkuo1aUXA7
NFJWbKDMg+vPGDzsnbwSLP672KI9u5UiLG8auhK57uqaPKGDOMcXpIhwqcXWpyw2XAGdTXM82fnZ
EKR/AW1ptV+zvlSAsaxkn0Oc6Lmfu+eWsXT7kcjKLaFB5M0dWqKzQHc2iosvslsNR/lnoDH4pamK
3dOTtcnbJ0EaWBFXXENbcPwMjfPNjT1baPDJs7yV8gE8Pw5jCjn1hL+C809o2NvK90+AF1loyZzS
45IZCdrDxh6wEk8iE4xMUQbyg52igfwZXiZCv4bYD3hMBXZMc/AJXM5rv60Y2KBK4Eo9w5EVTmR0
XVlHQBPSqDMFi88s8eUCoN6RttubCDrwWjgLAJREDcoSV1yMbhr9xp9C8Xzo7ML3WIVCm6+37cIR
lf6B+Q2TqixCo92hTyUXUUHYh98RBJ4qALVBtoLRiYEbUrZON+Ucwm8WKhF2DcvPIPFhCOgCU5Ok
C0MQjwhTAH4YMZg6L/Jkz82+zwQbfm0SANKJEO0hqPBRhU4omVFxof/6vSGuk7MmXy5LDhhwysh7
3AF2JPl/Oj1vTxVk3IhvOBi+Qq/XmKukA/gCnfIYW4dsgR4ED7VcSV8xETve8juJxznAylWOdou7
ndoA+wazB/j9NJu4BmBYuBdrCn9YISsTi3tcjAg9Qs/jEeTujQdigInbm9NFbvoREc5QBckbk77F
KbWbVy9OZ9F9yTZXqtY97XAYAZ9lfXZ24MsKNJjfYZuVdZMbS3nCpEnlNlPWwD8rdpk/btsjh2Xa
drm+eWY4v+aRZPD9gyzGMgUkn/hkPfTMP97zDoi95cGbV6KcFuOiTeeaUn4HqUm17im9d6uXWgQc
iWrdKI/irRZUNgUu+/H51ON9Klfz88jH4+kbfWqfzOlELdYMEDbOjSdc5HbfLlkZY8F0NN6G6jDg
zkRqgQr9MXwlEgwaGsToEHz6jSRkxKOQw0BRkTQjIKQX4NZ//bOsCcPX28xyx3/P+UEGFHSQ2qWt
IQ2yd/27xwbfPA5d9K7YWqxeQE4Q+/PUP17KBOB2CPdxzUPXitu6thasx9zKMQj0twryVjk0d2RR
NKaD8Z4WHjt5OCfoQhlgES5Ou7uVwULfTwNYjvUreS5dysR4QcMMblm4HL4dFGOunBTEPZxeiR4O
FQB+uZxAsHyDnLatp5+Kd739xmddcXVc/74MdaAk/h78aka+kQWWgX9MR//SCXjOtrb7Tw/V3E2Y
OLH4t2iC2A2K+8QXen01xYKQLEm777c9PfStugdYBNF/lbkGaKkG/ePiZ4Z8pnJCYrte2zXaZecL
/CXYCREJTTk6MHDEOy/3RtLBp6Djqi+lnSFOpnvH9pyg/8VwSdwOMTA5wIQrSu0Dm6nmz9yrbcw2
Xdi+21jTw0pgGv5/wvy97L3kD6i3IUq7IRiREDzVxaatlfurAvYzmDncOGGt6smLepbRgLtqC2UC
lJEVMjHRZ/i1HU2wog18e+nbWl7x8aC1aLTHc4XV/+fuc/GFKxjizaJL/Z7gy2Gvw87Ueh3LlQqT
bmutwnkC+xdgwXmid5mqi7XrmTusok+iSTXPVWiLbtOvgp7BE8C6kjtoL+Skzwb2urzb6PygPtq3
v3SuWu9Hb64iqqonWUmFZ11d4gGD5OLCybgrmBxBeyTRkIists2M1+JTtX9UODN5zhX98zEPGZxx
16N9kL3l2RxIy4zkU242/4WFmHkBV1NC1OpEipKCXXU1OQySwKEmifktXsNr6Yt0Klpf6y3gDWyx
8YBmCjEr0wfTA0AICqjg05ldmj2jvd1sQMhuc6YnineRi3M57WQf9voCB4/Tm/uBvmrgBfrXCrl8
dRpaDUZYARyTKGgqxUtWoYwiOHznkAs3Q5ChfUVQF8BWex/P0KYBPr+R2nyTKQ/Kf7lco5iX+jlO
MJsR/yajTsuaPxCiBlyeI/GdHmRMZgW9n1DtcCTQrqgM23dR9jN54UKchjJS97T2NVpw8JOWw/3h
m0hUlpeUWK0GedqtD3tffd6Zw/RBXirbQStQN+zXDYNwlwbrSOCSXIH/aU5gnEkuuvlRf8Z6GGxq
0VOJLJ+t0TGTpNFtrob2LUf0mqPyGxlJxbBbAyzjH7YS5Bf7xBcqUQIUe1CG/nIZILZQhaaNeJ4h
LEOjUdkE14qb8egEuhVQfpK6394dGTE9G31KUZ2x6y5Xt8BSP7boVMlwi1NwhH66Bd6Lnn3xJEdp
JpHlqQYQMg71bSSNitXHwg4HGWuxfVoTNNpwKkHWPGovKIycY6sAngLcWZ6U9Z5bzBhDCNVoW3k3
h1P3egrEsyyC1URceLOZZgA5VmmtEKtTYhgfd1g24wrGPw3+2BpdoakoVLIVyW7yymwfyX1aeZnd
3d7zAmmFpXuiAPCH3TWMdlKCFNrS7ZU1O54oqnD6RFc8U7SeDqIXeCoEZaCcG0ac85BwzLz9b0nt
gibf1kp31YTq1tc+WMFTn0rE21k59pAE0EreNswvw0+oGYoaudKz/ao7UDHiEkILr5aIhwffBBNx
z9C95peXCNscTdxvm4gf+7FZ+C8IvHnq2ICqMyqfIbWNoQtZVq4R5c7IDs4R5llRfIz4ENdKdeCN
po785y2Q7eaNzSQWg44ri1ocbyUAe5vivF3vbRx309WflLm5TbsojytBt5uQVjz4m4AnPb2e5Mks
GF/VNiUinRGcn84wP0FOQgdKhypiSJSBmjcSyWODpz9hqMfdc83Zf0ixmcruf45LgYH8onG4s96I
tPqLAJDjFwABS0Xejq954+cfaLW2qkSEAq6up13/dzrPuX1ifQoM9uunkGLwzmetrrUwKhyUkMws
gf1EF1sZKmSmZjsx+EArWMrs2r2kqd0PLUh+/vSMcy6strhq2NtjbJVyQNRSU7VwngsriMimrnmF
HdfoloB69/X4b9FTvzbsihEcZ13WTjyqv+GVBE9aEntfLi8AMz0PphkYzWj0b1bozDnqPN0ekVFk
req+tNrpulXSo1q8eDbJ0P1pgLmlh2JHxuuR2M34AMYpxudbrAoJlzbi5KfA/Ha89W6pAC3ZDvxI
EAh9RBXJrx8t3zkSQ9xk5z+VYv6/hARSPaU4LzW/fUhYbveXJ4No6zziEFDFmSmg7xRnQw0iuDPA
GHqQVgAeKvPfuE4HOelKa0Ccwi1PyzvmzL9LCIoFucpAV6u5Un1GiIVnN6FZDgR0TcvfXE1Y6hB8
eP7aRbgKgkWTemKHrd1f4tcWV8xFLO1g4036Pe3qOmuB5/5glDVb+awJTM5IpqxeyQYurS1rH0VW
3CHFT4sBV29Ypwsy2Q07LulJwmg7K5uEroKyr0ppoSY8KsjG6/TFvbIGJ6Fju7+CYAX8KlUkXv0A
pmNsIZrPpmQAqFtvighnd15r+ioKEenNgUoIr8sApFtO6zAtNoEw9MDsKG3Qu0GpqszWM8RWewB3
igsmRnda+aZaAzl3pWVSvRRRcPFhd2BrRbLo4SoXGPKdeBMkIMkRyemCj4ypT3vuVTKi6ciu3bHq
bsVeE1645Q//UaR3xyP1uDCR2ABDadJ0Z1BkR31/vxzRUR4n1Lq7q7/cpDAHwdnPvLu7gql9ZXfD
94JRnJbQfUjU/yOrILSpm0d7BVwxi6N2QulEIYE8sjKIbfIPocsGQGN9ce/hvCYy+VHiJC5dz++7
Vlcg/bYildivILCCQhId31DT7URpJRAq6yMpqmE12ZVVGHYEWCYxgv20hA/cX/geD/8/lT1Jw4F4
xrAT35Lcl/b8mQWUlnNQ+pWQWOK+qkvzUmtQDf6dNaoOC7z6FYoRL+EhPGcSyqaxkP6WzA+UddZH
Lz7GNIXziIVLhuGfm6Mnwr3Nr1pV0MR2BcapN0RF0tVQUfGVShOIpKl51veNlpT9CwjXlZxvYOV7
a9B9x2/hhIeL5r83SB1tKT8tv/bhobg2AlSyzBqL2b/Xh6By7gd4aVjPInZNAi8DqDSOhhvcgfix
qULByw71C/OWCXaAEqKeRWT886qDcuUGK3Ncf9WBJkr1KbN8CUFvrJ7BaqNH6c6hyMI1jakbYhxe
w419GbSZ4Tfy5SrsYosrxK/jK6TCixAqTYlWYdHzvvgaZUGv43THGK9nCvn6zSlupIsslkujJOr/
HGuRqzh/amHdDsyBv61eXVacoSNRSu8UYh4rHmfrAsUh6noitNwbe0s4CB5SArntNuC0SoxaqXb4
5YpcrWRVF2QLdgwU8TxxpkVfyKJMXxmRXiBn7l4VI0A+2hBDuWmz2OAzNc0xELcRp10dSdWrr4xD
Wqq/JirZ6u7SuD5SKw+rFxLrjZIDGboD7GjerchO7q+ndwa6ZYAXLQsxQOUWk8pIIRKEwck1Qv0v
6XB+kQUPqi7lqAqsTXYv7J1Jppv81Id5RPQy5cRWk+YW4SvQl4G5pTuQtNE3tlCSWQb2pC0R5WE/
aHluBwzvwamETzBc3of4grxMIJASQGncytC+ii2K9slf5x0KZVWTN9PCs2tlNQW6AxolguSkPLAE
yjqOqJTE8tEQY6aLRXfgcoEMhc7O87D28KegCZ7HjMTcO4VZ5lWkL6TkxM9wiy4Xo6oKmi37zuWQ
na0QmWZqdxO2Y6H3e4W6TDViAjONDHcfyUP9834b3uenDDt5IaiS8TZwz/XqbqDZ3CWTjbBkhkM/
P3jhKOVq3Bww94otwZ0FdoYaqDBmWADPc6VnXUJjL75NGfNaMIOYzm010vR85aFxjKEdd4iM96fB
pjTS/WNB5A/b+lnhHILNIx+/RKG+cAueDH8bYXMjRwc6Tqh0ZAQ3tTGY88+FZX3P1UqoAuLXeABs
pNcGAe02wLsHdB6AFW3qAyEJNtEL+4iIFYwYajPelRgKkOJfRGtEcCllqHtUvkWMLOug7R0QGM2r
Hh9mUbjfG5OICY/Sdu8HU/Do5QyP6lEeSWxsjPyw6Vridv//OWjbCPsq4C+EvaWB3exMOZIC+Zqc
X3Z89lA/Zzsao7TjpVFJa9dbrHFcK65gdiGz4bW+7zvrIfFIfU5JBz80nzwgUdmrKn8zoRjGe93C
ccyP4Tv4BbMkgm2WE5cci1oELxSxno/sQ7Tuul7DI6d61yXIcILKmwqShiizEJP1uqFCc2cGnH0x
6fBoiA6PV076ZOkjdB/H3o6ud4kM8Vm5ksfVjAsFB3S4ztTiJYhgQZiQajYsxhPja4+NlRAZcsBb
ZbGtqiClNyYR4fE1DZ4AGxbAAppIFWrbUDq5v0UyAR6VNWEDV1nm8d9AmfHGzeJmFGWDNd3WRDgu
gRtpp6KYQgVgYLetcqaoGuFyl5/KtDzW6XZyupJQ28+ijjr+GxbfYh89KcB7CUhor+KQznPDoGhy
77y4StK3yqoRV2zUIrkwXdFaqOcbgdR8V8O9Zjneq7LyHZTtfOMuXQHl/Od76fZI2ASFsh5QPq88
6yu5sXRIV25jU/N6s5cAKbUsVOOba7kcmZIhMrk4jd83LHkY/EFtVaXe2gGUwxjk/VjcocTCWlTl
9E/NtCKGqxZjdWNJHQm/bohkKDs5PCGZr2I3yBXGeLNiEUVdMwfXRSUlE/qCxiuLlS1Og2AiTXhg
8fKUQai0wbQQAb5mxXCeBnDFDV0NS0HZdPZzkfKvj5BCconH4UT0RCkOSvUf0usqEn7N0LYCENRM
qnKXDBlXXQBc8+bSaLQ7cnehtzty6lJLxpV0tGmO0DxEF8Ka0jfbytr0QEvCzbIBjfxd2gcLzA1d
HAbwpgo41LmsLoEJFxu4AyIquGG9v08HtDY8fJonrMcdy310dbPV6MtqV/IKshciQiYy4iUBwCXc
zTXEdljJR5gwtswtwj4QbJKwTNvEag3FxBXwbiNsUROsj2pEEJeyxpNRmYQNIf/b8fixnAlllCMc
PDn1g1zd4wiyLEnYvzVURKBMkbMKoclM2fzpOClHi85SAca19Bp+N62a8yeq+BiKOa4HSqCPg+Or
gPnUE2PkF+OpMiIT9YGczvDGmHibR4T/wZ+Q3z6/OSqRPmLGKwcMj0vVhOF5TwL+uN19U70gzO1X
j7WTELSKuoNGUH+wL+zuUtbBdAMf4Ffo4vAF9da0xm2Xo/6WMArXmR1wORXFLI3wZMTuFtrrNvmT
Pv9y+VK7cCnq5z1+KFuD719FahgqTuINYJBzvEMmuyGfgWNRLlDgsmVz9FimBltSHF+xOuUkOPKT
IebYMmuprBWuc6U1HUtkyJXxHPEvZ4epbmk6Aqlx13ObXm/Fvd29tC9vCYd//WsUzX4pAOzu7Yvq
FzagPsQWvAGMYiYiaiKZMx2HzSMmvRb4nlfyhfsoZoH2tJXYJDTTix0WutWKoiCXFGGh1nrbmNaJ
/3mlL3N0yp76ehL9hLd/jBX8js283xw0ZFMv+/MCn/MpsIsuG+UtV6EnMr/7Ou16IgEjCOEiDKzy
EQbGdxGSlzN6Vjn1KJgQDBmBKCE1EL1apxBPuYFhPaJ8XvJ2Pc+dQe7EGjphJgBSjwl4TkH8MVpa
lAKTJKfQkCVpuF3NbJeVM7cU061eCwZfzZZp+P3x5pP8ZaTdmfI1hw2NtKwsCcozAVOup2M75QKr
qzw4sdIZK6UeA1RmA7cx5f80ZV3Flcc+Z1jeKB/AIDZ6ovQlwhqojP5KYXvX5/jjiHNBKr/F5ai/
YNXvs3F7cBZAqdqpIY+nQwXTORMyHkHWAT27RCd3JTJszWgDlcNdAEoDgNtnaUjZa6Vp4J797WZz
FOB71ExxHamyCMtS0QRCF66Ym4THbjHFWi5bhtjeILHv80BqUZ4B1C0Nlr6J3A8jcCs7O01lYsb3
/Xwt8QgKezwMsYLg7ZsviwLvodsgcqatcigIkaPZY+/2/gkYuTwcGj0lCswTIDgYqN31QO5LU3jT
IGf/m0xdJApK/snRX3EX1z0sSFcDmq0h/gt1B8YHZaicAWOCPjthySet8iud194iqmAxwvtLHApN
ULTY8MGxy3KV7ckCUumQJ9ZFe3ys2uSl6tSNFe48doXSlI3Sa7mGsrNxQc3CVFesrSd4S6XE5Vvy
eJKiJ/XatKkeN8tJfbbwK16XRMvHMLGkODEfQ72U6iSPV5hxkPN1kNTjU+fPMmksHk+5UTgMqlQN
/g1okSbJXfYWbjYyheSraDSZiSYob2qfmxzafsEaVt3Ec6lyaTqsybmTVUZfadwRNqhZla7GR5ly
nB89V0conFutXQEu8PF6Row0PBW+RiazKUGcmgFLvm/ptItE+q4RHiJYsJCV9YGBi1J592GY7JpF
i+Z2yz+3SjnVaktBxeO5d47iyG9OgpqoKkhUqztGHoIF/g2Zzrm5JJ+/Uye3u9CZUCoHv2b5qC4h
FLdFct4xpYcGtTPus/9qdp6H3PevBAMVhZU//1l19gl2FdiD7AYBKYvkphXbjMC2XdzDG8qykiZl
1cxW44EhanizjJ8BaWXtyTOhwQSpTzgVMntHdLMYheoSZw3pWyF43mC0U8ksYrcpR2bwEuJ210Er
URd9ZdgStpG7sKQBQAEQgVmnfNJQ73bRG6CopKZcS/AcUr5kyHkszgtVWdxUDOYwU54wYCtEScUj
YucCoiUXVK4ACQ9SD4LwGlSDvidZkVBT733MwvKz9MEy5hjbHcsfPE8QoBDYOCXNQmHbQqRWtm7d
bbzqnYqY1arKEOwK8qw18QacxfTy3mv2ZlaD1dgi5apJjTHJSDfPExmR+2MD9uRPYoCzg9yOyIcN
od8twbyY1F4u5xxQswvwPIPcb5+QTbcCBcxafdjoOSrk5IHScCKbLeINVJzOBbrkEyIq6S0oFGN3
leb6mYlbJDowfTKf3oA1fPELWB0Cm8d2eLiRJKPxuxfFqiL9inSI4ruWrJQSq6e0x/u/eo1cGrm4
oa4+xfg6pDagwMheV+/dtXDlLkVRSuOEngT5TFyYwiVR7VryJqB+fwUbVIJzWp9Y7LuSHLC2UZEq
2iPZClyJ5DcOkGvJGgRCdCXm6hWNVAEGYqm6hyDAhjBfFE8NhKZAHQNY9ztHNG47MilYqiHfLFup
mC5xROMHeuElZuTHw/Ib796MbYakkNnwDQy5Gs2erBwm6ncZoMXQ+uyDIUlbj46dsBdB8e/zyUWJ
5NdLLZJq7zuEno0ZA+CldqfrZ+WdAkjVTy0KnEvVYilBG7uOGrOi6OxE4Bw4BCwWY7vUpguwfdef
iJbFSYOGUpaYy0EJdAtRBGyU06EqOCuVKo4UtM6tZEGNfz7LVmAlb+WkEz/ImQyNdWM1O4mxAiBQ
nsFErzx3mVW3nd146+p8EPIZwzQRD510PxtFTzN/bbl4XJz81sQApSxUGSHnKR5hOdPXhE7RzvZV
BROYeiZubxHJDwEujKLFsF77Xh5u1SYTgFsTMurWKiZiJ6Vbnz1u4s2Fnpvfm+mWfhJ4kSDW8z1T
6yPYn1Jujf2Yd1iXMXUgkF7hkxDWkpViNoxe/oE0G+oCsASQnwiGpkRr8NjFaKBv1R+iqiepZHQj
XaRlLRqnfeOkRPsHr1J3TUbCymYhC3bFmcfHx5nDAqS2FXsNEebIBgUpA89UI6t8SxHN0B6F1wSD
aRp3rEqXgvTWHA3PbGchrsbZ7gxi6AKeY5S6zo0fELCR7UMuMRTnzCmxcZiz2y2YaFvgmUSPsjQW
ixvEa5kh4swd4TOCU5T3OcEzdOxpdNCOb7EPVRZbJVeLflzbV1O6JH8HgBQA2H5KSZXcfwWScYp2
jI6fzQjVnvh3kxgSg/szg56djkUlSYUKZ5pTpRHNzMNjR7IBzK1/BdH+Vss9/B5QhlAtnkEuKAMS
baXNZATybkC/0LUocFsNn9U3nkJZonnQQ1vKLx01EIuLMqbOMcEnToNFdhToJYJ5kpdpBPMRHe0+
NUk+Pl42ITtL20LQDXwMLBgPaw7nViOzuy5hLBetGDGYojy8OhXLI2C/yzq06DOdAwDouOlbrUmI
ValP4faDtCvdeSBXlZxuftNgDJWW+pqaX+jZZLp95yXCoQsOFvHVuEomo8nDdOd/QffdLbsQdM0m
tS1KkfqpmHJW7aVGvnI8FDKhNoif3oiUlnVkoyy6mEsdZ3xojzWwSoptJOqn8XAsytj6kyn/b9AN
smWHZGoTxi1gK4wCCnGfWYiEHgqZZE5JB1f5lqU/2wZpA6X7/FF/e0hIjMvZ6S64lu1ddVZ0LDCt
BZPirklWJL6BwM1MIC59e0B7TL13skoZPzzB1x1jUGe3L9hBJVEIgKI2skWcCigqJ0WH8ief8TkK
u8jpFxZP9vcNWEiqwrHjSOqi+VEDSFC9utQ1FKhmppbRamFQF7dzd37eTJLoYF8UF+jCLvASchcx
XPfQT3qzjhpXyr8Ve5czuv61Qs/kDweDIaEPKZBIo0X0VPD6rsgkJJH9jFp5lFar9cjKx/xEWkix
he2jbWmGb3NfU1vpyRQ6NfnU6bsojDPpBJKzkIk5z8VGHNZaJ7Kva8WFtxSBC6iMTjtH4NTeagZV
bFuc5NmYofqcbboTEDrRFEQXjJ2NVc8pJe0MNkLHFMSOZUg4f2Su7obmR8touA3B+TcK3xtQxHGA
GQFJdYcCwXTbZ3zcmU22C7HftO4AFXb0kglK/k4SHt8z/MQyK4FR/YTC1iOrqUVDmqZPLlvJ6ikf
CFlu3CgH7Mtck2hNm0D6IFFiRHYsRdXKd6XbpUB78kE/uwG8Eb33DQzsZtWyq0tmfAOR2TBrgTox
II0AJWYPcdz/FQbmGQ6EiB2xZHVqXjNsMEjrpQnbW28FCrrYrKAAZCYGD5PzflQXVxfkTP0vy0zE
wjC5+G41+okXpTfbfpmQ13uhMU7DQhQp0deyKOVL5CD0EHoFOG/TJPcj3R6Z5gpYqjV1fUJu3a9T
anlkAo93XPom3ZsvTRj5kfGuN76IvHhHLElcYcdzf2cv5QOx34Fpl+Gqg7oAFYHtOD/mgH82x1Ky
jPy0f/SMBcnlR1EeACrB3r58J/ZlVXCUrG7Vjgal702FTMijh9Pna9bh8hquQuAhb553in5SghYF
c8iR0uxPrY9q9YAU2wJDgQ9im1w7yiQz5txPCMQgS2FOmxy1Q/x15RnnzdREyUVr6+YPAHuU4qVy
xFn83nf0I/0ANNwgi/PckW77pFueEmTuMdf9+utl7znsAEQAAxPDBaYXhCJ0aQRLrkjFOiZT17rB
ckZjoBhK7ZIpd1kLaQDuyHNbG7lJrdYmFulin8TCLOLD3L430U9x8ZZgHu8TQxMVPb/NEzBZ7OPT
dsdEDGcjxrCcyua87/7/xL9C2/0ZBZY2gYKJAEhSW7CpLFL1brNhhvPctU7U7KmB70bP1HOh+OCj
erSny+2hkz4bK9tBJmR8OdhsJKqW8ybrJg0KFJt67THiZ8B0Z8b3NilIZrPZSoN+kOPCN5pxoJyw
f3TBQmBNkA7xcgpQvhvXvntk2ejVksB70d82vJV3Mg3v5ynCkjr6IWZ+IMKUgoBkeMuzqtRLr6dR
i1j7G+kJHuW5jbbTqjG2xkPjCq4TbjAgvt2VyLjCLuyv1tyEr01YBxP39FWJRHXr61AlTLs8S11H
xzUb0nJOfIeYg8f15p8TM4meIKZbnLmbBofjs9iXeIXhNCCOTEu6L/szw7EzWZIhibiz0eKJHynJ
h/gqpTqe2dsYWugwBQIvH3ZLihfn6AM4poY6qDkHjzzgxO+swYiOKyd8yhhEscUF4wZCp4J4Dxav
IW0bgjzXz2kvpTu5aC8354C1mghsr8Xzoj/vRUcSmDEG2MI8Suf4GVFco6e3Ji8hpQHKq2pvCUR6
YlkZIgVqp6gR2bfzPeLcL5AWQV2pq6Vi7CktOQa7Kdglk4akQEuii3Yiwi+/htwQtmPsCJE4q5SH
ObSN7T33R8j+SbxgwkeQe9EzzOWB4ICIBbpx/Afu2ea7M5R3xBblE+JE9pExkF4BKvrks8P7Qe1W
yXvkiRA/sGsjTuvLpKqoyo3L6l6TenJt5k6L/49cq7l8a6y65Ils+82aT6/j9cX9hEJmCeDk1mvd
b8FYAQXOXO5zXgDjvrcX1Sn37qaC845hUKN/W+Inj0OTMWVjLCCT2MnU0y0d08VOfiAjCUd94FxJ
zvTYRBiQhC/iQLM2mU2Y2GRo6FZtBPlpKI8CaUQxTcjnMkgPSIkMVWl8vQW/afSe/wHYHIFZfH3C
O5iQZ6onwTAhA7sWL0KFS23zCwxrVMFwPyFeupq0WhAVv0aARHLAvXCXUQNfGxEc1HAr0CUNCDtn
bY7PJo3+MFUZYyDcQ9MBld4SzkVJqNUE1zaHtVJlU4kDPyOiva6GUKVb4b6vGgTVrClIdlNe74cO
u0aug2e7G/74GrynkzB0SHpcciUEc3EthrN+J319//G64PK1EqnE3415ZvKloYyUJBlJccxsvx12
K1TxnV/MvJ0tF8bSs5OsTIsyNu2PUAfe5BWyz+26DPxTdVT/Gp/Ofi/AtA/4jYjAOwaXhhRInr9t
49qOvDLmvPCAfA4Ob0fQqbdsgg/UnWAXhUwThE3VNXRIcD1Unm9ZDc5ueUKyGk9g1zrx/xgU3Ejj
Z3mzUiAKwdbgaswlCwUEu2HdbLlku1vSh0hfviS8FknkpQNyNiWkiv0ZMwTmoYDY1vnR4kvZvn8C
3kwrxsqJX2+o1HSq7JE0xxWcZjkxgZRpQ1bnIUBSaCaMZbRhA9VQd7UOQYOzLobYebR/kmlFPKrM
stGGgzJlXfD6SKRkaEwGAWGukUcuH8XToYa3eSJMI7LcK/PDvInWcbOhKMim08kwn+P0Ca0HvRgM
T90b+0CZJrrZkfqC85RSd/WgxpgX7csvNXiAmPl6ewicj2b1ocUMzrutJG7SufTMztOrLHburSzS
yRvvuerQNQpemsNc55g58QRMYrlzBLLmp5w42U0YW1HdMi3fz9QyhUDNUzHxESaode1lyCm2WhR6
Xf8vk/c94bxyZDy/JzLqTg+51srQKWUbOq4jOx3Ny6G79bNwoCH+x1V1rpSswyoN4Rf0WNt7FRpv
D+660/8pUJRuusZgT8VmOt70X4cfS01nY/PCqc30j4n+tkYE35TX7xEE4ZFFjJL11kItGlJTUMnu
0Ze9cAfknsu+gMeJclbms2sebzmkujGjg/mui2FHji1EVpiguCT7nrVAr0j/awHYtPu51m56Myw2
St2GpXjn6EDupII35mP8JnwkU9OOY0il8bZrkjSYbmIi9Ct8fcZpfAiw9kuok++oEo/jt2hzqmxJ
WdC5aPAYp/wmZ3HjWkM1Mzr3k3yFp+nmoOcz4hkeSgk0/bW1JTn7VI5vD94zHayX8IP9JoIKxSIN
UBraXWdNnQHMPvXd7ry76p7guODJjBnIq//FV12LEBDYtehzvnJQ5274kebGTgFPgVWhzidHimtT
BxIZgMLUWAMctZYgR0ApdhsU6P8s3YcSH6S2hDxnKmo2LRkifP9I2YJgkEPIthIhVYZdiF8pYEeL
OLbuSW3xm/T30RLXbrby7rb8ZGXGsOiIZRSWiTHfRKEGZGoHFSLqZoEYYX7NOD/YBwtCC6KQVo7p
9s5fIwk8X50n9xb4xnQOFUEBiLUgNzXWTbe5HCFx2rIeYKho1BOP+TAC3/Bm4G5S4hnFkarhJ+2g
0WrPOZtOFBY4Db1SkqKlwPXrA+VUDncLoawxIoK7AQFJjszdNtrQyASARCd/LScofRWFOZ8HnVM5
OKxXRle8IJJ59KYfiw079n+DAQO4AwW4NsqU7KW1OVRkdRInEFFV3fVh0yQXkQdKZIFH4zMw8Euj
kVnxnSQTj79suVWbW1GN7YAoUERuJRYTKgzRUc8hEJmJCjfaAKQeqQtHn/jiHArKOH9cErcEVrWk
4PMDe8JfnZ3JA0xj+HpcEpoYMyOww+YLMKdJRE/YWgICriCHx9r8Vam2+bjDZ6viODueYhZ3vP/W
8EzMjD0vokuzb+VUCM2faFpOnOqxFIi9Cegsa8ohs3+CGoSojb6S2EEMeBi9a1YA9gL1Lz39bHCO
x5mVnmRZjlpEU3q+9Zom/hy7KaoiRvB/R0elPiq6FygpWSDTWdUNdfJn8bi6Xtp3HR19eHgZI5sE
PJbTQldiDc8RWqspr0UHppGYjGHsRPVh2vnCCfFMWAQmTT1pkWVYHFRMsFajpGzwhaodCKQe/Tdb
XpNiYrbd1rq1JYrzV67c0vu/NHuhGq6xul0stGXyWwArkXjkcjd12gS5WCILcWLqHE6HY50X+Ddx
LIb91h/hAvgw36ew9zyYjh6HMliANevVBUoi/F11lzESTxOuJS3HSlzg5ZBwjOgi32lslYNdgLPO
KVA6oJoe8O82uMusL4QWG0VUCQDabF9U84WYOufU0EpwxO1+EY4UD7j2if5fTgKbIwyy8rkf73dP
KG99xazrym9YmqdjrB/95CGL3kRdD+6ZWS++WurGJITtoOGXyLrUFKgsdBA8kLI9tqsPeBban8gt
FpNi/rnJjkFddLFiEAUeCK71vVqPocwr+pQ6utdvxfM3Xx+af8N/PVEgrkeQjf/pTvmrEwks/vvY
yDjiqcoqySrBATNUYr+acmKmfwt/3aij92jLeZskH7/Tv1OY/oz+Sr0dCFDJSgDMx57hAc84ypcE
s/ft559sMfBxkRhWWdxZFmu3j3flJAfF/RxRulGrzMG7h99hclERgUHFsV9slxDhkSU9FCu8N+S4
rjr2GEbDqohN+Z4+osCBFckp2VGXpZ/rQp56h3JCgAbi4D4XBZtt6uZ2jpBjXMEuOc4/0jnw9I1x
6UqxVDbZrEKTccH/M2nLMXxYJeRS1pJiFsdnGQmbJiXGio504d1n7YjUaPy4dCKqTZ2J+lUqryo0
IKxV2Qy5TE1Sm0s+2BxvkeYzz0PS5glCIsw3ZJ1Imx1iBHrvTIImECGHMQVjA+2BXcp1wbQ9rdZK
iFjbSUIRk2bNkyda5EpebUO+HFgVtpVaM7GWCQgvjoLAF/kLWswKM6evx0wcxeCD8wZoWT2GfR/b
Z9rtyTxpz+7GLGdNfC2/QRXR2ehuv8faykqVivS9T/10YgKvirpTeIlJyCYBRSDeV+paZO208Yph
sVm9E/d3GgMcFkKeH6k8QduH7cmB4iMc3XRUJykcM0z0/ZRfy57LIMtAnC6GJvKc0r74X6vVrRru
IuJTDP0BKqM4y9JRmnDn2QqbuN5eqnWcHFROuWc+rM5IF9gW/BkXu+zqZ4sPGgND+fQ6Lh0qF7fM
p6Mzd8BgtormDcewNXFu1rLk4D93YSvZsyjDHyP6y5clww2bsQ+jkI6G10opODJaAgUWHLThY9Gf
eOkcnbBZRyDzgF4XFrLN39Af2Dk7LZPuyyFH8SiC3k5GlL9Dw0EtTtL3Qij2DUnJzI8DW3z0dWxW
pL35Do4k9suwKAP/OJ3tMUfrqC92qBmnN0RXMOelyD11kKOwsqZBInSMKBKdlWpfp/47oY9yku0v
l88sxXjw56QOYWLmYe1Y0hAKC//9PC2f+iYBujq+vMtDPYX3fSKf2NEsZHMtT07JBWm7F+nMUOjf
MwakmCGmoQAYpAVUFtX87z+NqU+BOIXVbW6TjIZi6uX8L5F8CizM/h0VOrt9m5S8smxfSjCh3xQ9
dH3vWvR6abdnWkLUbE3SWUcblr3uccIRCdSvYOC57BY8CPJYZ/GlhMQ0y4m6ZzUrAliI5BWEusfl
0znPUDkYhzK+f7Gug5icE4kvkcfO9v8IkF54XTacxbAgu+9YBJcAAzE6KRf+e8B6IN8gJb4OxKm3
kCVvrskEeqd3h7glI5IbXoD1mbsNOf/vfWxDqkV1kD9MaArbpxCEmwXCmqE2qlw2OHpL8J6Xmyvl
cx0sRyJBxl9WK6/Xq/lNc/W9m/KszSw47+P/24J6d86j3iXc3E714G8nVLj5hlc6ts1QxnmyYB6X
fJLW5/sDusvqKK4bn3bcvHAGUUuUQjdrrsNA4l7WRTRl8Q5S0Ro/CxtMXIeJKiaULFJ+vqJIqsiG
kRL4u3OrQZNd7ZtLaMB+k8hOlPZxDCFBSjHB5Lf0VBAn3E52iu3Een6DDhyx08Wot3wtkSgkTVDd
u/fkxAEhhyfDMZfzfdX4aoX1+Ebl3/TxCoqUJE3VOd9FXceZQnFHk8xKBKFj/9z5AdmwdZ06nsLY
9jiVZxfNAOS+sVPIsU5HIhw+NQfGk+KX2oVS0lbNl5Ka4wkLK9rHU56+P5SbZRnXQm/+HOkHrpOs
uKMcYLLmQAiNksI9D0yaxiMXM/0hRw2PhuIBZSZ4zsuerc3IbAvjlLxjfvzaPbPQ2om5YNWBC1ZN
krU8QEBrW8w4Vl9Qb9mwvXhs4x2MwSKKzTHU7MoppA1YTbxCY9GKtRNa2HNFL6orqWjWaBmmCZwq
4iRUuf3ZZX319QMaMt2PKOlO6ucuA9spZsYjLJU7T+G4E5UJGjlhAzi9hZXbHBIqxpDWNkx/h9K1
4qtqqbM6WguLPFiDp58BbqMh/D7EMDjNCc0M26HjjgI+yZLOwwz5gdwziJLggCpOctinpoAf6/F1
64qf+eAVuYc37NYiCx/HO3g/4rKFL/5gSbqmcbhYtjIbaEOzrnSeuUqKdrbjbRlpYLpYs+qXh50V
cBhbCC9xml8sIE0GvA8a8uy/V3sg69ese9F/PL5GiAfCxBzI+/LYS6ERf2xTtwZIrbAr7mxURius
UrZex/FFgpfeefYIqzVwqkdSsY6OtI7ADuLQct36NnUIKE8/iYWFPGkVI7xG9RW4VqV4H3EHRxnt
xHrGn9PVePSkCzyT22VgkkBrzYCZW1l9k0mfPflePUUnKaJ3qnZCaNJDc0r2QhrhLYfKF9YLIjDc
Q6fhaiVuA3otjGZi+V1oT+6uAyzIP9B/sgLtvcJIdza7Eo4ZSbIk8x2Js39iK/0FI22k9dxCuS8H
ugTgRotJXhw9c0ZaJU0dWtZFI/UtB48588iQpem62j10AIWw4V0PLvDLCmZfyIIFABVTZi1mnSIB
e9wpOmACvYEM+1gH1uzRMD3ZY/2em7LUo5f3fXlEhzVjgU6b40++VIbyJREMrD9/ANDgQm5GRlLq
iMZZXsOfP6QK0k3xN8YzujZa6tbnRl23RXIrnBYeAxdbbSoUglEGLem+WsCwqKeR+ZBDpv1Sp+F+
NnGuwGeEqI3DZ65NNiOKVVQqtr6+8tPpYttTl4XcA7eN23pHA3SJlfFTSfkSG7prQUMTdMJGum8U
7gm02UBcFFX8RynCWfy2Cx987dPOVLDRgDqLInwtce0bWMawzQpoHXshj74T3Zu8yTkrOD+VZs20
QVOdeuv0rp7ey6A4jBGOKJC3R0kMB1u1O1EaCVDmsElroHksTUN7kgoV9giolCZpKoUjIJoIllTV
8ilZzEI2NoepMYt8jjWhaoKGKUlaCfTBajFwozkYPM03+Os+aRAT6xt6sjsQxpwPzNteHjZVnPOe
UQUoDP+hoDVO9Tlj2f3nPDh6deU1KR2j1BdGMxnXgmPTdMrDq8pDEID4NfDjVL9OjrI+IqCKk4oy
phPNZE3rUVTahZAI58r1OwoJclfkx3UK8AmKMmTSOdHP8vLmR53fi5s29TRKpzM6TeWYdJbcChoJ
ciSxw1VKG1flgxCdEt7lXBDj32emZmU7rwsmCnKr4cIs7y3vmG/Sjn2hET7MYQdtexMWpRcx+Enl
7fUVcqTPf6OY5mayleSvUdpdX2irou/xxv8IT/P79Sen+lo50KCtoQGAgUe6AS0awPvFYmyx3PAQ
1pW7K+NNlUXq4hiQlQuZN9Omg8mrYfzcBvXJwV5m0Zf0Q4q+vMQZ4bwMRpXGlGILql3HSe44tJff
Y3XXpk2L1XQ1pZyAvmDZ788UlnzyORoiQsLmzmkdUrkqOyPi9sZQYxhELSTPZpVUZQX4ncsgTeny
ZQKzwTJYAKr3ANUUVEe903xHYsdCjBtGXe1bUPw2SUXa3WVg+shvaech1PSYFCV7r1ZAeAM8zcuO
uiCyT0j2CFNwNsap2g245AnIN+Wv64U6p0oMqOUxv43AsURlii+GyVnaOkfnOs1/4VzNG0PwA1mH
Tue33HSPu4WEa0gprwGslNs6ghxvDptVrZoYInZhKR75UzC5/HABqH9gDARE5ZLe+gVQZ5uiB2nr
EtSxDnAtsohn0PhJON/QVgHEkZDWKtimXV77O8Ovq2aMRBheFo6y2tPflhlH3Wlp2RgKfJiqzNl/
RrYzKDu2fbAlZHNonkhFKJ6YTtlnFIz9df3G4Vnsmk2AnDuS4n3Mv6WmjeUh+hQ3WuQiRU9q9tfX
sN/zWofbBpFLDCUtX7f6jxWsJLMIt9umGCv6Owy6AEaR/Msr9uU4fJ1x1nne21kVALM2PT+RyMU9
2mLJnysLtk0tdICghuzVz4cj1w1MsvNNoIbxc8ond4QuPzyxCNd2Zo2OAs/QvCJQZrv+xmjXDxt5
dN8rTz8SxXirGb0+hH+gzqsl4hW1Lj8VeuBXfDGO2xLFJ0dSpQJengSu+dIrl67MeQ2ObdKg860E
djZV8fciXydRCVM8WvVvbwda5gvM9mYC0BFRCxKEHiKVmn/H5XI/Qin/nTOAzZWMWULJ/AwzYisa
SeA0EVU2IxxGNpjb3MoFREn3xwAOvJlJdw+xAMMlUIJF1Y47Xm6s6VpY+HhKwAmqqInPf24jqjBy
tp9Vh4lzwoQs/4yH4lMxdkm7bHYnM//Od4UerdA2DpZYQDjxqviYyeOBKg4p+eHSw30Ih2qnJTVN
OrpsM33vGMLFTguZz0jsm6LSKAHEczCrhS2cP99IEu0uQcadwLvvQm5t5Uiv+XVRW19hAA/8oAor
irnmVR5WS5nSwUi79TU10sAwn99+kzP5MxdKVHLZ7qerjM5c+1peGjYuE+n6FvC4YbylujltHtFr
vGYCFkYfQYOBISmuLeKm/JcYdb/6A9/YkF+JNVgClgCNLwCsRZ9O5H5uhp7rkN/9ADNUgfCi7M/k
8iBiiHG8awJjTxfWxKLRyYvGotczX8skmyA4JJel2PmsbemhNGyCKwenWK218uyMW4M5htjUzFB3
wu7bxFuOiGzTVh81iXNPICTQhdr2Yg41ORe6dGJrlIuxHIX10hMg1opAVpTxvvNMrAcUOziZpcoC
LEkZqVs/29d9N2lssKg27tHoGYTf4/fpJ4VbTHNJAlDuDhgE1Mrdz84jzQARdrKtGeM+8dpt3vLj
2UK458b0t0T5vsO/ebEHSKd2/YPSzCR466+XPzGUwNB1C/CPC5FtnoUWDWp5O+Z0yv/pBfUCM7Ep
maXip7xncC7UvTeTe64Sj4eZuoO4u1F4TmWxRsKmaHQaGBBjlF81GCzUZoAtCTkB8bRU6dULhepj
UOk8Uj/0bmlHMb46VA1WFBG5GbnPiFJW+ZIM+WEYGqgW3OzjSnXELWoOxOMnFWwL55QtiBbWQm7X
BNiKwBW5tRvZ6XI+zxoNOO5d1hX/faU4sKBGWlvxP0mHIe4SL1iyEs/Ry+CFkEABhifif8nnVEiA
eTHPP3SCNuYgnXrWPNHVT1C5+YNVrDe9K/g9GtiEZaDy1OYZ8SqTpb6DUWiPq/BgAGwRDyBdDzJk
tbG5fGmghjIoK/kwUmcDHoO63suUZYXAtZKgumjyiAQjybxFMKnPX7cUxMQhYv+7raiyuPhyqENo
nvlCkMLN7zs6amm6KnuFp5W8lKrJGCLO5nZxqQnBFpKr+6+cyBMP9pmDLZeEo1Mun3+2Z/QrxuxM
wBGxZj8nrd0gkwymvuyhX/GyCtRRnoei9H3vHlhHyWig0t08PEVqK7T6pAfxk2sxejl2HwLPpJnj
gl7OmW7caCKJ1zF5YP+sI2eiTAxWdXkbrBuy+NCRkpmXTUh8rTvQXPg8QG1X1URRvza/ekHjDVPk
rjOHxvlo8Cy2ajPY4qRjeJFD8Thux/LucNKWzT7IFYddN9oNdiEea6KOYXagvuBwFjB57enlP3nq
wjRXx9+SeCrm+sF0Lgw6p7Imr4546gIdxSOjGPfQonDiw/Gi9F7Jr7lvJRf5eY6eJBekFhCHZ7aT
7qSO/PclIQjECNDQfVV57kKvwHWtjH+NPz5MlYQ7cJqGFXaqHIqjS0M6KuVtolgtCLM7QH82Dw5I
37ndFkeUDI5qX+h3qxTcVbugsL8nZ/3AWuCGZQWf5iIqEJRpPQjlk+pKv0sMoqA+H++zsotpNi2K
ObVB2oTIVujYRxFgKZW1QcrHUnKDSR9pRk78Dkm0/kbv/qWEXSb5JdR/mPxvoRCbuuXfW7KEa3ZW
EZkxK9oC0eBrFLF/wD7E6uI6XPDr2a83Rg5rJOrz9m5rVlB/VdfeLU+R9jlbxkE07uHdcwd7D/sh
2mV8873lxkIOnG/boXX5/2urBr4uE/P2gDxlJ4w8c9C1VfpMGYj4fGQaz388ee07mFpKYriyiQ4Y
He0LDuXhPndCiomfALH1WXcSXLO/ljt7+OH3Wp4Os2hgvWSUzt/E6xovPM63SLWxPQ79fLfIAFsV
VoYD/VQdBr7OshWGcKWN16KTd+eIC+J5R2QcU1qjKcBmTjngxLSiROa76Feolz46GmwTghg/qSa5
sgzvQM4s+1B6xFU2B+7jq+UZWsWD07j4v2sw4w675PPDo0fBOneOqpphB8AkTdgmhYv9F1ZtatY5
MzWsrVCHBSQTujIhiv7WdwAqX5ZP2WGvqrkkRWcWS0QEzKasxaF1Ev2++ntsz2K8rtWsbgo+4VLs
qVWeZh6yNulhmfDKsTCKjcDRNlQsHwvL4wbkLtuDuNoSu7LgqVWmIsEMX+a4zMZksRFrSjZh6YRQ
l56FeXeXHYXK9zbVlIZ+f8Tn4PjWUYktsmdeuZjexJ3lMfXukaykgSrKMJWvTvXT5pJC9J6fVFiY
4Ho/tAK01uXE1S6xsywOhg7G4t5A9AMhlmfieEChX00vgWDyaSnn/6/M9iwW93FerCZZVGHY9aK8
sJz+Ha7yox1+mDAtkViD821/ViAY/cqxqiR9P/5yXbM6OyAFFInLllgHgwyG2xp/sArFpemCDh/A
Nk/69OhHiHUg60f8SdQqzrxCWwn313jDmNeaTYPlSkJC0DFFC3KfYd2aGqzHXBBUBYY5/eqaDRHe
5HmAK/unK0liwvstdixuETAdqtzJ9boIHqQU6iF5dXKH1JS3cGZGaZd9zLtTyUFuSZYjUCqsQP6o
fDMm77bnKYcNiVZM0Jtgdy+lDntJ4e8+PKx8E4JbaDDYeCIe/h7HSf6noT71TVa34m572F/7Fonc
aBvrc+xnfL7Zzl7yLqw1VKSHXKQltiBqrmS5R6g8ZwPRS3gBT5/FLtIqrDVEgaVvJYySXtKc0kx+
Q0IJ7xD9ky9Dh8/t3XbkDz8dC1Yt324i/h/z7Hc090NzaA31Th2bYoc25zRiybLxsCavZHQ3yhYl
KSR2apg4gReS1VUar1BIC0O6FMsN1rGbFifWdTwb4WPx4APmyxa7luXPoXd7xuki0yy4VQOCxQ6L
3j57uK6zVX5JacbaUv0+o2w81OaVSpWdI9yhIDuu//+tTHRvvFKzmSNzABvZa6Aw6ro6Doq+0E1n
xnnhOVApArga4BcZXZYQFltSSSrNgGANQzfFrzCtqDJz8cCF6FNkk4K55QjgSn9GhrXs7yUrwL7W
CEhSHT+ACXqcZh3KQY/jb1N3GSNrdI182hTe9GJVNg6DDF18gsqoRjbumR7Y8v+RPlJONopurImW
e3V5pDfXPuL0S3F/KawktiGPkD8YTT2ILQM9WVZYACM152CX8bR1EsvjP12SeneuX9QTU+UJJYfA
b7v6w7cTLUBWlPOspxJAWXLoy0Fzb7j7Sdn77e3CoNyOHjEy/fJ0qC25wXX0W4iM+eXTqHGQ6cKA
koj5kbPhQfwx+0XK43qr827t+ualx98oNERu3kIw+oEIpgefFwFDngPatXzrofHFS2OCCboWqvUT
eI6YpfcyNEPC2nyjooP9RjoCCHxKFgOAPW1Ah04iQIUr7GjLCbIALRmY0ZGMB2oU+c9WVN6A3Bbj
/YpV97R3//GyfuUv1V7Pv4PcKLkQG9f6R4iRGTZlPexF1I29l+mbna8L6L7lNCKPgD72T2782xyC
IRb2LdzgTTI/9QO8tqVu7Q8Ydcu0xnNjaDm2fMOp5S2lxRMZxkREw7EtVLZjs72vALxN54LRu82q
rEghUqHKrjUR0aqDTqOAKasGJuorAcsqHBNEPn9aml/pQ2jTHIJnMLh9DNydJGO+xBUHU+xP3Rah
4z5Kz7lj6FC4YFSTY0MTpFRtOm1G7hMyUicJej+K8sB6KxQPboRJoghcEwmzKr7TawEHCL+1Yura
E7QnLbNdsENxbesarfULO2UayqiU9Gb5sEt2cRLctu6ndcdIWuk1X4mcBw1fs2AUWXlC0n1kDftK
AP7WP42hxfF8ZRwJv7rcla5/mdn07ACGO3WqvcESAhwtqv9TfpB/VUGFyFxds0WeOWBm/wc3Zmtg
4iOWqwq5jM9P0dckPUCKJoNrzz9SUfFKssh5eVMoKnOyKFHdlFFueUyBHCHWN0Vxl77HAW5wFMr3
IDrKK9TfO+3rm4e2ccPBiMTxDlBK4YetFLSr69P9JTUPcozpLV5xwAi0hummqgRh9Un5Z1Uhb2ty
mwyMImyVJbx9l7JrMCJrgKER+LC8Z+1mgLwIfR1ArjstbGudut7PKKuUbiT07xQ6+jffmYwrEmp/
ev8aIuNrWjv1H4N5RZiTAoo+KSOSPAEjQN96OaYIguO4tIuikMPnBi7UOGLZ33ZU7OOuQEw+k9JQ
/NFxku2PM8TgceYbo+Kejx3RQcR/6CNMdiGFd/DlPTqS1bms4Hj0l0N4i51Zz6wUgamnZZSKwof/
uocOn02QX9Ip09L5DksWcM7to56WHbO0TxHOhpjaFUW46EtoxoPXR0gXCFN+xgUhIxDVfAG67wao
FYmcLaZA0JPKxG6OengKrpBJjIslFKMEeboH5gohaLeEOjgJXMqevDIAip6HvOUfNEc3GzjXPka3
/tAIvkHTGJykQa562vstmAzyJW8YtEjIErSWan2ecZM+KS6yfJKp5lwUlmnsOSsam4Mfvse0ZFel
SKfXIkaN2PaydAjdMzOnQbwlwMkriuagw7UGZuvFPBbUMCf+Bq5ozsdIfQN/HGnpzDMDfokoLBby
/iDas7laHsEcyu5IFsWb36puBpjM43ZOPIYpJxKsx1g/DXVs+lB6ar7bLDH9mKKHOX2b6OfthK+U
BRFvcaAtHGoyfbqIFNwbU9c37iCsZhnwx0NnreUIgfBuVo1VHomprL24r4vaW4wAYr71+UVhI+Sf
MvB8DVoo6uM6EUVSI3nGu2EuDfaSl0lb37uqqEhPMBfryYdKwX0EB/dTdCSzM0hyo97TLh6eZlSc
szusxR2EJDPGgrmq4bMXvcZASlkxd+dYhROG67tRrcBTZJjjFWNMJ+ksKWw4zcwd2epQNQxF96d0
k1XsKt+82+0/t77b+X7Ad0fA11KOSgDJCWdX1khLGFoEP2tnqOykEFJ6Ifv9UaH7AXEMI4MwIypG
bjDttNqnNGfl8QIC+WdibXVjUfkD6C2Cra6wW0Gl8sp+EvdviAUXZl1NmFsAuGBTbOLPvbbFy6ha
ReZAr8/O4vIJctP0Rxz05rwsYT8Ggx+EoOCpTeruOeQGyGEyf26YaWQXr6yl8qdeVSa4IO/MMe2d
zl+RTqYt7AGlHZYSTwO8Xsr0E6YA4AtRiut1eZMca5fl0cmRYrqpJsN3f9cYBxhTqYgW90AbStfL
EEUThwKbhMolu4xNrP79uRKW3HIerkVGzetMsG7PZfayS7DwMsJoLgtxX11C3jmPJdaDYAVaBOEe
25skTgGuDPSFO73Z84LEmAj2OZPoatqpEfY/vRoDgvNh9+ms57K6ciURQDb3MzExPHK30/PSyFge
hm7pcr0sMdAJWzToRDtAc6mftiNFkmAsyVej1ALC9staUTNudxL5L+qQN4oIQzO+uU29yEQqBWGs
Q7q1q5UqJhf4KcCpVLBkMdq6QgkwiY/5aSqhL56ChBuNCUbOeVDpQ9q5YOx7uAyk4me92+mPkhmr
iMJOBDTHQjqCTfHhsEdR7OjKM5zMiW3GHZffiyjuVm06deScQ20LZMd5ofwFMV8yOg6QY8dcibSn
aRKzTaeA/ocXuNcjrn0TvvtcjyUejW26UzQM+HvQLvPnLWOYtuneJmICD2Z32jgO0ygDhuWlqSd5
x17X23WMIx3t26qonDo5B6rtCTaUP4bYdTe5mRpFgSeU8qoeKpYltOXHaoulq6P/FzYhpizRHHBP
3MC6hMLsRSU3FoZd9Hw/LXZW6geld3DgOu6+0ryehV7kFUNX+xnPR3R1FvvPieiY+LZkBdwjaUDf
0bz+rHyBRgAMSDfGF+10XEMOnRmjoo8IcPWEHKHOBQ5aHtED4gEZHNU10hfw531H6ZJ4h5BxCIto
749uMHjb6S4H91BSZcUGe4TJG+r2MPGk+w5t9CF+IuNTND+jA2mjnvJPdy1Gpp1q+4UA920YTLWc
/cifG8zdHzHi2mD9qkt7+N5JU9l3hvgbeGNIzA1ZNW4aXNXKleFthbssmKiylDWZgN/MndFrpkR6
3TkqixH0/p+nsXpUTIvMDSseCaUodfx1boA+A1WevwDbgJcvTj7G9WuiGehtgZuzKsQZzGJunWUS
pEGaMvyiAQSl2Wi1aN40EE18xbrgsGp+U4zMXg619t45ze46PRqRxVUMFjTbuqz/dKoTVRt9nKsy
juXCzfKi4BPGwNsZj8Tx1SOxetUtg1nupBrWi+2o8PScwXgL/5fg7qbDNWzRPJuY0jJ40u8b4oPZ
oSbRVJfVOUIu5+rMtpucIfSntuR74H9MR+RVxir5R11Edb3aOBoLETnPUOZWS68ALlmPP9GijFu8
DIciXiBQjXznA2JAXkiFki6C6Cc2rnp11hU2YeSLqqZvuznMTlzc7wDaEOLZP+QdA4b/26Vb2a35
2AsGhkZZvHDmwT8RQ+Kkedu9I84ktXM31tfm7pXRidrojJiPaxemETWsk84w9eNW44L7bvmLDnmu
B8mHdYQAAU4eGwsECwW9EBza0xGt1D3kevoQUsUDh3OpqYsDxadZW0Zxfs5834iQwg/D3DqRrKQJ
fk/+4SzORVuqYc1lKZeoOmCyT5Rab1wGnZ8VM//Mxo+F7liHL95q8L+xqCOnR4ZMS05oAT/0VYhC
om1bwbcuIJWK5/uvtcEvaOxt9MOPrd99kJ4YLImuAKj8yApi6aPhXExohe4i1d8WGbe8HzTiZCjZ
1c4zieH1JI3XA6RJAAcz31CKGYwXUrzeuzEI3UJkJrlYuHbfcBztiI4hwdDL7pLWfgyLqqJGWLZk
J0PNp9gjKUwgfsji7UZjPgLSVQv8lajd72NihVoFggpi0XfO2Ut3jItZt0bgXK5dPVBavu/JpK4l
IV2nuYGLme+kLf4rNtVvN7vPBzRLUciTq+FoNCkSokWMzDynNPIJ0Pama6qExIaP8BzQuw/Aig63
pGh1O+0I2EkuvKo40IOnsrgIUAVJNKH60/I9DFV4e1J4KBNLZ/O/cg9KkBGzscJOIPBtZNvzWRex
a3jcGvP9fBHt4fAn9dqURUGnM04bJlEBxOOw+43YDg/F9UuTDlABPunq1BD6s1gLliiaGG5GTiVN
eV/oXVocjGyNHdwQkIay3N4RhvbIkkF3jHD+MbZtx1+OJ7xbFgBCNiZ8EWAo3d8bmK6vpACZG6gm
r0zfTqoNyMLt3uMxipRkJpycdW7CjHXriBtj5fAx1G3fuJoulzBlPcyFqWtUcQlo7VztlxuZwGq3
Ed/ihr8xcfj0ctL4GmHbSgdZSObGYmHqnP7FPANnTtxQwTM/FzkP9MweJl7kvxNJwjJmCc26575x
RDhV3lytCJdL7IymcPXZuOy37g1it9s8WCEgMA4axpSKutmOwhJ/DO0xwSI6WyASJpV7LSXgxhKv
iyd1Yez00QKEOoxG2A0aMmN+gixYZJIhQ6zrOjw28+Kn0MbVDDw3tncxO5BPnlKHwNOB/3I96HR7
cGygHHj5JdWulfRc72qiRcnWFiHHfUal7HA+btcb9Mda53XK5lflmB6/3vyZsQ00W2ExKGEKRP92
LyrmoZAsCZvkL9me2N3/v8o5vQL/On6UKugrCM080fTXHX5qDKI5QhKYq655C/pAKDzzJ+CsusON
nsEqJDxPqGF5sAibQ/fBTxBhl0CTX34QqKAlP0WgT3G/EYxgHGH25RwPDRRtVy1/UL0Z6z4SCsti
QssfuOBueZk7Uy+qvMeD1qDCigvxp/se1Fw5ulJSdhIbodWuYVFjhLQzzpQLDP0/gE/R9pQSze7o
Gx/DKeFsbeYGBzhb+qAkFi0zzrUk8Z1mEIaguY0w8gbeLCi0pbV1oruyMN3E7sBdkzZ2ZNFeXV9g
DMbRqdVzkCcGBu4CZdiKB+wp671+gP7ZJ2x00VV1kndnJnYf+4Li8Yd+C9rggySxE2FIqsWrj3EK
jIznqdSTZzxEFsXcC2rZ2stP/9X1H1xemEfopFPjY+yRDMW1jJzVNwxQ+Ht7i8rtv2Dt3LguRWR3
6OysRu3OC5N335oVLn2ah1QdbLns4q94CCgE6sXY9SNiF3cCpoie588kVuK2ve6+gtcFXxdhqgdE
EqdJaN/+NWZEB15mN8aZw9v08mH7gUBY38pnWCX+ITAQGIGzF9prNQlm9IGNlXLqF8KOqgnwwh3Y
sbuyc4IPRJfmmvvWc8vsMF08rVGjXRRTCxfmlWVWMObDqAdXNnHQbjFKmHD45MYFAMwMJSXVWKA2
ARYmOkMYwtS51AOSYIZtdOKGVr++DD+wtS0wPUef3lo8iVuBWPLDN9UW7tZD9uxtSVhrITJdc/cM
z6V96NoDlME/NDrebVYACQNGJhUewRDl4eLakMqNKyaPWq6KDRQQq+gRp0LjXj51R+cT5cOTs2UI
8w6bXKwUmT3Tpd+NZdzwD1fzYJeijHTNANaQGj/Vp99N7UNeF1jr636bwrUXWiPQx01AaiOTSruG
q8Y9odKKcrI5KVhF1pLjanylQWQEvL47+x1NJTUXQu5VfqogLehxR4OGd3BKBSX9hMRX5sC5qYT6
kgPewCAK7lpAT3cwda3gIE4OsMt+aYHK5CMSA5ic9iXgKcgoHglaDEVVTX4vIDWXZim+HnfhWOnZ
OAoH19W2EVIHqu+P255ttGmmnOWpE4pUx3LErnfMOmx5zhlbT3r0MKEYJOmvZWgpcu6PLU4j3/zY
buHw/BWh578/rTuxgA/p6czfe3lY4MA0H6OmYxPbb8FehgDIPw9iuXwhkA9Gr28w+Yu7kfIl1xnN
QXq4EuMPhUT3+HpN/HBKgBd0m0PuweoQbPwLy/Ugf7fqoyzS7kNJzaVwkLcfn9KVFBxEAoLEAnvE
Is7ta7MhwUwbYP1q3nSvun/mev9C7QYcxY2NOfdcsedFJIWYFT5fvkEgyFqBkEtwWoLF1aA96uxr
imJOtvkfX9Cqs2+NOfhs/KB7lTkq2i8EwRez7e7/N+2ukIiNjCQpEe7oVZ0rX5vhUwlJZemG3o8J
1NOkv3nlAmbD/aesatv+FEad9M37DC/FVTt/MlzLwxIdIl8CQEPdDriOWH7QMA5VlvH9txPyIxti
fZpKbgCx6q6d1QX/CQQNe/Ctlywjhu4NxuV4UzBpY97CckThrr1U0jSl8MneRSk41qATHH1f4zGO
1qMWLnYqJ7CpnSzx3CKBobhaqWhf+zzybK45heS/woj/t7C/W/jEvu0xviYHoINsfKpdDyMa+2ol
Xy+ChYOxE3u+ojLr5NyvGGn0Kdv6acsbvFvm8GOEGFXbWNi2dPEd0wDhhXetclaiV9uzDS7u1zT9
ct4suwrz0wa1/z6L9G7FuHwqOBZNDPHMbK8SsswBNd35QjA1egmbro27wkdlXPaUq4MnfWuK7XcV
H1WsjNIPSPiW1e3LwbUgEjDRjxVQUdNbNpQkNomjEYjFKM+CA0bP6gRVNAsevqU1ooub2kMAJ3sI
5j1K00u8UTYpd9erKk5EPDVR25izdTo90MicrrS1OZMZZr6GkPe/kMzcD0NFLdejfUgeK8YbMXiO
fc9rA2sBKk0NvAVL2ca5XVSwVjToBnMVqSMiN+J3AHl1EkEY3Wg1XVZycPmAU3NqzKdFMrFdNKJX
b8eiOjBHg40WwWXgGFN63gUvB3a23nJJXhU9lm5EcjmGV87J3CpZ0YZh9vv/x1Bi9cbtFvIpzglG
/VsbyyebtWHMnNqr8tnQn2muO1NQjwzRduB9EB5EZOuLEoQqkSl34jJe/JDIPYu0UqFpu+MLdRMN
18Z0fH69lJnAA2R2hJ8BJybCcAeWtg6Fbsud2Lel2I0yTqlA+0MrYmQ7LK/OBYjSbDC1wy68729m
2i6bn630Qxp35SG4KjTQrR9BWfi+dYVXWSUVfeSaDeT+oCeW3auX+rqs9KCp4UkmeOes9xDv5rbc
exV1gc8e19jqDrUWAX4khaduy57e+FV4a7aKmg/SB1M+eAb1zhBYozYcK+5kbcbpC7w33xKPY7fz
XGhnbqo6dFUgvHNUrSSXYt9gjhWVmktRMZDbULP3YKVmBklRdJg5qzpWHUNiJo2fqwzEx/vE0qHc
QTOHIK8+Ur/YDvGNtDMCRUgwbqWcoGbH5ZwGqrqYsXP6ruZQ+zxu90FqFiMEmFXGlLmRASSQEgyG
WCvgnlKZsxtOF+rR6a8vjOtgiaGKyklO1QpEBAcSAbAjodXAxt8jLiehm4pHHvW0yvmtl5gj/lSK
0LT1HA6gatOyyPqn3JDEE51kHcanyh7zrTWQKbqjQGhp5sc/YkL0Fj42ll+YSY7XbUNH4dd+YYjq
gUeCRfV2p0tnxLuFJqack2dafTag7lMdYHFigxXC9BpziqIWWvH2zHqocpLlqYM4XTcZlZnGDmX4
qpkA84dl0M2KSmFxY0238qVmE8QmAsW7ZP9wTt93smuBFcl1W3BZnnPWxqxtJIfuRU+5aWguUYJn
gMVu+wch5m/p2peAm+hAA+kwoYiTwApua9rLYZyaW5cCs4YOl7peDY3luZvM3QiUp49jK9gkOYR/
QN/m/wWmfQXgM6Xun8FbtVl0Jt3zrswJsje5M2HfbEdRUCYAODYxasQYRM0Aii5IgzErthcdG1NI
yeNT/t4cpC80shvpCxdyFZU/vq9EMiQp6YL1ZtNk5Qd/ZmqJfBUieJJhraLJMJiJublULe52Na38
DrRErSNYLQPc4ThxbzDNzMJUTEfjFtNSxOto0fz6de841D1FAiyKuDz5dgnRgxWWxtekuAEQiR9r
KNmiuWyT8jRz15L9Y6Ad/xrL07CclHiWd+p0pCTzs8+JiUomgtZD3uLGrxnU5VH7XlAfRpFSLWAG
mC2CCzJPbVIV5YErj2gEQeKsNmA9AJopueA7v9JNQrq0eduYNv2PTRHkSR/869dia3sJWckQIAUk
0NSKLsl3T6iw9zBlDOnfYITF77Hjynd0Xg+eiWyXa8AGVmbM09MQwKrw+dg817XNSscfaib5fUFC
/wtnnDgqOuXC8ShJFfPB5WEqKCjQQbUePIzmnKE7hzt834YyCaAeB7fi+NZuElGgQj8Js12KFFZQ
q2oL5SOu7lpuGqm5yvNBMu70keH8D83dvjWkZF+hdglF/SXZtPeQmsP0/Ckb4cNydyV+P5JqJrhp
chJIaRvzXscxZE7/k3ORdWkrUgRQc9KyxVgUkJ+z/YQ2OdSc5kHhQb4D9QXcnjPswaWs3VhFGyVc
4ZTEsa7MyilvYt5dVLlnxRKGBNU7Zue/PN47kOzw+j9T1A+GhtcOKFeFf+oEn3v52/z2cu3OZfwj
h9wEKa86/UJBv9S4UV3c2NiUZXFtwISh0BNvHnhb+HEpGSPnEuIPY8c26nOLOfKPdFZ+p8hS1uTj
CIg+jQSIzq3jEd4zzHPrS0hP0EEkI50izfae5yvDf1yQ0CEJgQWIHVQcF9I4V8fx6nphq7OTFjmE
kraNERZbjxd1oUJIgNdRqdy5bb2lkxwLL40uxWuKEQRgiK2QcU4jvf7y9rzADd7bxqlKpRMcf2Nq
+GLC5VAjI4uZ7DUpvWY2+xBSbphuaUtk1G270oUR+yHhGH3KHWUOeu+EsvyU4ubNywC3OdEkMsxc
Bev3tDX0I5ZNLbPiDd2Pm0sLjWgAeygyr4FeeCxp7fVfsmvnjER+5drwkWs+M+fEmKDgKlGNxXtv
4sqSDXQ0dWx1lxsOiaAYxflK6ZugsSOTP0pXduOhSsw7xlcTTBvovUs5Zmm/uB5T3TMuxOBsnPFN
mpN0PuuQweUlk8c1FILCBzsqHWGNguCxCM0jA9T5+IdjacSlJNh83uav3IRcNQ/wl+cyLvAeO0jh
SB5E2k6NplrY7SMIhO4r+tde9nt0T5K2C6rRM89zpsEpzaMK42rgOXeTUCEuwq2CuXqOjCCra+65
QW2UmJQy9HjhK8ST+b5NDh/vODFcXl8BNmGzpOguUh2ZZyPsedsAVY1A9jHN6rFUj8rX3ofuBPuY
FVqnkrzGZ9n/8uok9yYMfqi0lGB7DlgdO3n7jl6HYw358lJbdaXxGZGlcdclp5Wp5S/yyUXBvGDz
d3tIJ2MquFDftZ2HLk5PhnKssVh7MGSVD4WpY2JWZ3EKLg9IYAz0RWsWF7pMJoHflF2TvcH6ftae
zkHdCc57/+d00qj1TVmqQHou/MIN8EhOPv70Ycpq4ZBHelrMf8xdWVdRjhIYQ6GJphfAD4h7erIF
ZaJWVruiWC3pC0peBV7k+K3oUuDDt377s9d6kmSkr+14GWia8nEaxsRi0/YHq2rYM8uOfBqUDHS4
Gylz96H1/4BuXziW8ExGucn+Apgxk86+tux6lm7nLhtvt9lqdqDKSxIGKoVeMEXCcEaMpxpJPZ/7
RARLWRr3B5jAPIf5YzJrvQe4YPryeMiUCsjnI08ykWN2880isMvSr50Lic2won8IRfDRPkUcWz0V
qb42d80NckOow+4dxkuvTYc28D4frGGH2J9Y3DMFvF+HgVIsH8KKGXfC95Xcvdn5O21Ra2T0QGrJ
AQQJ6d5i+oBv1aq8z490EfcnQoOwO/eYn6qEdv90hE6bh+uLKWxBVRxgJirj8IxhXRltpSExMRt0
LbErxYQZwwj/BMuYvEN0zoWK2e/Exl8OreJE+CI1X6WGZDDGnq4qG/pTnTFUUn+DnAaN7XO65XZI
YteIOxbQNiROu3W075CmUs/0wwIcfsikQFe8X9s2t/nfACM59h6uLQVwtcg7dyHlKwKdNJcIBLkP
GZfLNVzMaHi13WampxqUWwxOZaztyYIoewJPOno/hPFm8E5oHK4zSB+rFrtWi1S/vYwYP7bo5ZnH
UF44El27icv08lT8fbmnY7U3ghqXMdy3KPoVIytPSbqdwZSymHi7QVYwjO8njXMDcPxLcwkFpkrX
BKdPPhX0DNjJqrXZ2Gvv/m2PTW77yFtZiYszAZAQa+y0YWCcykakfdX46CZgDAJWzzEwWxUy4Zb4
O9nzJstcZIiqDaYK3MmVIVmUrL7OclMh2BnZPlxlq1haeT8pQxhJ5QnkG25/Sw+X4r6nRW6TOMLY
rvjQ5szZo4XCVriPn21JPBe2OxcetANd6FSZzXl+XF4DUk0DRLSPG98v8pTl7hUCxYZQ9J7Rw7OP
JYwhmPyneVv9aPUl6JMLqBybi4RlcSLUNtZq0ijE/0TQSVDBvtySsIIoXB9xED4kMwK/S8SHEfbA
ZLcOGEDTxgcAKr2+jfCMBSJut6ou+ig8GwRqTTsaiEJ8XyKKd/5ulZJRLek1CbnKkFQUmLC+jTAi
5SZv54LOeQL/ey6FbHHSXET/ujLqZviaRCbpL7P9tS77pubIq5vG9GQvBtim17EjiumU5y8tPbXN
GGpFqnoMjwWq+Z//1k5ybOPsg8Ur8zWWcN0pUNroYWzYvGXIjRnIq/9d2XX/lZY3j97TO9njlhGq
lPMchLr6jpwWxwno9oVdzkjsMIvfElU5WYm+Bg5A93qefgANRK7vR5tGtC5Z+KUBKjvnEXmpotqG
YqoZAOyR/Jys6/3++a+iRyRGWkhAtYqvFQrn6oQA0AUN09MRIldmNTT3ZcxaoTPuZvBvX+iBPPNd
Cs18dZEdhLs47t2rym/agGELx2+YkK3YnAMYNYaVwMDD2Hsdk3Lr3SESukb7yPpRU/QiHLdE76cE
gksiLgs+Ord5csYB9WtjkFyorI7j9oive4RnZWtW8FGJ8C1qOg/gnhCslz+8NmDCtLKsqzaW89wa
bcFzF3m6UewQH3znizFzFKx37Cxrsq9I8G3EadhiCMiueDYngGUVBsfASQo7FY5nts78JekPV+hy
ZPJ9reW9du0/7gGYXLaegVZeC0nhTpMF05RHrzUIzlDwmRdrwuUL6LM1apTrTGt3EJsys++B3ala
fAqGPEoE1boLcOsLP8ligyENn61/6EdkwpCtqsAd9MVXsGnBBApsROVO5S9pHBOne2eG6KphIddh
N5N5Mq2aHI1V8k+w3ltNSHMjZ9idBeZx01wv+3/p68lM0epfMjjRMYVshJ6q2HWWRgVPevsSUnp/
MwA0RzNkywmFmhVwhvvdWB+Jk/PkqcNdcFfSjtOYsQzkDTm0BJn6PyLoWd51Bz9cjqcGQxYm7sDI
cNiKPTlj1dQ8lIPZyrXXhrBaLG0POg6KO/VEA8Q1T9YWr3dAloKhYQTiX0JcxRDM1y3MFNfZKGqv
V9zDx3tYtsj7wgfAnblEd8UsVvY5yKWFwDPnRo336oDUa3g4bgT2gEcErkGmEI9E3I+YAijyU81L
pgJ84UDhPDTOx2TnQyzefXDVKN/waxUcGabWBq5fLLru8JjoExMBCpzXeDBR5haE98Uq80wSqbij
S51Lk9nDc+9artnAWic1DrGGDq0gXvNhtVOZyZbVECIBhMplbgvJKD95t5D7MFMsrYwTdXFwMbsP
HVNbXA3Vc7yWnwESBVSlWYiT+Q4LR+AICkLlLbPC75yj4pB7bGRfV9pAsNsZVJuVe5S0CFEOeWun
xe2RcByE37l4c2e6G97+/UOwhcb0taj0cjF6x6F4pFvryjgf3Kjyk2x05C23a2Pqx5kj+ScOssgd
deCq8YeGqZ1Xc4xdWpTcDLGdQ3YU8EcDnNe8wlsrQg/UBKFDBva/ai+n59J/Z72FCA3VyNO4ST9W
w6oJ+TdC0aJkDA9QGb61V2za0C3jBZD1RqBDpvZ3imt5ajNbjXxh+x9+nS5vmqU1JDBNoCiLJAi3
iWotqwjJpCkdCxZp67xNrHV7+mSBzFLX7FwdAL/65IroOaBUJOBal/W++ZYhGpR2qIMoMw8uw99V
gRSJc/jlPsLpTjTw1x6gjwIZEac1qQX2OLC03ev8z/QjhXIqibdP5xLA4ynfiBbV8XY54v3UzafF
oTNJ8i7NLYcQ4l9bza/ullSDeWZ2wuewREkmSYRlFFIlsXYCpUL+8LUSfypx2kEz08arUyD0iASB
KVu8Zi2Dexvokv30hiJLm4+/EFo4ZNWJbBFIsk94P6v+Y59EBrX7tJdzWZEiFUC4XgaRyR6ijuA6
T+yYEffHgw5qkOXQm9/Mczp08L/ZI0DO2HlfFdhkLBRDjc15bsZb3yXLv+yu33jqJ9WlQIhdtyok
77LvnYOwruDEz7kdGHS8LbZBs03wDBxPFTfijQAR+4ktN1z//dZtXqb8EXevXUeHsorws9tsTz+X
YTH+TN+nujUV9lXc9XoKiqFl55EbgVy+d6HPZ3mSZ20eOJteC81VJBDvK6rKUuR803l2904jRQcQ
HXQMubHflUnWtDzKfDHr0c0MqXeYVX99YuI0T4QgkPMifvO3anCOh3x6imZa0PcW27whtQBw6D4W
vToMx1ba4JILvjhVokqV1HdMoiaCAMzByAFd4ngXncAgPmyKhauFjX9J8JVd26nMtod/M4HC/PQa
aYU0gVOyWVpXUAiR9yvR35kokR7w8SuHkgKBJi7tSuG71NN6z5XrZEG3Yh7gRps3TQLjZ5Z75E0d
dePpX97SNwkUZqIPsX+E2ClgMXuFV5cNe0mcA6MJCsj8GLAmN0rqa/rbnVhz0AFmPfUoltyK5rCk
w00QxSv9qeL/JEB7yym824qInORcxvHls94TGeD/7VtJmp7iuSvyqN38mEpr89XEJ0QE6In7PRKY
mFAR9feszOcSTvQtis8ql5m8EGwWf5I0M9GO94/YA/tffigmYNsERPihfksw/BqgTPXD7P8IFel9
dYlGsEIVeNQ+imT4sVeJIHNS8H8vysfG5SWxrspxdqs/1kRYug0j7qrAX0EkWcvZPTHcav6BObXK
Ow+l484biPReFHwxiKrnY+UAcrRdzslpK62+nuIhfNEmit9QepDZAokCj4RQ84GaXKx/ZnE/7g3L
ODR5fSJihYHEqg5xT+T7bsntKqGQcJzI3w06sbzz4I+7KTWRGhuxr5gIuRmZkTcwXyRFanDo4mRg
QBnWaTw+/vqKwiiApYDMn3Opnk2FbchHVzvW1LQNAK+W0nqnJx5LEpc24oaX0FSrVUa0ZZS169Uq
K4BN95/Z1uZe9cXM6XNeZZGuAN2Tq/POx36o13TvpV+BFXvaQIhkVa8XoPFgu67YD1NU5EW+zcXq
N30kMOa5L4KsBCaCh9cjTpsz6Yj1Cr5zLHGJ7yIld0jThJau0qIJO/1sHby9BA0ZRHG0tyaM5PmE
v79r1vrQIrk8SaBpX9rrjTsjKNoC9lVwUM2tBJqsl6KNKSFzGObIUXiYzIsTx36bstPbsQLFJ2bW
VviAY+9n2NB9qu9PnnREmBTbduncnE7ZOGiXsJKTNCdTmClCdYjCvJ/v0lO8/jXu4rBeoZtd+D30
YVHVdIhEvJlSDGlPh7cUSrmKvD6lYHCuokNnerJY9pFRSn0XSB4uHEeudEPY2xgpxFeVNUMHHNMA
8oNcVkZmMR06UCzK0UKKT9GVIrRTGQoPDF3ylHt42ZaU74IImbTsWMG8SlOXFODwCC7AxVxzqVI9
DU2khBu/RN5dO7UIANx4/2JlqbJAsSkAyERDbNU/UYknKEnU/1anGFvv0M5LkMnWQ1CHl6SmYWIN
dFDDozypCvTP6eARjAvgXGhkL8bPqg1zL/l65gjHkZb7vjMpLIxx87+Asxa+c0r1eHAxU3HWt0P5
JVHty7Gdz75fdoLKB7UY27+hlhYrsV3hQfgLs9EpPWbbbB0JFplyEOyiUSEG1Zm3ILAy4tzuei54
I3jJvLFDqpDRW9s9vILKmOSXAwFERjhoPheqnAt9RmgpW26UhZK1sy+OR9vYIIJuzlYshQeu2HTJ
JpcpV5HB5fW5oAvghIo3IB2B5mkjmFmyTWS/A5aGUaNx0JPk+7trsrJ5wD7VFcVldY8C2XMLwkhM
fyorQBaD3pubFJvUALrYa3PEKgBew8n7xLvhn57Ie9Afu3IA8S8ndUccD4hYtsDYWVin+vL4IC/F
9+GA0JczyjUWkFZJeZmYwD0TquENFGsHG6UIK2UbSxp0fLEbnzlTy6EMeCgFIbqcrWgkJaGmW+bw
Z28RMNT+Jphpyhkl/4OGAXgCb7dnZKJBLX6fVol0WGTLlLY6dg5NkKY5fM9qwr/D3GgABiwau1VI
yuoamQQMouTj3EstWci0GnWhVaTW1LqhByCSROy3s/xZOxDjtjD3ss4MqAukO/T85Pprx9mOYfJy
NY0sazFv0mtcxwsosSW1PbE/wNaDceEutdybVPzw/dTeaEmCdvNTxSd7RZQEqFryjNmtOV6DSAjZ
ndEBgx5Ss1zSoVpmDRbtA34FCh5PbRvY46O3ccfhtZ6uN4Xl9j8Rb54l9PBrS0zKck3lngJ0C36b
HpcaOOwY9j6uuAxaxhQOfUgd7TwxSlOroEI5jqRX2H46hyhp7stGKcuOqNkXcWDSlSw2NT4Za+2c
gIsnG6rahkDZFppR03+a/FKepQrRFfNZ3JplZ5G1Ic6MjTBrx6j8q6UdJ1Qw7trq5mZF+baF8Zbp
4RCvXaEDqWyLCLWf3Z8KdhqdB+ypevGoPkYZJXT20wCcrZ+gJXi1I0DpILvVk3/qrs5crrMel145
rB9LBzUEc1C9SHkEmkReDgoWgkhuTU4V2OiJ+jx1UqxxEGoS2lQefcLEAqiF0f6iizZ9odMkAjIR
9u6R0W9x/UFmnfYHE+QOTSe2NPW9Z3taAnXZJ/fro6nPLB3nM3uIAi6mV7HMnlY8RiUGfXGHQVeH
Fepl8WZjPeephsv2d5Z/GbmDLlmyNGmqqLLZTn2CMJVe2c8QMB83lIHv81Ll1aPWbFLaLz/xGrvn
MfxdNKa6GZS1iTm0K7iOVxg3tD1VHOb6A1LOIWjWyK9sa1Q8CXxrst6eXFH1ExHJZT/2TRYOASYf
qjT41lVyi57XP6eK8L9ruURZGWgm8KPKFi8Jx2x1ds0aMat45IlHMqaa+JFUh8PB0M+cWYiyo5i+
m+JF5ER/ZpsdFXjcdXmqyrJwgC+RK93ERm/p4eMqoXxAj1dgjc91ucrBE+VrGBI2VC4IJGqHQJgK
jKhk6q9W5HiPz1OiWh1Ne17B2Yo9o4IAWySteAhLKd18HLXPh/pb+JaIh6arUDNc7E8Oeb+nB3q/
oYNjkuTmrMyAa5Rx89UsBDCvOgCefcsTdwQxEh0ovYRa36KItqWiL5Mu6AcuZpvflijJz3tWSF/z
AgsbSOFDIej55pdc/T1zj1CUD06io1/leMKUTzRDHuIvlA/78ZwMHQWE1d7BAQuiheh/iQG9iJSX
LbqHydFuDYAleImJidSo+bx/8wesFAoz55YUwNoU961Eb81F17bRSATkh3I9uBbhAJcmuCGhLvSh
8uyLWzkfKNHNS9LTLD6b1uRG+Fsn75j1qffKx4kKPKZqYlrs1k49Bo5ocR8kJuyZftT+louN1p6v
R3Cyd0qEYAdZoSuNLINUEZazdWmJ+Cp1nQX2m/onwCKH1WONZBDrhpdF76MocedH+LxW0DnELM1V
VhYC/gW8KBkLwTS7zBR3AyG9YtcLNQJeylfWHn/OJ3owRxpD7VZwOjJ+8ZNlCYat6fI/0fK+95C3
gxazOamTWXlPF+ai0zcwC8sdCHre5T/CDg06WFT6IZZAoJ0m0NaYXpOZmnMu6+gsXZGyol/kAGzJ
kncq5IgM85GLyaTXi1g+p2NAMniFtxDICYDFbJ1NLGSbQJ5VjyLXH0zNJHB/5HHIGdQa2j2Co+vW
A3EYj2KuWc9Bh4yELowlnwcWDeHBRqXXZZ7VbB6E4MP+cSraTrncneTh/UucSw8g0JPiChFWxiN2
ZR+FHhTRp7DpQKOGqrn3+zsOuCaSQOGMdbZOYuwmub3x9OtXw99cztbegNCvXIL32NPnd19PcVAQ
hMwkehRbP7B4M51Hj/ypg0x4Ax1Bzo3eM3LLk2Pc0r2uFiGUC3CyjxJQn5M6hDrWhtQVGuPy27gb
aMU/Ugh0NTNPdDWuJQ9knoeWOBOMlBY3PFCK0y1HqgrRy2jMzSQFVV3L5fkBRvETV+pCCvJM58zR
j2ZTX4njvmI6uhu98QAgpIBo9w1d6bXOkn41Jv5Sv6PV/WCW/Ehg7Ir1LgOQCmYEFbAfGqjlKeeB
E/d3sdxOMN39P0VAvBKuKVhfw+YZ/a6fDJxTM/l7qBHom4w4jEYVu3yaZR1b9PyWzbAtC4Aek5fs
ZsDQkLrxzLuPX78+OhnJGLAiN7rbT69Vn2YpoHZhmOj8sQeW+xHP6V1GQ/yi3nfCRrkdirS2JZzf
wOklWL6awPQzvCpdblZWb3VppeQp9ryDjcgwAA2CpXQdFQRIq/Z5TwkEyIi6M2L3NzC64svRw5mb
+ELI2bJ6jxnloPI60fTsuF5A6Mrl/BTsTk0rasETiFDgjSbzlgxE+8GKi9Rv1+Zri5mPLWERLh6s
QgdstSNteD0HopDhXdGKeZ4e5tIbHl7YetN/SMH00C1dONW2CIeZSMGMN6YrWLoLJgQo7d7t2n4e
wXWCoqSgy94u8ZSCYKaBlzTXIXEAK/nOgNB2+cDuFkiZ5dsg9jlIKelhkk35ipuUuZYqfEcfYnya
fA6qf8Tubqnr+YnnZn5MDGJQAQz+Twf8/Hbq2QOneKwJVcUy9EVCvCvmsFk17SVKSk+gUsDB+TfQ
IN4LncCwXtwbSP1ur6WS1BmDq2SZJs9lyR/AjHRb1PRVP8IE/n7WotRUeHbA+WQtiATNHEgCiLVm
PsKx0a0ToGiAToxQJ6+AAPtXGKyya2naFH37Jm07EtKuW00d/Xg1sXLfRfpZweIIkeXSUGDOnXcv
WAjpRv6ZPMDZK2it6k+DBMCWS/4c8FVvFWgzYRsGlVAYePZsWkAFksn6UpZA0H8nbhUIblma0JEO
1h7G/bbraxPMtOHNcBdOzovX3nPsFyVt3XfXtc11zJVk6rjFzBnqPFGTX7s0VAxD68m7mEaFRwRe
St1JZQgmWCfMTK2tz8KV6n4opzbRzdFyPe5vkoXQXIBRAP2H7qxg4DMRVdb1YoDemxjTaCQa34fe
A8/irOLZwmC+djkMU9MGwz/E8YRh3akaOzpW3GsZNfogYwJcfOrxS1OmdgLf65ShUrSkwc86sn/f
Zz3ku3ZxpcHP0BrcDesi5YN/ge7oA6P4w5qKb6WpgAaYFsTXH3hPYgCyqx4eJbldfTZ910rMD5UR
401aJ3ZzgvEQ+/caXeS001lpdbyEuUNeiLk0JgTF9saqwQZJh/Px0B6VspZ8+J0CHb0AdlvktDks
kHZY7oMuT8+gRa0xpBKbEZda3z7+PbvKYrfj4pyJc/CwsHSk3iMAA33pF2QXFh6eSdvJw7PDpi7h
W5A7JHLTimAvNc10JYlj0nFXsVwFD6QmgIUq7wKqKgEzUhmRaZdc72ZG1pj7E5isoecp10MupW8f
0srUb6HC3ZbiyEPLrd2nzgTo4WEIe2R4eoytSxsZkPInNK+66PW4W9ateQM3S1db20esrtPOqakF
E10f76kiqwvF5AsQMG7ZYVaS8M1fQSdyX/3a9Ius5WcP9rPwdN6E3Xu3sdluV3yq+6/y7kknhxBY
Bp4Ka3dnwhZHBgF6SHmzX5amnvNG7aSXL7pTesbCz8SlHNULgDbbZn3wp7o/bFJ/47QrxeAcYhM1
cCObtfNq08+tgrC8ZdHeyopwShICfUQZ2YZRn0ztGzzKa+vRJVZhidfX3Nu3s9iTQk8QCLznu/2K
4xQBDSVVyV43OMiDxjBAM+dIKN58BZ8JiNsSTA9fZD84+raTjyoANryvBaLfalHsH+/JFhN+lhGi
v4cKMO65vUobUgca1kMCbdNYjBbfaN2RmxhKN35IcVQe/d5NBy0uDga33PqeZ4cOrIFs7PKi0On+
ON7UVsv+GQjKRl9nEsvpNuWlwrodCKa5wny+McKo5jQFRU0PpYTGEo+PkXtElMqzKglfX9XeFTwC
B5YAjbl1eMZ1zHaZsXeIJ/wb1G0H54gfCtm3BKKKD8LCt8/2B1hC9e77M7Inan2DJ1ti/CnbTH5d
IuiRHLpk+YSsdZeKzwGF7Jjx2BWMNSNVhB8FhuoXdLRWqgIR2qlfRxP6qn8+E8aOarb0XrZ1HR93
l4jR+HmenAbzQ7+qzXP3c0FAFZqMzaL5XT5YedJk5vinFJIF4/EdvVAz8yDI9X7zrQ8M+JEOSPZg
gu3IJzPyU0eQ6Wjotk0oBcyGwvk7nKNYlMHgHNYtb0U7kW0bQPsNzMf7VJHvhFxH38OlcDO0KqfC
oDX6wED/54SHKiES45fOWNyOx79/SBTeUjWUTxxH7AdIueH6mv6u1Sa1E216k/VsXnl7si9Tap/n
bhwCYom7Mu3E/jTpdJ/WIUPP/bnNxBnm2oMtw3Y+fiO3aWQcikN5BK40EipRZwL/ncnBJVdHn+9E
gD+clCUC1HslKPU/i/Rb635ENLrd/Tdr1j9J8WBaCXEiPhekhHyKQ7N9PHdPOIxK4k4DPlcedb5m
v3ojr8WXXnU1zxuVEcTpc2nxpfhG1zyEQBowzfrI3aJh8uUTz9wWyghixu3ZJIzA/S61acuTMEzm
VQy644QePmi5cSIJ8jEOfy9HLu3BS1+fIX1wtDDtl6kYqdvPi1B2S1S9+ArwQDvMWy2cwmvkAv6S
b+1iwoKsnDDoZoPkPfQhoeidWcNw8IRwaEIfxhp+6xigD9gSfwAGkcp7crgePdFtN4WlqXetre9d
N7bRfwBzYFMBaoswsskN2vdnHEeA1G8TzftLGceLDT0Iar9lM/dZ/UMd2brkdGHCTbReX6NIXjDe
biH++35ESpwR1Rb3EIRYCMsKfDmSbLoIJNbR+wZ0Bl8IrjXsmRFIEYk9Aa736XaLCt0CT7rHmWSV
1vHGmnNT1oK8Yx9L59EgyWVKf0Mt6vIDmPEl6stpibhyUkidFn/PSrBMWAiIRbJ7xuOZMjloFbrA
yP6/UXB8UHZq9mYgZohNCOzVegFsXiPWnlTRb8kQ3V6rOKY2+vsJoDYB7PbkeOyECb6zyJ4CtEmI
KCho2fiFc4q3y8Lm6dtuUhuSb3wg3HqIwfZGtX2Uv6C3oLtKE3qK5QuGEaBi4ERhh3L169NXc8WV
ymi2kTdeof+rABYjWsICRsvtGTzwbfPM3jRDBPmhzvCtW7OpSspQwTtxzLfDecrZIhi0CUTNe0G1
c1+seRaKMghsLZJrPkXo+3CuU7MVRGwzMUdzWG6szE56PKG+GtEuwHha9YdXnZU978FRW8tCMker
WImtJqTYVcB4WmU0GZk17gW7OofcJCjm3N9sP24xg0kfy57xGo3GbOaPJ/wWPdqVo8A13ey5ba+g
0mNQ8sYGZcn5hBxgEEp1p9ZeYyuEpxQLn/tn9l8kUf+jNawg/FtH9QzQstZR+K2wzHB+K3qDNmWX
CDL96OYIK2bwYev24guA57gYjyvNbFeWkg3yhUXnXL0wGEaJUczu7dRY43IUWTkLPs/DkS8BI61s
6m2UnR+nMy7flGiGrCQJaR6LheLSr+Wp/2go+cbMu5PzAk4YIZlgFDx2LTwlnDtkonuuC++aDCV7
h7itExVl5wGE1qCgSqJzGSKmjaXjxTnsnPCK+WS/mqJfoqNruXsSk4IMUah7G2w18m8FlSx0CQ17
01qz255I0yEKLsVujHeAn6T8JOfgjE9fFoNfN9YE8DdUC8D7CwjXhNCB7+vNIbHj1bmKhjKg2UMn
AaTmHb8H05StSimrLw8qtF8pfhbk0X1gDTI0geDLl0M9fDyt3BgdLL5UAj1gSFvjMWU20v90wxe2
N9fXogGZoCAi1fbBAw1/a/LcW0hE2MWlJAoA83j2hjcRlJiRbNGQ6t58m3Wr2bm5XhoJTvc9JtFW
aOX1aLtsdGVNtl3nBd/lsMURRvt0ny4Z5oa72R3USbdZNHvPzu8FNeEKfMGpyaJPBXIkXIfZz66t
aqcQB7WRBID5ZVf1dhNGrEcbfpK0kBcAt7thonqtm7AOfs+no16T/1d9ECTsQGam2N1Pi8OPlX3q
ixr+wnApq8JEb4jo9Nye8snP30Fb0LLHlnfyNO+gyMQzg6EJVTEy/2g2wuN2omTOqG5/wiPP6xwi
e/G+5i92Z5f4qhGq8N+KfuFhDRijKbk481SbW9TmQq0Z0+HBpl35SVjImuocmWTaEuDLTNL/DwPq
BzbN55/J0kxUfcvSmFEsyFAIfbjR3LwpFNxDCBR35QlGJpLJxJ9ACTXX2Keiwd6wGZhgix4SJ7nO
9nJ7HF2pxPQ5OdB17cBDJA8zz3fXDeoTjcHSdVukl+4xVfn5yiQdg0e65I9MDlCXHn2gD3JnnPdX
nVrTiNjv5kTdQrEUBD/Hhr0yGzEiFempk0uCcPaENiLPEmT0yIUDWiX93bGTjxjgnuNt/SXKLuJw
eqpyY2axpeiGG4LELsms+aSVYO9sl9Nj1jEslBc8pZx6YrvaZDmuYTCITUGx9We9VjPp8TZw+AKn
Tlj+S5JZbaBop2yse2tlPDy4raZ2hzmg3AfoUm4/ioeGlKhn25L36/nWybWeQWY0F2IvRBAN0lvX
4bC8IW3HxV8RDp9rS18DGpZa9xMC2LgX7CK3l8AUWVNlu/Vd6LDYA1OERSn4bYQz6+y2O0daOtRf
7R4LILTfs+h0UkzTl5xJ9V2mRuJ+u7Lhe14l85uFeY5eMVY0S/NPbIjJ0f3Rm6ckGCMKy/2JO1ye
oGWTbo02lC+K3MjQKU+XXOxb9f2/2y9+h8iCTjcEMHV8JEHfRBI9dAGf5EDgu8eERUDcH80QN3Fr
z6pl10CDt9OK8b0A9nCJoRsABDSFAOpiNxIhLpy8KbISY5LhnpFD76ta8dhIGmLzf0n0LbcXEDcP
iQkGm9r3PqctuuFvyfvS3epbgaCzMIOHs6vc4BjinKsEskt+WfVc1dPYogl1/O+nqVlr2C4Nnmld
3Tj3bIXXcc/KrLyEj7RMdhsThmK2oeIPJqmqemai7kZxA03va76D3EoCAqLPvgpiEV+9gdTcE659
jzEZGL44Urb/UxuFeIHuFF0Lgr6RVMkPlQsEt0xxQUeWr/G8mE5BmJ/hJ3QkUH/i+Jx7e53D2nvu
aWz8TOa5R2nGewn4Qp4oM/nqBBVDTkTUMDruxmzZ2SQrLOnzFEsfaScX104c4qjxZBRv0brukI7d
XsLhygMRimGDZS5keRgF0BQ3E935HXbpxat9rUykUs7sRxk6Mrc3O21d30MJvkjPXLoxIhiLNUSZ
dLh7W318zeVjHYD9jf7sKu9Ap0HCfFeMbtujfLxBrYIPz7RHJy24ToRm5hIrABzAfaw/APfuT+FQ
gl3/1rURCCSVho2zYpn8td1x65RwVFmswNiwoalh9o9/Um31y+CIKY75RFSpX0ltjnqvp6if/Iie
mngNDdnOboEG5FYJxkDdLZ/uQkohCfd4IFAEtWOw/bL0P7tnLfVv4WwhwnJS5bdYRYqAEd/QTKPK
iFU23iCQI6eSN1zEJ4Q4BxGMxAEJ/zU7/HdJqkEG6Gh9noQX020yiA00O5dD60fCQaH3oWF+8WQN
wLPxioNiZEE24r45GuEKpq7JcIYev/1oivi5RFZNblKJ8ZabI4tp/fXPLDvjcO4u+xerMfl+MKpB
LAD6Mk/mswdKElpbirQpzi9j+QtWAsm1hU1IJGGDR6Qth+FZsVpbpH3UO4X+RPv0ujddIOLrvKbB
MKVCfze6Qvm4MlDqfG00dXwW+uquZAq5JoJCAHplwILui7d9BPn/uK6SDUuZWfoAg8Ues6Tw4Kdo
tb2yyu01S35bsp2E0meLhLbeMAmu/dazAzqS1REod1/cyZV/MshSPagbD54BtvXeAU5/X5rdsOUQ
FGROC+02xBmIxbwTA87EmBXMTZbU1EAQasn19WPvwfqARA9BCuxBK1UNFH5YSm0Nzg1S5v3jQFkI
aPg2ahk7tPq401A2i9SI/Pb+n++R0j+heK48jEysfApibZ7L+T8gQ4rru1vxeC8TL+i0OorBtqOn
jFBB3h/r9F8BQW0cvE5WE1uh02cJPSrjLzalrKECAd+BWz+Jo7Xm3tmZmbNgotAOEjpVde/OcIcK
PGQd+aZoJWPQUcwS+CtnN80syYcIAE/oWARpN/W9WecDDKJVQNsTxB7/5DeIibSVkLzJpH8FCuyT
KgJU+hODh64rARCuiTPbSfWRoOsHVX5dEvVlnao2fuNxZDf5u3L9fK4nS2Wwzr3Ojzxzc/lshPtW
3V7WMLTf73f6McOgTD6tmItwQXsfELmRwOyp651aS82KghQgzVzLyDZxXI/Sx+FsIAarOFbzgLIw
LdpkR/VzEv1yNk7ibaKDRh34oS5nrbOMl3mcWo/QPR+dqevBjyhy4ayFnv2BBBe/3sFNDv9WIv1V
hW7OX0stvg381LNzKJRui61FXmOmUgM2+RV1DregvCIZQg7YU+0YZ2IKOy6+zO0K3kB4NtL/nm+d
cB4diH7Z4Nq2bahaTOgrKQVpuO3XjL1ZfyeA3kyU8P3GzEV5f++bUqDWjPxGte8I1DfoBdDLL6cD
M33dkZPgSG+lARt2y67EcVkaJ2AHem3mtdWOew6VvE24Gok6XFk/7Shv8gMf9G6kW+IprwFSeS0J
61dVnh7fnTowwS3WrI6/H+KwaR4hOuzDFjSUIPt6XhMS3uhxVz4zkJhjgCVeiZ+5CuFUXy1qRvjN
zkPXl3tu1zeDgQlOvR5WtPEb/izZkjGM1euyZfydcNT3IKJDrfdvQnZAb0b7KxIYWQAzSk2pB/mM
FlRfSMLWlQcatPreCuwhngwlsAEkxTWnr8ul4gehgU+rOMAtUKbQSpffgJj9HrbVk4WQnaI61tV8
a5NbIokHLHlvUTqjrMPKf2oqx0TN6aSX/EZ2QTFZDi9I5b8nIgTo/D6nZpBhTXEBe7dYHFJglZyW
QFP3NCpMZxBUtx9Q7LCf2TxX5ypjJJxAqVe+xLCkU/PniY2Ghp/UZ7s9DsLQPbx1jA++TSS0bOF0
wcvTcTi9guCVzAzouShMTGCZ+Y110F11X61lEz8hx+Iy8qJxYCnp80bRt434QgjYILNw1puOgSnB
v/4ALmeBwaZs8V1jHBlTmderz65ue7cDxV2c/VW9Je14wr4HrsutMWC1VKufMD4V2z5UwNqnIuo4
kC+llCP5d5OTUrulaQ7Z+bSKDv/cziMkMcRtrSjlzZw/ymf3FHasNTVmw9HmSuxy+pO1yb+1LX1V
Yh2y908kbnHmlihyB8n8w/stSj7Achu2b/TD9FaCcAcO8ZKAUtHXWINXPfEQgJfhslEB415becWe
ElSa8UfNH5eVf4CFCzIlsidCdcVJWOCs60ts0LJn765Ec1Vsh7++9WmkO6RZqZD1qPZVA31JFrYn
yw/10QkFjkJDNCIVqCMgB4/igsZULELJ2nbTB/YCPGgmrLnz4UVna+hh3Eamk6exXFoSt+B8JtY2
eIsAqgEYjiuwLnMyDPwxFAhp7ckEV6wC9VAIhDemGdygPPikQ5Gp6G6KspX01NZQySn2BtifceU6
Sr0StVhcSM7zTDSXLpBRmmG8UsT7PuY9N8bJb3nJUd0I8jNJBbFpS4DXH8DVN7J6J43trQEqdId2
QQAjeKJbtGXKEq8im9m4eb8Eu8yzvxBClTg36mDc/0P8w0C65O5bjOejQMDJIQUDbHBkVteEYFyS
7wbaI5GF6w65/G9o4GUCLixenI0kZ1d/SuhQog/7+8E14XoNup9xrZi1OYYFoaW0Dg3cRsRT7E7r
WEgvxhWnps8cfRwSeMilsOqIDi5ia4vGM8jn0saOmoXz6PaOq1CPv9jtFj789yLUxyzPnmQOJ1hH
5ocBaqef4YwcPrzaebjM6mRTCe2enMjKbu0D102kXWSl0cTKA09gIc+ZvEBQ+lx0SxWTsoPQy+kN
hhcrsA0DrUtRNCISbYIOqOyzpH6M6ckpy/oBtggJhZmV3jssDh8KcCOQPat4ZskMWOPVr/qAJ6wK
r7SEh/179XPIsXVghzVvK0tzrcguLxHzM+tgyM3KJN8LylctP5tfgcDoJNPKppzlSGbkSuSnqAOc
Tlqp6q8Gblo7CVJOo9il2syK63Dd7pYCCVh+NxjhZU32aDKZ0dJk8Ahtu3rNfIOIwKXSl7jAy3Bw
9f13SrQc0d2ewFWiqRbnyCt0HC5CV81X4xrbxCj+n1kTA1j+4JyiEMtIoFISQsMaUhdg19xFiP30
qzEm/mv69P02Q0xwrAdAnh2YRCLtuuW97O7lf/s2p/QyaxRx32b3pili9lefKV8CCDZadB7rdSJg
hyCimtA2aLGKFeSIwZE1BwwONtZCWISdF3426JD5GnDHSrGJ0/SjXtErebmugaR8JHbNYubHeFQY
cNa0zlTFQOLQnar9cMPfcbty8IsYZRoVDucu9jsgCsJyfJwYVyH6cgkREp98JrDv1/Z0bPpSfMXv
XIYgYx7P3KTMEAJpmpNv+PcLaastTAFKXSkoSBqBY5kKEs4LYbGV4H4jeMd7kebKG4F2h6G/4FyF
6XCpxFcNuEZRf8nK99WwKpT9Da0UQhr4xFx4mpi14MG07dr6HVkNYzRi+AUkMTQDwqmWgZc3iosj
rxZQG4dlEmqa+2ObwMU/zP0K+gJqN5AFbluGFYOuzs65ChUOch2rBIDoMDsaGA1WT1HPeCs+w2Js
RuT3HHXyomUcYwvSnQ5FSheFY7Q45Ql6bnk3hwV1bIUxiQI2TA59swEdw9XDP5fdzI6jyoXYa5rX
21DnSDoOdLzGQX1yfL1Yc/0MT+Sf9oqoRBuCo9MVWylZcd6UybjeK3H9UJtt3cx6VpxzdSeXx3pZ
x2ubOEtb0qz8XwOiqWKZJkw4nmmjyNBTosNPw1WvAD2IBPl0Kh7Ifj5KbmguTvDA3VIySRofzBaY
ihFmeUszqYp5vwwo7Pi10X45hK4OwU6TR89EhDeX7kYO1FjlE+ddRuhZ4hZYs9I+3ncUwIjlito9
KOMDwBvMLzQ0sGUBgUsVfxMSrsX7BZOAigXlV8cmQW0yKH7XsSjDKBqB6eyn9GoiaM41Zv/wbyJ7
ZpDrX34xfP/eobuDLLq8Hmj07glg4X6od2CvuTrreYg9UzW+PgWDVImPx9IHqcLaKstpfR8zYwMs
2rfGSjtUrIFgV0hsA1y2LH1zZb/1FbMVekL/2nG3Cdy/+U3a4BUlcU3FgO2yENbDLrSH0Fw2pQ+5
/gRJ9vN9R4CCNfjh7ZQaJcfXdk1AqFJQc5rKuCDhSW20ap9//7y5i4NgsuycHoxKvL13b+eJye9B
mfI7Bbf4Sf6Pt+qhAVQcujCOQQYKfsOTXiUdNR1VwVhp5ANvV4ri4EhqhfSwdZbnjiG8mNNi21vf
wK4oxomw2lPtTRf5RP6T+n3qiZzk+4Ke+mCtMuuhu03E2R9g2M4VwtKW/yT6OWx7oylcLdpKpjNi
tuJXY5tAd4ntZlfpXO8zv12qZXeytb7lUNkaeXbeg7yNtc5k/JqJWNjns0Kf9WQU8siAT57dLSah
qKDhh1WfegvrTD7msJKIOBVJKNX4ru50EaxODVuOoqZjV28p12ZA34qlBPPvXt6YGLD6oc1wYp1Q
pDYmaQUf8N8hQpGiFPhW2O5rGkiz7a0jgi5X9qPA4lFpGCpkHoIKb1+mRNiFOBnE4W9UfMLF0NGS
x5QGWSCaGhUChxOht6Z5zTgndSCkGQdOqwudH/bacxSgAk3+ZSDRgFAT/msdQVfLLkXcGJ3PliNp
xaTLY5hRi/0hxs5S7IYkaqfOleElNOcN9cMGvTurgHTx4jRMKf7FbkjqA5Hdownj1WxwcTJvOQex
nGkuYsxALZFmxj3prUJw81qk3dQ/rDgsauEJPDZWqnuWmjhcSt25yJG9rD3kjVfYXbszYiz5A73q
qUxgcYqwSXZxbIJEu8zu4m++/t1NpmizXpkTlUE/fbzBbgVB02ksNXHGu/3Zmhyayhu6EGmeZlbU
Qq9/Oye/TzhKumr1LARQkkzEH42/NaVkqKrATxewM4khwKsAcDyw1OmpDkCErXNqsQO1DuHcQd5j
TfkSKhyjLf0gwxKZBwBD8AeL0o2QEXIwiNkYwxRfQ72vGfqaF1yfS8IV+lQNNuJBbyT/ihSbh7qT
28SpNUYup+eIs/08q40KVCfwJBfMF2QmkZm98g0fL7QPI7+/blTlrusUdwcVdRUyR6KjxMW7SLjU
u8pHKYy09+Nxwz435A4Uwt19Egmd/z66i62CjPLdP0j7U757swuW1B9mekQGPmEGhqcco3neC0D9
cu4jUkYb7dIPSdjAPmSpwZDeatPaeMBC4UBPtSxeJFq8Rm9KuntgOXGRUUAjagF2OHhSt5fqOo0d
mXwqO2CeCJUvSZ84Njnx9eKBc8So7xLX9aMOw/R9M+zHWINmUoSdYKNbEH/JNXn9ArEXnnYlA+SZ
RA1vbgRNSu/g5IKs6zIG05dh2UZNaRpq9ICUWCGTg/nDSk9FU/IvXyjarKuLPLw0e30YNDPbMLyI
U8hlES/6LgK8WtX03rqCGS9rJOoKcMVex9kSkBeAF65Ie82ZKhyuovfMOCf8q3ABpHf3ZB9lzlqF
nBOe0VbS/Z7epYqGf11iY8xgqZrLWZcMJT/mctfCXDn41CDVkEl5WCANGOOQNemE5qHlABZhIuZ8
Fnz3LoA9kmZm2xDw5OaJx1tXTOB3DAwHU0ThoPqgFE4GuNc=
`pragma protect end_protected

// 
