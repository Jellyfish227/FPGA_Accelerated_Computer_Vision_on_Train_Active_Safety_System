/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 912)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnMYaztJr9jY99iRo8Ll40uHEv0EMYecblUuZsuLkd72l7WcoUwxlO64O
UO+++pkZSFcWJd3dABenWlZxGWkpL9m7CMwaqMgu89p1ZMlbNLzZCxTxOEimrJ1y8KBwMdacc3Am
s6zgR7EzC+/g0jqOXS0ePlrTBttG7oCEYsq0INpkwF05bs97SbDSMmZUig6TAXvChyId00DV6duu
kiVbbeVB+oOc+Ckzi9fDpUbi9oN3I9k+T7PCuMOAGOdHKGZPfbzizw2IcVA/hAOC/65SWZrNrDRL
SMDaKnwJMaRaKVARgMkRml7GqTkN3EHWq7N8r/1fYipmPFc3+vLA3oCfaui9tbp/DAZKxUqWwBgp
GlaAoldlqgqmh7NRE9gaDr6dBIkBXHbdvdZISyZgiYH8mqvCBdZxvN1CAU7m6pAYcxT2ISlenVBn
KztRHzg2FDKaRr4Oyyf5Ig86XCiIgAczlbxLGWhdJQvpdsGNLltWu4+j9XbyBjN0wNgplM5jmTzI
OLo1WppP77OqrT8Oe6VGqMPtDCAR+nvAlWOgRtovANPCxNFUk1V9XDbJUV32KpjVQxpPDrDvGNme
q89sxNzMAFJd/oMrZr46G4jTghW6jMJIqGqW6H063LjyNXyhhzuTZsKlFjD2e9cXgahuyMVuviRG
EmEP17YbGgKWyOwseeS+ycflSyy0qhLUSct+E5wGel33UrSiSoseYCYhluiqITTHonsl1IJDwWjH
Qibsm+cpQRwCH2ePZQOpmnZb6m8lhydit0ezbVgyi13qSBb00+9KDq0rEMqFWuH/sed9qaElidTK
dBe7Uq3a34DC3weVVuRXWuAuB6US0rWPd2qSLtbljYZSQVhPts6jjwWHBGKnpbu/oNdj1taG2lIb
7aYBBbeDveBgj5d2wIb70AtlNIrnH/B4a0tVUeg0KQZVMWHEWb1OYcONqvnApv9LAgierTXvM+Bh
IcTdobNuOQKGQABMQM4+b18yqZg+y2Zd8NruFnVaYiN4jGrnxDLciysIIVCtQAt4RW54mgvOvdrl
GUmGCdbtR+8ACYLWWR7Gr0/z3JZknikPkpsJUPLjSda7ygRXvGgGgiQK2m9V9GIBmE0liJ1hGLMO
SVKko4STVKG8HW2qUJhV458CEV+74mW9ksBntisdHowzSSWRijSUfYEyXMY3lmlZAaEhAdDXjezQ
`pragma protect end_protected

// 
