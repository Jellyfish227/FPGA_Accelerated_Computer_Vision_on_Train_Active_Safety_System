/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnNRDwdhgvpw1C2OdNnItn2lTer0lhy5vOjhpN6hwvvmCo3Sbvbn0JxZ3
uHxaW/MGut9KL/LIeaKDY/BVVnamT2DeIVuzDh60iNsPG97+wHY8EGxEjzvthn9zBSImVG6szRhd
IWD3TDIJV5tww53iV4BAXXND8DWqn6yHrRgshlruXwGqEYaxCAJ14NbG04Co1BqLl+ckNteKcXX7
xJtqYJJsq8cgVbBxDsDfR4nD8TMJEYXYZTZYqXL6bmXp+7VtpN+bOzO4gNQYxrQAVsQy7c1wRVAr
G2iJYHd0GyLbof0lh3gb1n62rypgabvsQZ5RiKgOwQwl09Cl1iFLV5NE60csupEYuYmF1ATsAHnF
Q4ygxjWqvkJ1KD1yGO/luCvzFKtWoysFecEmVLRaXiqCPFdynzWNUBMixKYViWHBIRC9N3hWPUhv
Q1lERGaZ+A9Znv2uu7C6+3Oi/vsbE0DHFsN5V5vGexVQtNPvk8yj+055OetZ1u0MrRm3zzSSRbkc
8v1z5G+5ut+bML1pMhi5NiLaalsf/C+R93vEXWY7c27dtoWqszxirt/PEL0bMbtnY1tVON6aNzdB
cZu2phsLZPhgvJis5jW/5EA83GJwuEmWpEs9uGSzKg5EodAL411PYwZhFHeteIkdTrW+gP9o6ygI
ulyt43nvwAamHx8JAdUTECRX/IgMdfksRXlY1DsjBs8hCetumF0eihNfrPKhRYuVb0wHn7cVYdAe
n5eI5LZiEfWEAn+eeyKABtLejanVoYeIRRuBe4ZTycCoKRS8vswjPC9Pxw7TyrYmQAef8QSzgs8r
xwO9msdPTMgETCcUPO3kQgdWhApriVxp0EKx+4Kqnp+TTZqQGjBCA1lnrbXVvHJqYYVWsSD/LR/q
3TpTLQu1dVHoLS3bawnI6j3nczzOZF6msdewryLA5QWk1ihFhPhHhGVXtj9FeIG/EtCNTU5+1YNp
YwVlQOl1DTG/uHTdb9TDpBlBXJs80P4+Tm6risr9ItqCYkyhV5wC9yBkZhkiRBZX5i9g9P6I26il
RNW4m7kRvg9pOGxay8Bc6X6UqtUWMlcfQBZPStdUZd8u1Rfs5Kli8VeWLVdXmrzAOSpxTiSQmPOT
UARABPWJYMxuPbsWHIgOsTHIIyEWOsi3Jhw9pXx9HtV1QAadKv4vrXXuoAI2MftMBqfuSj0vtLU4
yjtPC01IwbUG6ahlDHbUGQkMAxSTLF1gHiiY1yMuNmC8GHU/8IwFlYAdhunekNuMtc+FRrTz0iZC
KYBW1pkrpS7MnhKvjuyO3ni8/DVpOdFI0BHWGB8b0wSRWpqtjcKI18trTIwH/3/1vrZJ6Q9+hZiQ
MkuEyMmKGkFiwICiROz+a55JLQrhVUjL1sv/xmpLFPyv0BNTRaX3QbhcGUFRMCLZZUyRCHTMyaNa
Wr69e7ug8k9Ve1CLHrgE1pKVXbi9tyYyIjTFryXfubSd4lpPZg2FBxTT8HiMYgL1jet+90W7dUhQ
QzFgRkDUp09NX0y0xEfAlpCYY3HVsLBphtKdaM8odWTm6ox2n67qoO34iSdg4pS3i7kR8bgSptAt
3J4dWSrTk2oM4lRsFmkxuA4o3VPLBYCsuunrPCzb1AJboWLPmKrsumk49lscFEudeZ7GNaMx5ugj
JwCPoDFkWth9jlHpURlWSMRR6sotzcqnynSnK01EgX89gT72msuhK5tKftWBK8PFNJY1W+PwW1TF
aPcAGarKcFoVFaYC2Sh12FsDMOFnZzJ9Gsf/smVC8mpmNUQkTXghFCDVmGJ6dJPobGsB8ZmlsMgT
c9h99EMqQzjOOpzX05y7w94rXSB3XBAE0G9NifkfxA42DEUvwAyURPnrfL99R6ahTSM+t8UxzVpS
1vIAY4bJlq4a3orhmgS8/IP73F7qDpkEOuL4dsvK58Vfjb6ZN73uuGStYIVBsxgSU2X6/36T9Mci
p5B6WFt0i0efq0KXuiGK1t50iYqiZ+OiilKxWXflbzcPRpET3gwq3wFVoUQ+SYbpzUBa5obGNBHN
jb39UhYMegPfja0P9MeRLZiO0PLFo2+6uXrTpCI8pX5aFp4m0RAN7hpayka00a1uy3dxMo+6pf/V
mFmxJrtAqguUCe7ugM5WhUyoXZZOHRXVPXEOCZ1BMj5K1L66yLaABfb1eQ+LARNacY5vesvFGEr6
vXzsT/HkPT9dBIWjjd7rP/1T/YQqn2wJNFnP5iAMtIlaTbs3U+dG9uuWR+sTneGTC2IelaEu1yub
sBgsGJoaIHPy+8PC1aYaixHiKPdvugxbGzTsMOCGioBbr/KCQTbvsH+cJ81cUsX21RrSrjbCCuQ7
aOscS5ZETawIgv1L1xCduNey+N/OmooUPzAKcX9laNEnBEnYOapdd7VIQ2rWu8NQwmJPAcanrWjG
lSSfxwLFq+Tzes5k34glcmFuAifF7aOJVi2HAkYQ1nOZMZ0ajub+t3Hw2O8J8/TdzODTnV/VEmlt
4LERyB+Qcbs6NNwS5ne17N4QsNPfI2X1hSKHxgWJXchmiJ/JVfCKBsbD13DdW1TRJHcVozId2RJ5
V4hQt7fKEAKXOkjmw2hqnRwfNTp90h+L4+IkXFw/hnLVkZG7vX/OPCm6xSkhS0P/4Su1fgdvfIkR
XYqry/ym/vh8TZ9gfbAvnR6fjo/tOaaC29nGhhGGjqQmXCFkkbCCyUqJWxSxozKngaqTwxJKlL1l
bRY0YukUY4d4+7W7jsZ1rg/qVteYUlsO9RtCHJ7tRRMTE4pVYijjThpNUA97VnF7BA/WkRvTcDFE
+axeGzb/pznDqNzdWP0D370hjTgzku4ZyYrtwyLAwVMvpvtBHDcX8BhaB0jsRYERDpLTN+/+BcUG
yMSIxZ9GJDFCXSczDcu40aiuyq3orO1PJ0ujbyRzmr/V7ginOgCPjoMBuLnlXd/Fgk0/wxoIMzEn
YM8bhMpTNMHmI6h62K1OOYe6kWqqcbWSm43Qma50d9VsUAMyhJEJG+hXNzU5lRb/xnjYnPlKyiKP
9zY07ES8MomUYRxuYDWIlbbMdWPhUsyjYam0JP3HEum3mU8J2oxZgAZZmi62iqC1q1Hkz+RLgyq4
d/0kGglKiqi6A7qnoXE8+NIf4ZrgzCXC21xV/m84RoAqCpeV5Ks9BMtw/VUHNzFC/u/2vFsWiDIM
BJi/XwJ6Zb3+DcBtj1/S+CkCHCjiLvqYxjAzibrxBTkMC0lFApTVy7kAmvaCx3VYVKy8ZAiAzsb0
Izc7zfoPduFcaYNtnqe66V3VRVICUnwQMXJvQYF8+4yj758r9+lDBxol3c3dyJKaARZkjMiiO6hD
XXGOnmSGKWzQHoF8H7X2Tbdvk+X+93+mRxr0FcCpCh6IOE5znlH9tGEu8qR5n7Pm3HwEYVYnWord
biV+htC3tSs1t3Y6j1XL1sX+kNR9/oI1blJm5369CKLGBY/lA2wDt8kVrxjUQY0NXcn7wtlYAMbV
3NGNbVdqv6yUkglncmefgc8GO/GV6cC3YEzrMuZfX54eWiq8XWHMzqNsqa6MG5cX6q/y6/K96Ukq
+XsIIUi3Z4GRTio+78Fu/D+fXbD4PMV48XwfPNvyCF3oH99OTTCqnTSc7V5pT7A4ZHICLSXKfoFc
uBwOCNgr+N3h2PPYYtApiPHHVTwDOxOXBPKT8GGyTBlxdiHrdWeN5tYnarOWen90D2kHFKrDWzr8
ZeNj7xrAiCovG/B5Uce9nzMiU2cLPEKMJSpm3JWQiIp1/INrTn68p2RD9jVLD2nbzi50OflyW/OC
9F2SMkLpvT8tF+dXD/2Y1u2Qlwb8AQD2Jb6p0HIeZUrri65PN8Kf2jDavAi3nVnhLRLAbHo8QfdJ
ujTcgTpsal2oWnPSZSXx6Ap3sNCde6/IwaW0+8mQQRzMH7N0dkU3JsH2/sLgPUcSMLnR9uLtQ4+T
k4TBVmWgUUR+XjChW3nukrdBvnb/Yh2SY1E/XD4OkIv8FZNRUIxhcA4E5TE1TNqFQroKhYW32I4A
9aqFmSzrxwoKLm7nmzbPB5JGI/1pmwh44RnNzO2BIMqGEJhkzH9+RtpDwZwDsHzBcS/tevzr5bUf
Tdtj/GvyIZbG2vVFCCF1yXVRhTguxU9ypn4CFQL09XX5/G1xSswOQDoBkiHnO2NwGUsVnieiCERT
OJNtrcqFXCS5D6zMKaQE//ye9oCCR5pfEyjWKMeEQOo7FoK+E3cKe25yq0ch550BWO5ajnUxlt3i
XkXRn/+Cgpsydykn8+b40pNuYcHvBrQ4nUwxP47pnTdm8n5aLe/otdD3yajDXLHekj9ikdi5PjZP
Rpb+J9kYE06uWVxCReBswIVImYdaDObjVqX67Z0jOiqwHXwOvO0+EwtL9befqLamXJUTwOjn5W4M
UtdlR/IDSqKrI8wpKIX5AcVB3sq/hjO+bevpYTcomCO7oVzv76iivmu/tM0S7XaA1Ki56j3neHBs
6VIpExBsOMEqvbA1wUqhD5VW8rH6vNnvXWC23ts+W+24Jn+AyDFi/3BXLr7BcU/II0nbUOwXbqsT
G6dacoVrOISZ4aGF+lzileY0L0foRr/94NeFTFIHbdvC/Nh5GXNSAY0Uc/1mDpZDbr/TLaqba6ei
HxqcJm7lvb4tP2ExNpbVm+MNW7KBtzCZ+JL/a1+Flsf7M2AUSiAalzzGSdJnK76NZVJg5OScowMe
cbeUvy71eISbvSxXkdxZxeGPx4CAK0/dA9PdmJDK5wZFhaEK27cDN/5w/3KgrIr1UtUJoMNYutul
N0G91HGNwV0Jij0Z4RMAKopyoz1VR/i8+zlSOkB2kxz2Be856S9jHOFquXZi3wga+RWKvTLPDkI5
UmUL/MUq431ALddtAvmUSY0yL+ZUrwOZm49+c6uaTpGz8Drq1tkDW7JqIReh5Xd7mKXmg00gJS4E
U589R7cMYlsEhzDozkYzjuGrxW4TliCAmAtQa3K1pPadrg09JBVTbfoVf0VO3W9UC9k1pjxKHtLk
SPBLQ1iUAKK/tI2hQyOjuJxDjTyxmcOAt1vSC/3lfmsMmdIueMIWXyTcfvoOnjm/OlC47UZUa8X5
XyQPradW3/eehIF1OxBuRK/s5o1S
`pragma protect end_protected

// 
