/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnNFv9ygviY+E25ORm9WIdE2JpGZs5olhW0jOP6uucB67Qnwi4MtkYZj0
xzODIFoK+UxbU9vvsNbZaM+z0738jvUzWU1LhqlM0YwfeP7JSiqHSWmm7HwDCgAfHueCVOogjKff
zNjIjDMBInfPVRdzg+tnvPX0PH9oEfo0imAwJaWC/fhrkuiakRCZxoqH51mslDC283kf/HuzUr6w
yqY8LSQd6Sis//5vOsHHrv1ki9kbMLkedfGfmZ1WMbO/TXAiB456deKpwSbmhNbE6emDu+ztdPDi
k44QUwAqsZZHGU3V1c1UwC80D5l4arqmdwflnVVR5DmN6FvO2fZiDJOcDM2qH2zEyykqvu7mmByT
MHWQrQ0jKZH57CTzxjQLecrWPT3uAPTfEpSBUao851t8RC7giDeLKKIKmCyqlI4tlhlnVa6Pco2s
E6PTfGqN8mS2MZ0hrGzKE6lSFStQr5dQjmVuNFsnKsmj9LYSjqgLZikm62eKPGhXIPQQ2iUO7Qi8
qCUtznjUUOmD6T4vkf69CEdAszCXXf1QkfQGW3XpXlJwg0J7a2xLfhfKuos9QLxkVe33Y3N9LnbZ
u9hS4g8VMoTI6cuMD1U2youtAaAGsJsWh+MTkf5lKzix9T4xopHf2bLrF0cWUUzU0lxccWSRh1xx
Q9vPomI16bDHUyOU3EqsT2t9J0qS/Mn5zBSuuX1kyR+FgRNUaI4GmGXsQmSG0udcL9tPgZ+6VkGu
Cw+5oZeDT30gW8188qfOuasHGJ9m8JjBJ7W96TfaTZAlwBZXUlUaYyejVEhIXLMVqAx2DgjqPWag
tGOCmZ5El2Y10eFB02aGjyXLWgoOBqY6BEG/0rwvO+jisbmMDbkMC+ofXm0Nmk8EgNDQPiOymD8w
q7gAiovXEqBdRLMVcUrxEfFlKdvYKLFQ0IdoGA8Ks7ovhCyVpXVPoQJKz6w7hN5dEV4cJI3KDtY5
y1c4nW/Rot3ZrEWC3NdN/Wy30fyx4Jhabp+YBmy3u1PpFHMJvNzWVcrpVUcoOw/3/YMTFP4PUObm
/m56Bo8F2I8OJ7nwgswSBWAnbN4XeCHPzSiN+aUCI2McxvTD8+If4YlG3uGpxGPfoSdyqOhPWikx
TXzD7pJh4FSHN0VSlNB+j/Ysis8qmcB2T7LxPV8Ce/RxLkXRn1lo1okGgE7Al+fb0nWlThL3qEmM
CsI0B7PUNvNontQm2wmhgTHgTfVt9z6McDQ4MHZfk3zIcJV0tBfERMIZwx4R5JDjg0DI/EGSB49F
wgy5wHxkASHZgvtRI8muLDBqNk058FFbpPp8sZV/DSDD2ci2W7E6TQLUPJCddE7XuAxyRnfmmS/s
AODSCChgaKVgp6z8R4lm/7HQEH0Z5/GE6I7FcsQlHiC++7X6EvzEOzp+kKXmTBVu0jjpJeiZlRql
/wWO6wg=
`pragma protect end_protected

// 
