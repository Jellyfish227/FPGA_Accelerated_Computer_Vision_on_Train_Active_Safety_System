/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 322256)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnJmU9CFjI6C7s4MBSKz3Ar17k5G614SItwyxwmFfNqTHzzYcHFCVI85q
7O4TL8DNCWZBeIWdC8j69gnFzg/YgwJvSFRkh3Y3eXZOpmrUQN9qGB2By03XWslWV8HRxRhBzf9g
IgLI7IlHmCEzBpjhc05louwtvmCE7JTBXDIsyWlIzXweB82sgnmSgEvQ7KrZUpN9mKUBm0s7R4Pu
lbo4Ot3h6WEVShwAQVhCuxjs5NMmmhMHx5jcDDvOywVBDboO+xMgmHgSkQZVo3rvKhRGF+681ShK
4icmwZIY9ayAlL0NxIh0Y9ifBpXD5WQfZshmMLmLIY2dqBIskqFzZMyUYoUYP1AujFqqt+4Fh8pr
9KHyqEQXm4pm7DDepthEIak8rE8hk6k5U2I3gLVjptwnhuH7S7IlLJAwvBFZHJ2kI6RbwIYJPgvE
5Q1JYLiX87g+vKQeEKB1sUFoul2JjUy0WtKKQsKoiIWFTamoHuTBThnQdhO2n4NF1VnqgWMnLE/c
pXU3IbOERzLYLsqCWkMK0+MTePJ6NZvDKmQo6+BivTWfePgMekU7aNPmYxtlGt5eaL9qqi87LFgJ
ZFI+e9Zb3gzQHQI0RPwxjL4apNfk70HdyQCpyvzTnG6dQ3EyoFpePYznKxhQqRoF7w+tRn2w7LtY
njKnf8kyGtYjOxz0pxu+479Ibo/o1ZMF/8oKe10ZjK7LwxH98v5YgKy8N8UZX0QhXpkueH5Z0vrn
39MhM/i3IcLBBS/jk6AMgq8NPealvX2M6pNsRA6i6lChqUofepS/TFVKB/WoA5N7KFwLxcp+VtXU
UibI9AWfwx5d8fACUZZZfxPo8pIGBcF9Rm6JrwbzyKbhOort9/nDQ2+yoQ9/8VPLpPjK4q2UkW6n
KmM9iH7XSnCgEU9k9A9Mwkowy3oBgL/25foRq8agFkbEYK6NZ38mUd7B4ReE6QYFeCxQvnvV0tpw
cmE/KaTKeVCNIvBLzq3znwHKShcZzawfuK6YOZ73hnRuIPgdtuinVUHjhZCGhu7oaJAGtoHUN9Qk
4HOMHuiTMC9zry0qd7exm0qGolV4L5pyEWZHFf4doytbTkh2j+VDy65PH7p2wcVMFg8YkRuQi74c
FwatqYsURl6qe5OJeYQbq3X7hHmDIRbM4DyxBa693W9wZ9/uFGjpIFT4E/bwCi4reGsSJBWbGBeu
Me+BQk0JCpSscV5d4NWOYP75Vg/tNJs01jm4wLr/8qFPnBAoEf8JBJg7//fAVAOkcQ0ZlD2p56Cy
nFtux/OpQ355hcKLndfCMDUV1nIF8AnbpRThFwoaQhy+g3B3676ioJ2ahu1AwdYpxmUi1e3KtBMT
JBCFk3UaOkMV3E0NYkXjNOIA+I+lHbg/WbwALj9B1CdjGaPlXkfYo4iw8T9i9sidGIgxxRXRLQBO
Ob6Vh46Iv+G+nA8r8erYEmFQdhp2J9qksSDzLNTWy+/9dsqxT7QdsiDozcpT4+5iCxkaKZOJkxUG
BUQ75XsviwQqaTAowu5cyI3SQO+DSWZzQoxuEnx0aLbv4PIFUEhbHJs09eiscgb3Rw4415i1Hogy
6zHm5Z6BFivpZMa5A9Goi461GzCJ2L3tsud9vYr6RrvdiYW2eNiDHc2znOtwNnF5U1rBgLvP0z08
6sf9zTaorFbFXlN1p+46X8YFeu7hpibYeSkfZ+ZjK8eQVe6XR2K6pktQhFBlkxDKrKcCvb+Gj1E7
xiRi6mOTTRsF/n+DcJ06hnH++ciulxImuwHvXcY9xhBG40n8cWlwX5NFegGfs7mFEKzu2ZngmGnP
YREnb4dcEzJEgyG3jJg8tdotBXL9er/rqSr91C4hFIHowerMlvYqvKFrD4eUXek88LVLtXsD2dFH
JN5nfp63RwX6hbVFKN4yCgZYFO2TES47mvEmQtNnMpWktrBtmN/gjrpY7YA2WBnggObXu67w/0SX
Qtf2N21gZSvrTxSQwrFdaYMx1F+K+F/p/R5MMOPhN2ide6TdP+WwGkRALdmpyKGYBnchM3JekXK4
KF9SVHg10cylMlgOK1TFrI5lBPh08TgMGRosHDmfA54xxfsgZzlj3fSmDlpCUrEefoA9J6mw2fSq
xU7IUodPabBLMqyoDENo3ZZ+tYjpCHbHWqYhTMp+7sT9pMyjyJpdrlqYG+OEzfhcaelhOF766FMj
LsPY3MCApoVb627+FVL8YXnZEnXouOQyv1RE43ywJJP2O19k+7uwHLcsNO+hrYOLaqMlRJAyMqBB
U0SzozlsnTGW7ZZ3L/KDx+bwz+Zh/FGoF+zTN4K6fBo+o4KRfPhUs1cB3UXor50kETw9Kfb2I9iI
Td1PXWxm4/no9YkE25CAdaSiEeOuIhfTx2WPZIURZ4b1P2ExMEoTueWRviNC7EPtuTMvrK1ELg9d
b57A/2GrfpsPMM35x5r/PxU43zHh3blFYQokLOKbbTjQus9/ogyXX16r2kmMNaMNjXPyKOy62rGt
l/Ut8ETPr/LN5oNOzJkXRNZ7lfREDuL3GIF/LGrjbUfQRdNRap4RxbMi/OzTy+B7F7/oSW9lwkjM
CmiaCHP1TaUrbb8euYyR6tOFHcoOMBEjfIhgyiaMF0JWcBN8sEu1CXfkiLIk1tZyNftIOH00xyo8
V9Sty0sFFL26emUpGa+QRMKITVS3aFn+Ne48bBxbR/ehR7TY5u+4VnGTyubUOwwJAjQzFxTsRIw/
iWZj+Gb3XM48qHKlkO3q+vocfixtv4h1SzXuCJ8toggvvF99t4Yswbgs5ShPmnkmBC2lwSJkeguZ
59gC+/3qfSd539tQubtb8RGdShdgYHSZRCf0PBixADeuDLCUFM/NS+t6O1dTRNfj/3w1bmiEdSc5
DK5lJYU02oq1m7cYt5wSMN82j19iLUD6dKpevnJSaIb/z/E/vuphMgj7iq+sHfxOAHKRyaktIKjq
aw5ctqaozKfR5V9u/BXHHQmjDasVycpdit1efks8Q0P73+DlUqu6taW0MBO7OXI+IF95tdC5GQF/
BKASgQYyGQ4fuJvB69UmnWwy4SFbTD6evw7YKyfnvyPgCCzSPwq4j+G66p+6aFpl6H8Y8UMswpeQ
/IRAYLIBHbqfbNBFlkHd8W+0sgI41Ip2mspQvpLFLmejmOpoHN5ElPK3v7wO6w72uvUoRLDA0g4J
SOtdP/Hvq2BGFVmj8r3fDRVw5k84QLCaII8V4CuHTCQ+yNBRugSL+TVUmuiSg8dG/nQM9AhIY2hC
0A4X+HEoEBJ0ReYKAjJPoC4H2Z1WZDRdQS11VIGJ6GHKNrK6dcYeTUyFZg+gcHtk8dpHDH5ZykIq
2qO6UdYdYvdSQQNWbS49/aTgaWAB6+/pdL4FQDMrqEisyvhDwMEUVlF9GTBIG3zCQ9G7sJIyx9of
7emM0lGa9JdenIIhwVBBlk2Jcv/gvae0H30dWG2BEofMJ3szq2zovHIhYpaLE+Lf6kUcFuIFC9Ef
Dh1s0VSuRDD3LgiaN0U8t5CY4vvGJpUP1mC1tcIBTa5LlNN3whzTWJyuo+V/9Lf55wScq9Pp0w+n
KkNFVZWFzogfQOuAHl37RlxbvtD/cos+HJ1Ko/TnM/feBnXryi/Zf9SEVRqbHm8uA2ESCZ7OrODC
lUFu8Or9wiGKFlQ1/5BqPuRgy41YawPxg/+bX1sSTxkM+sHitoNX3NWwxPe5VPFAVBCKo9GH1YQC
cBT1zaeGAmpMsxg0rP+h0NAqriU1W4ZIYSNU4I7O+Jx95ZHZf/3UuPM6cwmswmyOYcqHu0/BRdAv
h9RTjifdtZFKXkeUpHWdxzRemQiLHHIHOd9daBNRyVpmNZyGOMoIP3vvQjp9ynbEvl2/FDruOlvH
7HyhTOetxcuZLhjWjSazyht3p792nrEsypxhOanU4nDdY72591W/a07HY50VrkWjP/dsgsUzciPk
nEAMsdBFqYG57WAGzUXsS0EByDv7bCfYIWKFr4jzT3VaffMWv4inxtww4I899aHQvzh2SfV+pTTQ
WqbJNDyXvxu4zFO6iSJcGFiqBPxU873cEGUIV/kQMyDSrjv0ZajSxi/uHGCUNuwAZzvLpN8psGXQ
j9G8Z9Zg98KqnARWTULmcs/iTwXsmSYl40EcrhkN8r/71Uw7snlL4aeQRqxeW3pKU4XPbcDIUwDE
xn8pkxS2w9ty1rEZjAHaemdUGBf0FEia1tdnJnsQKbHimhIKu1Ak7thX9cHPqU7Rk/ItDcSTlBF2
0CbssBWk+Q/or2StummxQXUdNCCLZ0715Gh73Cq2HwSgvhOcKfuBuLP1KqiQNYCEWB/zW3avdS0R
tMryz+jCnPQQzIzhqEgaDIKZIwY5SrBWOirkWTViae3Kig2C/egHdVeSixhq3+fUenS7QjHdcJQj
+66x2HdE5O2o6zXTk4ALYlNoImZ3lYyLH4lq6lXTV6FwK9vB8dLNDcWYn4Z4DK1bPV5HNqCQ9/N0
KljF00Xlk1LZOzBZJPDGv9/fL7dyP8OwQhi5x6gPrq4qD0mFk2WUY3afAFru9pCIvgFAtjlZP7eW
zqTSM/ZKMs9271a/+p2jDYujEWkgjQwMmeomVs9xFqgb8FshbFS2bY5yDbo/IWcBIFtnmknzJEWr
wOGfP0/gITYuLoJdaOcsJjkt1qL1GYzivBrIf1Ps9Z8Hr2r/Z8Oip+uHqAqWZkRNtzwk/wMDSzNW
pAExWsWbDqwujPdF2YqAhXxnk8agYIzsndQ+t/p3EwfvP6BI4dz8C7elgyuo5dAwKceM/gOKpP++
lPp5tOPhyOoBLIhd9Nz3vebbHz7dG8GCo2jwadnNHcy/DjdXM9duPK8ZmO3kp8auuFPmjBz+sVpm
b2V57iTHLVDo9eOv2CG/l1P3AJ+dnJx3skbJVrIVYjuZnRidFxDR8fEgO49wJQNECKjneJ/QuNpz
f64oYm4BdmFG6vZ1uBonlACZRzThB7ZVGmeXxmDwyalNTZ9ptJ4kih54jf1AHSFgkbWTP39H08P3
osNBiz3MP+2o2uPINbUqk/uFsxugPChLuUk+GI/GrsJHx791yn+n+/Wn2HG6y1QMF2h2NRJb9IdU
49AGRgZAOvsWazWqbg4Vox7dSyckW/qbWF/CQx12wvMUn+Gx3M7EwEco0hl4UWZufQtvKWw1uPN8
rzVk8A3UctXSyziFD3hPIDjWSHVlKn0GxUbO2gZy5X84/l6dFJ9aAxqfdBAIA3KtWCm/fXMeqNla
uZC8eMBaUA0fEFTqcPYZmoV8SrFeg/+M6S842AfBJaOXeP1w1yXorolC9RDjc6Sq+zotdOFRBS6o
j9r/eBArbK/EcAmcwows588QrQ+gsDBq/Aj9sYbfAjR87ZWlPG8QL33cCWzUj9FYMSbQO2O0NP47
mA5zcrpA7jEy3nQaKYgBx7oBbGdlxEPbi3foEYcI983pfrp9EeI4ytHAdct1UtL947KktuL7nTVJ
yDWAwqZLZu+aBLMcuXEpSr0P67EVDl69jrcmHqzGKv8IXO2riiZJgl+9Op9c/xHGqru2SHwk84ny
a9lFrYauL1s+TJioggPXpfQXyQ76ztV+hqJz5u1IF9INVlYOGbNcPjw/MYQMRletcvgsnkKeldw3
ndxddGbQ9FMbSwGUudh7Vmw+UjXaJQF0HLAJw0SrNGeNTKoqis+QQm8QIh/y1Z3xTCx+mViJ4keq
Z/sgobPi4kiVCCehV8WEBEKwuaQ9eCc30VwvFjsgkW9DXrdOmJGggvBCqbLAuIutT4BXAItMS2Jg
EtnOcpc6NwEQn+R6Exzz7OyiSg7xH0ZC3H8fRH4umR0EL2IBwDgWYxs8eqDIkPyDxJRoaek6e1GZ
BYJy+urxsIj6kNVuL+4LPww2erTsM4A4nBOFKZHMWfwrg5Fn2+LpNxkR5z3CqRENK4jpm9vh01Hw
XikmfeFl0hDj5Y2N5EfciK3OcYiJNeP0VG7XrtPH3sm5UiUh9yT/t7MEQEzDiiRhx7Z+53eFB07p
T7vUhs7ZpTG6GZ2FR5DYIIDKUq4rq7hNR7lA9FelbNYH9lad5OEjmQ4XXxIGTFDoKmbPh8g9Vosr
6vtbryj9kKL7eXiqcnH5oMXOuU7OSaCNBglRU6T8aZ2Hpfwg1vY0zvimeTHUt0z7XU7YRBXzV81Q
0bhmCDf7ZjWMrAQ6Ja2+HXNQ30sXjwfZIWS5jr0Xkitafuu6cT/tRTe+mpHusgB2LkJGcoFx3b8Q
cJiYrsaEEnz9lYDzyOrBrgFfWcZw6MPzFOejRjL3zVjtX4+GPVZpOlqEU+UM3FerK0T73QxLEYip
Xtc6Myg3K3egu6sBErUVOdr7x0qpca0SQ0InBiD0a97OGrHcUKsKSxmh4nXPtGa561INF7xW6jFs
TaupJNDaZzSSGXqxvTPV1jbPb6alCLuNMKY2vbNruTXQtk1hxl0PFT2NfRvq/DdKiTNkfwIJOeYD
F8KxMclmRoIZkprK49C95weFoqnseFusynqgOeTgbaJOBJO8sztjPbP7z5stdXeRPf20Y0vM38+S
8HvYdBLOn1Dg3fz1emcQTwsqAOd/9Kan98DwASSsWvAGfRsuXiPKy86K14+SSM9F4Ma6vH5M9Y3x
3wt54ETjwTdIgZS5KatksHUhw0BMZIAG3tbmKazfzRWOudUlNw9FAnAQLx1e3ZDtsj89/5tukixg
1VS7ku3oWcnIxRjMWZ3yQ2wbOxPp9iQaQrsudq6NStPYjPKm6KfnGzQAnRh7cgFXFhlSF/8EtYbZ
b0e1JPQuwS7NkcLWO9Lke2/IQJf3ZcqlT7MYcCfwk0cco09AzTDaqp7hRKg8tCpooxBJ9dsvh2dB
nnPKHaOLWXEWe+dcBnUl9ct7TmtHumctTZFT04Ieu2ugFtU1S0nkKgTh/1i2h9KOjlcjZhecX/Tc
jJY1Lj+7hCo7gd3taRS8uqvHdfdqjCTxtODEk0zL0Cu9C5WGFXEDhK9AdgRTRHfT+hIOG97Hwb65
AdvhGpxKQo6ojHykn5arLKpqXFqYVlF+I/I6IbM32HSh4+bJuJ62mB8Px8ueqrKv97+GHKoxjkPX
Pja4+zA2HVz/URWbppRzu7Iv1QaduDVUZnCn3QqbEg7qUpOUj9ScKdlkDlbi9Df6+jFwrMWE3p15
RFiJLtyUm+aqnhveSZfa/xTAcO3didRR3/eL5N9HhZINHJ0bQ0G53OmLND4XamnL3hcFU5NVL89P
eGpI/5niA2pt7iOZ2U9bUknhhZ6ZmfN67wYjDMiS/CoW1V+A0XmLJTMVZoUkaNZeRLuYloExHhbM
aF4FD3YVGDlAjtdpWpy3BvoUIpcJoH+ERo+ONy2S88B652rE7NbmFRdvhjppmQF3HpCFWwUzM147
vhCfW7bWAVS25yN6Vyj2zgKDOk1fY3GkTLIzJTEFZsEhBcVc1UVnQmNuqeGSZD25wtVL4gi4tYyt
zXLMSmjuinLJhFapKnr+6CFWQJr8UqWskwY21DsfaJWvnyuYUpHyfl6bBq/a7Y9L67dda9S8TUD4
A7JECmhpGSNiAJrwTIhyGDkXm+zNSlOMHAbnCs/SNCN0A1+t1QGtqZrmGqPMPHqmfQcFCBumOgqs
EPdMBO1HNpaeapJtfd6F6RC7naTo96Un27iMfc+X7AbIyLkXnlm6t7ob0a5h8eiSoSuPh/RUev2T
2lQYuRI6FeFWXBL4EueBK/rXB9R8kWpBBDN672OrRsrrnOF89DcpngLjCVkjEh9a+tyAULDc2svo
vzwPLbY3/hSsz6hIbdfHn3hBuWVUdnvt/+fQ+ZwuyP5VCMVz/0uIjiTkt1b/Xbg7Mhlx/m8ShLXO
hLk/CH07bBW/mYqmqzXoLsnLnfHkZ8+Yj400alkw2ORUGb19vNdzZ867czGN9I9Wa8cepSI5BORE
TuQ6dQbMJiSrqVwghDWnhDKwPNBK1kmlACxOaEJI2tJtZsWYV8wgij7ePgKKfmxtm7ck3edWq2J8
dXMyTmt15Ci1Ml2yhktDHnuk5rxqIkGpXgilCYztNpKy4jYpYJnHBwE2FqlGsrvZIddI90NyEbI/
FawwKx+e6GZ75OuDhk3vM+hwzEbR1lF4ZqHNW/oS++Dn2WTXBx8x1x9S6Dzhm1hWOdLcEsXs4jet
3Ajbu4to392+Tk8qwQ4Csgxi3aNyvluIvWMvWUmmq2Xy3sYG70Ww+RBFdp1L5+CZUEbZAO+B9YX7
Zu1X7JS9AaKTrm8BxU5NPB9l2+JLMbD9Vd63gpn6uVy0q1tcsQ+jfa/E9cdTVrUCR5Tx/bVpGsRy
THnf9igr4Awadg0l83ZXbetWm+2cHWxf/EcQYW8yv3UnEE2El6RDiTjYYQ3nbWaq9OGayTxpzaBF
hjUV1rcJpm6xtDcvMOz7PCL4S/BoGKoOz4g/Mk3Oh1ZpDTQVSyR9YilI5cT/EWg/ElxBUcSpdxA/
I6TV3/8DgoahTpxqxrmphQ0/VRYx8E1T6d9nc2cwnB6OgiaLkdL+gqPCf/uidLM6NGRSOpkDany3
6TJl4pt008+CuE4zNQEje4Z3juG6nCANk55iRFyy1tvojWDGoC+OK+/begKezZNeP7xO61nP/j1Q
dqi4D8ugJV0YJTrJsAOvFZHYCGIvYGvSNU93hdI1ntOibZ+KyvG8A+KORaevisMLsh5fnQk2TtaR
qI/fIqrFLFpmrofs+kwVvfQ09dBbpczZCIJzrPR50OeUiCOrNwtcHiPPQ/enasmanfxhJ1WLxrky
tM7bGgW8FK5pUr6egRkGF6nVzoHFKfsDw2OtPutjUaRsPf02a1LznFHZZJ7V86/iPyjDALwSbrdO
HOSEgath68toKE+7VEdgzqtHScS/j2JUPxXVd2/3rQQz5iGpUeMHthe+PtVgr12rHCHTJjxPLkk+
Qv1iApnQsNwNh+FIxONLvM8W7ulxgoOezoI9v2REGd4c1tYelQjRYyVyiotBPPbP7QSMsItFkcE0
VJjkq6dPhOu5Eh1KsCblv7N2rPaxDkIxwCnMGkB35+iMUbEDQ7BRe9qCibMvO5Fh/qROKE+nzn5o
4Y7G1Y/OyIXaSj4uzIq+u3QZhxjp2QTuePDTzfljfSJJQHhnhqOhRf+P9TtCvqkaPz3FuwYrkINP
ZldHJ9qeZyx/5NfBXhRWQjpL8SRvzaT2994Dz8At5de9oZRl88+LVK0L7pr+p4u6DHg//sIOS9oI
KutAnkAqRjdnY4mOw42xmxw98FB85Qouz1rfn1Z50yv+T211mZjv1xdm+GcydR5np52x3hAwsyOr
R88qmDK+TOtIZ0hWAcPfM3e6bp0+QRJIS0fi5zDnFtCF7DVY1J9Ten+8AUfyPRtrEWBQHTwqTgZ2
NzhiGl/MJSzZxX2w9iPB4YInGZ8EzKt8nSvsh/NH3H4jyWZ5Hln2jhZvT9J0XVdc4aF8T5LbQA1h
dA1b3EdqPDdY75t7UNcBjLdIxJt9ZCJ5Bvujo3QmME4PX+3uXC3mmSl2WNVS6naRrD0qiC3rKeNc
L6pDNiQurS8zOK+KVc7HWVtzrlh58yzA5cOfXYRdUpY3onOVVK8ocTQ4Qya22Z16nyJhKgf1HJwx
5RgD+Bkda3CtUUB1/A4CeLbo7+sfk3mAXEqnoOmqkB5YB7STwWVFSgE9DE7xPD0zfQFhLX5Oejzl
iJ6R5VINF/kMpOMdL7Ewgd8SzXf41pq1Wbbf3KFHHgwDAVMJvAgP8ndJl9J26u2s2i3p3CUeVO0A
k3s4qDRpjvBCoDM4e2NQUGs0F3OlvNlZIs/Xw6A3BLS9id7RP2WkNoKTttrASAxIAF3J6sRTTC3A
LXVoqZEitV2MvKv2HqnhRjrz3n6M2OyPuAGdCq6q6DyouyyivjUsFe8bqfuR3qciinti1tRpDy1k
LVSByR/VtfSKXVEfaZ+YnPdJcd3j/wJAXzeIDElaU7TtzyFcUQQFq7mb3/B56/zjSkGeW5B2gQAp
erKQgf26GClejDP+I8neEFoXD6cLRx/IHTquzdw6pQHGMYNCoSGMaXAuhKQNnALn5tLikSs/uCYK
KPY3DTRYA/5WgwcweoOxWeOtsA66L+UIEo3Hruoj30iReNa1Cw7DX8L4tors5AqH3m1ZJlvSbFns
/L1aaOCOMioJRGLItzu8nZ5YqCuwaK1iWCG1pKXDYVIwX1272iR5fbPKFOfxPxScYMyOaKKGNaIW
55eZXTWJ9PW5NK/IGoSxbrx93VUwqSkamqOWZrXtWKh8ecyLm4OUwXUACX5ZzYRtVg/Y8EzEPGLP
al32R0xQ1ZJ+h94ux+IckZ3GHlCJeeXcv8yOq+B4hgd+BBjXTLlrCGnbRM/E/M1zzSrmM+lozSlg
b+ljfgI7Lj2AH1Hu6SgFFEkjJIVaN6FKNSoLVZjseKDL4OlkZqCAl4Km2syvia+uPt2Sztxm7xnw
hMAKs6WKj5uCy1RMcYbGpUdDbHSHhvS2R5jONXfIYD3o9JkuYvX92MLLt3ypIwdWrunH15xepKQU
raAcX75wmtv6tzo0tgYmzO7LocZZJmxsPNQI6tonbgmiyihQ/rL0/4Hp6QMj1vaAOZqj3im5+XXz
frPooTnZNoka8WfTfHupj7k3BwNmjqE5n3/hiBh94cFs3BnPyXv2UucSaCLTY8oEVXeFOT3Zufiv
qqyTjBvNFZH4uXHWw0wI9R/OZ+7jN7+wZV73ZFT9KqDGaSiGffwvDrBKM33UmSSOpf464XHwWDT7
9yxPt3iLvpmord5ZZn1XEg09q5WsKfTS15h5k7216ddDr/rbpoCBDqu1MYTPM2b91GERHrWLSIk2
VFJhHiVXTWtHVeY/VfDPjaOtjZyk94BY6D2M6yPy2DBlrRofCRX8zU0x2hQ13iId/ENkbMy4G3Qr
/3X+nCT/7NMVmTjLtMG26UHiEtbkjfqQXY8O5iWUArUZ+8t6t0QfL/gyOMzVMyo9lkR7SdGICEK7
V0fBnYIpDVsWY4qfeQq/8Pc8z7Y8Wla4mcpV+8U8wJLMdmRQ/Otc02H/uM1wdyjJudMSs2DXdn4p
9GVycOd5cuJ2u/BPuBSGCNpBKPvNPhLeHknrMCxDaS7kw0/D38pizIwp8GogIRKJdtbaC4zoZ9N5
PNpKcU2uh/jzPDH8kS5T5uBY2g5XHplWwqis2eNrqWcohO5txR+Z0yJYxDA4CFhBR9UgJulHl9Pk
iL5xP5f3QSHZOw0ogJbk8ES9O91xyt/JdOfwyJ18dcJIHa4MtVIHo7Cqtp5T+HY5iCGDf+noky5I
PiJzaOdouHR3m7+MKP+uBSL7jmg60Ei7fZw2kT+zA112iNL8Bj1qkMlYdw67YO1z+tVSCXmRmRtO
+1wz5+FlTF0c2fYme4+VQvD0BBYwbWdnxgh0qGMcS8xbaoiMRjbepjtfd+AIc2zaoNqTpUo5CNJb
sLFEpKmRzWTxn23t4BGgVG2vzfGLdiARpvpGq3WACcvw07fHfuGPXu7KwFifnx5VjyNCDhM7l8CO
33v1WlW9s0IggAYlZRLUH+Z1V5uvv1Q+HWGDHyvLNmTqwxl38fJ94D6W9QMuKX+bI1RziIWKHthH
k+tYk4n/e6tIVAwuAogwwfjQnFmmhGpDXJILtir+nkLPP5SJU6dM+r9YpVQ7NDfdIE/+A2Uxsaoc
glHtPKayaGqE36k50AQLiLJa0NRVUncVf3Fg8jApSvoBEM94VdeVQZ/wzF4I8lfgWVzllhPoIY5j
avrn4khX8l9HSpWc5WyA2D41KMpoGNA/g6fW4zqgEihVlLUe/iyM0hrN1Ovp9VmohBju0IlcwcHf
uL7H2lNcOfQMVT5FwXxHCkI2RV6t0dYwQwnytlJGQntBe4DfKlroBLsxyAIfQrwz6YGRUQtH6q2N
J6A+5xNumvB1uAFUFgRwCm8Gpjyg1LYPuM0G79K0polOxTbiBj21jdPirD0h5xPtiFkprcr40FaA
HnoLtF+8yv7Ra9wsdh32jmCiPwFsjVrsxxDRUwMifHasc5RFq+GtZrakv0MzTtHgQkxDPvHCHFcx
Ha9fVaWL8hHqO5gVSr+i+fVnX4Hbv1g0+s2enQarRZqY55dbfmlU0hyLy6uZhT6vOSgs/nq6wChB
JUlqQlj3kGj0lly56Kekbz2iMUc4E6mXHlGgtPFUDQPeLVIQ+4IOAGTNvEuwyEn7PCoBtyXJmKh0
PHgjS9wj6mw2EjFDB+BAPDbCar5WewyANZFMIT8tXNRzH512I/o0OQjR1IaCTqHCa/vLhLF4v5uo
E400kIbvaLy2Ni7d0kXlM5jBnnrGGXpWWdg/VGzIfBoOslfMdU4Ey1CFGh1xdBsfHZqR2Xmzi4vw
GVI7+ftL+81kQqen60lAMe8Au5LoxTi5Qj6kMSdMbIfdvrwEkEOTyvTeD8zoXOVx0Fxs6gQXhG6y
ZVNM63RQg0L8pL/u6P8lZQFsjtQd+4YOqROuUl3uQbRSVtOARpDmucvgydOGDZyTpX8uhXF+gLOg
Kdl9ec9KL/qgeeKCTBt2VoO08nxaWQ2fDOhIae0i5a53moFT7QeaSYOWw7TtMjez0m5tKdwNrh60
wN+blQVKX8jSsDmomU3BDIiQrNdwy6wORuvowA7FC0rzCLiWhy84q76Q6l+UkSCyIyZGRLZuDpJ+
ztQC+IyqEC+ikFSLjEUFpp88mCY41tQWGug6bSZ3SoEVrhRXUqL5wP8vc7u88/IG4RB6Wog0bGhr
pwHOlGyTvzvvrjgm17lCzxte7bA6XW0J6KTwpKrLMmT293aVIcpcx0zbaUogkRXJlmIggdacoDyY
db/ftC0xGDGj8O/osEswvsW9cLg/uTjp74+Am6iFB/iZipyUqaKcmhNgf8+J+Rk5RWsXm/sjNHpL
Q7HYJ+E5jXRRHQXmWek0LWh3jhhYKzaoQUaZtweOa2PLnr80EQXTceQwL9GZcP7THUQ7374LReL/
z6SmLjSoovh9Nk0PPH6VEoMsDb5Y9qbwx8ENIvXZdUxbvHtAhD7CqkA0P4Y+ZcapB4/b3pZXI1iM
2MqWnmP3uc9b8ZvyXlA5S6tERzsbhhBslYv2Gw5hUJg8ewVDxhH1TuC9ASJ0CRFLiUdosCn6DCId
bpJ5367QHfyrcBS15DdPWjmKrB3jFan+eHnCv+JOBaDyQxjkEO11S3dpopk8oPN1rlf3LUh6ktsX
smKL7NObPZouwouQUGU8WnS//JapeSkwMW8KJl/mBmPtGp1Vg2omblEQOho3VS+tqRGAvL7swdpx
0+C1TbJ8E2cwZyPsFJdkg+VG7/G0nhMaVmsOEIpYYe32zf6uI2GuIe8XRhHsSri/7ijJu3EU2QWu
EM+b5jgNdKBq/VB3DJX+4gJL3VROcW3lf9n/ET/jumIeuuJ+KWL6IHj+j0/gDfcCXMTaEedLY8A3
Hmm1b84vFg8mDY14UUwFz8z/RKQhUyk8EGMg0xgZG0gTKnOoeU4HeKBA8xaxyJGsQIxWEYLlV+1H
H8yzDlGdqXPSfkMs2kTq7z8HJxdnJunZT25MlGc6dhwAfPeNCXGqeavjVHz7uDFDBkGdswhUu8bz
MEwtdI9mB7TuWCGcZM895OveFyWjvjx9DCsBZbL1360btZ6gcme8tefmiiZakymNC6qVbS7lq5ty
nYm6R71cSAdmIQKMZt7oQe10Mlgn7gVUbZozrbc+JrLOKmz5aaCddVqhaiJEnM4KKQX+X0DPzlBf
nhzYEJyrEvzEJWW+KtQzQgzpXg1FIqdp9CIWwFqobWmBjdLs7L7HCO3gE8KnfO4Cq62DxjtiuC1q
1WyIaA2vC8WgdMm9Xtp7kQ0VrxOTcqrOYmU9TFZIUP3YZN6WR/KUep7PPE5Nt6e5eEQkJdbV+HGk
YSI3nYumEJ8Ulg6uskmU22nbqM9b1df1MewS47tBVRlPjlI9GBSALKeyOMKypJmqwzYXxrNG4VcH
8N97EIDhMQccpsLukFAFjvDfBgSfeljAXBiJ3akEtx18+1HVVpedngL6j+mOhRDUmiAwi8kTQ4A4
9Z3DV6LNrVPXazVWPYyb58IxJnjK2GOc4SwQ15sE0M6mr8et3fIR1oRb19IJDM6CAt1ko4PXSJoy
nw+qZTUxoqpyzCDw/6k3qVU0vky3J8lp4dSJ1Ls2x1ktKRcWnlGUfnxo0gNPiRjJ8yAij8QF7YOv
Msow620eQfRsVHKvXYVaKNkdJ/4PSgECcDnV/7ooz7EtTx3OfEIiz6bK19Gcou4WMwXMbUQYEKZv
afmE6Bf+Up5XbKDRE+gIx3X+XZ9W/f0Upavje5gCzPMD+ZinMMmfZujCiypM+c2YV0nfY5K7vZrc
Ih04vEmGcYHieCcs+YUFLhUC5RFQb7lT3rnHHWlKj+dELvlOfvbtJSlR7EMQDJxphXYerHMG4Kr7
+qCKOdKFFCLiOYnGhqIyeOE0kjvmPuL/J4T695AvhgrLGXeSG22VDSsWWcpThyvFVZ2QcGUllq3t
8NGacvFfCUCi/Vtz7kcb2toZ3Sffrwol4Hys08vF7VozfauoBUIXyL3vCjDuyfNa1bZT/l4FTRxo
uNt9ZVB/Urn9Oaje4tSPKrJcwQjYu3ENGZPHfpq1Hy98QFiEhsi/DXuvRVix0L0q8X4RSZPbvwfL
y/P5a/kU8MTem0nyTNicgxXkPjPqdZxXl9Tx2QTNhAer1Er1ENUmi+rM23kuYw1+8Tb/UgRiSTJ6
5Q3+PsHlwFtmErh+309W/C/0AA3VdjqYl/OAc27ab1vJKMY/d/VhhRZrWREFmCClrBaiS/qkDLNe
ODxdLTfZJa7a2ordJTZ3NuU33Y2AI8IG3BTHOgsvZFT2l5RH+KVxb31BJFC/sKoEM+6rFCR66P8v
FbfdGM8dnAsQgSgpgfJSp9EYNs74kTMvrfD+S1YtvScA7IGLNFpzOk7+txuDiUQf038vBWrGtObG
w7ctK0whn3NsQ7BeQ4ssC3sLQvWtohlAzv01kQEullxN4UBH39L6YcSv5KgYi3ba2wdJXDX8jybp
lTuShPAEKX4KoQJQumeid2DN3rvrvztwLyRIZSuI8fQL7DaOMOI1uhrA3DKWy/p9E8Z3YFsYbf38
GtyS/rsJuvmKGZFMu4sN6STegvUPwRz25/l51aRBgK+jpanIeglKtU3Kn5+r25CqEdL0zCl35IYL
M8OD5w53MZku+F6PSmTkr6fSBy8j+HDhK5aFkKVmwe9TRVd+06Or3i674awsc0rzMXGZN2WjNHli
GoJr2UvzNVW4gbNLu8RNIxiYLdFEoc6izmMl4lmwl3Ki4CcOkdIHTufurpOHWSiL7pdj05VJIPON
ElleJKqVSpC+NphO3kyw39MZ/sUa8Eb2qpRcc2+p5kAl3ef7uzXPNgS/cdRxxBL8JJBd9GulaZ0D
L61SQIslIK28wLdxSWTuw/cy8ZIm5TV//pEvZVKF/XXZaEioSIbgcwO6xKMgVFKkbJlpJmdjAlyJ
mFAEgKxQuCPA5RL6DlZrjB4y5TOciw9LIpknq+SDtFfMQenX/y7Nm+0kcQECO5ypkxKqOwzfDkHk
Zd+rSuuOLmy5pXnEkhBo9oXMhAUAmceqtKT515cfP1uIHzBWrmkIzFEQ5MeaJIzpWoqzuzAnOOQo
AFV/dDnaLGOav9WF3SGXk3s9LZ7dMNJAMjF/039nwS6tMkcv/CGMVYP0HlvMGYPuN023BJv6WNtz
WR8KH6jjOWe+SNC+xH1P9Xt27IGyuA+CRRucq6v5dV2whgCBPTrs6rzI7bf7gLsL8/3XayZAX+XY
MZ1xtSBlMAc1wMtDj1/1hivLoB0ohIP+2WMPwaZGTYw47sA37sFqD1/BefWCK+R84hhJ2qczQLkb
zakCDsf3dDC8mTWYQBbJ4dt/M2nc2HZNyP01k/EgfJgUFQs5zfUwZK07paPM7PJ583CVK7Kbx8h+
vi2XxIc9IP9zvjE2qcNvXhcS6DFtzApIiXWKgRVlONF/TiJuDorNMKayHOYJyDMlcQVLnTb2nWNF
MJ3AQ0gerXRJcpw3sr/o95LVMJ+HergPIPLYXkTHX7xYDNIu4C5gMUN7EASqf9/40hNTihTSicLp
CG3eEmZTpVXX20dL50ORfb+4oZSTkP9f+eg6vUw/Souem7rdBqv/ybk0apYnaCE4wHsRkYOtzdyl
KgpyVKtkNUN1QMFOGjKzpaM2Zk9OxqYp5v1asTEkvdQBPHmo35PmKqwSg+a7biOSdwIClSWcDoR4
utAvzvsJLjP6LKoVwBByKNIr7Y6F+XsB67GkagzwCuspe+r3EATC2CGEiYaGJV5AiQzKHaOndUmG
3tVVrZbkxcmZrPF+MZrtLfFeeagMy0mRtlAMeKKtwHex8LEddHw4eE4Ss9Lw4AtHXPbIz2OioALr
Knqd+aMQ7e0knjAS+26y+pJ6uD+t7MC8lfIHbX767CPiAr4DAi+jOmKdfXluUnNQponDP/SJJ/al
MBgFuGrZVxjaIO5hK0P3Qg1I/U96DydZW+S6vXtv2QlObtp3WJcLFLVPp/Izv7ri7Dze250MQy9G
aQ1jiCZo5fwbSW1VIzB/AmzjNdVsZHxw9tRljT7LUX94XURnq5eRPwx9PF1D9uKmV9H5652z/Oe6
KGMj/3aHPWzL94jI0cX+AThDlMmMiOUl96OtT3R30u2qhCPnwE1X+X+2KB/7f1veOBYotflgcZ8N
6X+V8vmtU8DvrKKZ45VGzu/Ux4vpUoifWnoNjrV87JOS2LMLNsfY6ppG9hclRQfgiKo9BeElufwA
6aL6ie9ipHfl99RCcvPeBcE62X0yNTuQzYdURb4kR87xZly+hUR9jCYXcdlxZxvnVOLH0VQJkXLy
ZFGJvl6rZC/CR49XfKtWjApJAlBpzL+yUnC59XN95NPK3I3NacPZueszNTN5318Wsb8C7v5YnXK3
8rLnGv5PnKEA+uYBj+3y2c1bs3pzLYY407KcUhN1/olOXbh6vaUS8562zAsrIVhH21NqoNjy6LUd
aP+0EmUjtwn0hHR0q0qLuDge8efLbd2LXc2TmdhxPuwDC3fJTWm8TjT7EvWxIjBDB+wsJrK7P3fQ
cY4Znf4XNpHkmn48OQcbAjrdfDWZQyDV4Vn+mMKEUcSkFaHw2anjCMN+Dhph0WJeT4TcmK4sF+Fd
t4Iy9c0x4gTCrZzxTTE7s012NvIM6WmBIG9UBA76S5XCL6tyjHA3KoULlAPtOk5LYk/3hU+GXhhX
cgIVhJrRZxybsDv9wIYeTqcIxcuCufOFEtflbAxDGQHAX/E11yclEp7Y4PceOKcYa6vN0S1f1tLD
swDrzDMbC6RssGRmXmkemRcbyOug8AUDsXWrAJpBCOr15nvmY51XRv819muNNvsZlE2xTFEGMJJp
bV15PPB/KmAYR2dtWoSkEUj/jy4EkUlXAe0Bmrp043HmgkAed5/4pWcoCq9rg1uP+T4MoaWg4EUL
vtQTJnCniUegULP/NPW4PrGL7BAjklgEKmeRYQOVlbnyLHd/7Ij8hbX7AQy+VsvU6V5o5JBomK1J
kM7rphtfXpgjc1aRpHdHnxLlLe18LOXWRmKE0NzRvq0BKAEcwyR1Og8ZtN7GtnsVuremXE2FGZi9
uQOl/6LtJVROu6F65ArgOwN7bToR+iUXq1jW+pY2IHHj4qHkygRZ0ds/DoMX2Skc46ypOfaVkc2h
EEH6WuRgSp1eLl82TGpGd++F/wZn1/36fp4zNQdLQm21gfT0qzSe78f6pcne6Seskp0nzyXvY6Ly
90BH420yZsbF1Gl1JUAUKTZAbeZxC3dSm+Mck50bmIex5Y/NokJu3vy3ZJwCmjzMr+wGGVmqzAEb
pI3xU6T9bKNbiczEF2/4CBPw2x/FjmhSCOLJZq5d4UnqivanDsz/4C3o5Z3FhIPBBeIUt9AvdTiJ
jgHicvgeL9iyluIeIwOOg4xgTXfO6xJ4FLquh9s2dUpGuc68gVcB15wp+ilpAj6kUcdCsFX7ll+V
5EBUGO9FmOZCZRG16y4MLMPGGOtZzhmtCeLoIoOoB02R8P1RXnTA0/eHQiET9VDzCG5OotalOamE
4CtAx6aNdByrk1+7sHXMeaKZ1syZn2mDo5mTEI0zZ4RlxTeSpdYsIy5xmDvT9DRmu2SurUmSK4C9
lYs7Ysh+/8Z60Gf8mzvQKvPLyfQvBN7O44xZY1BKJ8tHpuebMS+1Nt6qw/hYtrTefpqaggGGkr2T
I/U0rR4ORYQNDJNFBfA96OrX8B8X1DQOYg/2VOjYpqxFtWZqwNTItADQCb3BWe7t3DBCWlcY/4QH
/YKaslcOoJJrIQaev+BpzyoaDxbRTYCqCKtCqTHQG46j35pHld0N/EO9bxEG+OYDlHXCXSBy8AvG
DD0GHizgX1zaL/9uOQYEiIwA2mIttA5ejXEjqcD6RO4FeK+lge3zfdiF3tr6uMRs90SxMftRsWHJ
JLmU1zwmR3z5tlSn8DDAutRnX4rikoVMZwBm7F+cZIUTEoaRgvz3aMhwPtVUMpekEegxIkKxZtq8
QX2VC/B1aSohKUXviGlplmPixEY9KlPzw3AjB7lQmM8obw9Wi9++HdFOFN20cRpZ6Gm2Uq0rNdcv
2kENYix6QBGbhrGpIBE/ZILGinOMS5jLOXfBwYEkBZlKpUQFnQJmHNar//1ccAOlyB1R1Vx+rQZm
A7QhZaNR4OcQyqOSO7fhDMldtf06p5ydbqYOq+P6fAbmV42YlM51LM8zykl6bv4I8EGPtyT/1dRe
dVgO6zaH3eptsPodan29y5WPoXiK+mpIbn+rA9wt9aI5fFmXw1jqzk/vUA/nifGBNv8hR+UPL+Kw
oBvC4LSxwjgqQ0IMWJpYG2yZt3nTt36WOwbUjxPF4CXS1q++GOtoPoa8F00Om19WTpVFYlvREAde
xBhaBMtBqDiy7HE7Gf2f+YDbUw8/NIiLODPyr2vOalqUppMH2N53xb83p6YMO6SuYtHhOqsyllx8
/NBnamddaVQrZU/O0MGRf16r5RoldMYXIhro4ckPu+CGwnnKunWhpubcLp7GWRNGgPTI3jvZrlBj
p+wiOMSsf1RUmFDdLQ2LDP+uP9zLfLQ4AMGBS9QepRXBOq1CkaDsNZqGJd9Z/r+do5MQ9sGrLFGY
covX6CFG4UrUWNqV/nSA2Xhnns7kcEdXEfjgO6G2txaDujO1w+vJT1Or6NHQ+yn2JN+8AmtYbuP/
+Hrr4fJBrqnw14KdENgLOCB2iv/xgx3XpxhgnkA+einc8okv3EIApiOUhDemTATw6urUZn+lgeoU
0NrV9TGG11h565h68/byEsEfPiI/uMfE9h9hrkd4Peobj/IikOI1pxm+RuirdlPNk6B9YW+NQn/Z
wwlhOMbriTxjDZjB+rpPztuVc/OIN5RxoX5pmQmEFCNxe8xiaNQ2zE4G4WXfFR172mQfo2n1QOJG
VvzVw4r0p+SMzPb5KCcQTdA2Xr+ujsdkIlKnCO36OCI251Up2kyA0fNg7fKIXDApMT4bNONUNHyu
QiueRTfh89X24yf8/KbxcCEvWiK7VSBs6+zGbwnJFlXW+nc9kib5ByO9mAqHDIeNnOYz1wjHmoSO
1I+wVHyroORNcCmMMGh5bWR8zr+LEmcS3YTFXKNSEwL4bHULUmXICj+r1FzBGfdt7E0SiQQcrEHe
MCIQxysOv5mmE93BhpeWPYx2smrI+qqqUaX2Bzg+m9Nka7D5lQ0cAkQTKd2VPV2olUZYUlYa9TSw
+hLnRFIUcQqFaWUzaSlotvOHAUHzVVsZvYzYd75s0Q1JvzW5uLNTH/avMnR7dPnpfEamt1Bz90BJ
W7MFUkNBcuQ636XND/p5zb9SUylrHvrZxQu+EMhP0ZG7SQl+FqBm+g1ntoypYEJIQdK9ne7sMwRW
n8uuFJ6jB19sO4z4UHCWltY8yPdFnjiT7JkE61HFUBptinNOS+OA9w7frpqfR49S7NDeuRUKrn1V
efuNoyocx1Z0jGxK7q1i8buPagaSGyZnHucx3DB5+MmK1AcByj32UOOEPdfxeZ9/eoTG7OsrtS7n
QSfes+K2UetdSQ274ALQvPtx0eisnsrwIcsjQrx2TF+Gp14e2G1NoWysAE4mIbo9CJbCzBspb9db
FJ0luS9KWSEEsYh3Oy5upBBj7VqcKHYqfvCtSb2zyoY8HzBOtJNHiBx5hiDxS6T6OaLjDhs+l9gr
xSd2tLjySrLzuxiA/n9N/l098NaWj1E6ZiLy3s72sb36EZ64qeLbCXgmolkXav6mcbKLIRHdA5zg
4SXRUo1ofZrcrs/X3/WBpYYC25rgp5kkY1igbpzFjdzEWmuhXTklrPoEQQ037ksab1N7MVvgHVSP
eOikItChxjaOWSvNRC51nRN2Pl85PCXlAFoNDkCDszfyLRw+FI5geECPlStLSSk1hGUIWHACsMJY
HZOi7IB/tDyzbHzr3xQg4GBNMMWeErMvPdj6/3SFWdxTGw2kUeByiIBr+PJzOySuXNbIWpZE7a+V
+d7S1zWehVicNqXECEvRMmpbJTgF/3dU1cfigzbNC7AkJJehlItRaRON7wlZN1YHHX9/FjbQXAD8
47aDNg6KKIzuNXpUM52INXIALK6jVs+2JAXpb4Om8mmxf9OvV6bjdPOYpS4YAeHAwk37W/kMn5VH
IoRRt2yTSebK1JwUq1//nId+ozBDlcov+x9lxn2daKOd4XRJQONwedJkfU/0fMNS1nZ7pm2mAV8z
wuwvfpfixX08X/uEsj7/QrRdN6fPgmmGiN4ZUwl3UpEDYdjbWqhAnyiOQUFUdpKzokGcBYqSkQzl
sXuHOKnmqIfGvCNN67d+CbPw+PIbvQwGG6XgVSmYMlF5iqvjDOK0fHZyr2HDqy8Xl3gpOT+2Icfv
uR3AF9YRsmrA6aK35Z9h35iabkA/flAbSDSf3JxXt1nOOUUPTgAtXIQML7B7MMfM6+hIqpthJZ7H
+ajP1iQ7Tr69o6lpWl2OXjRHkmXgbOULSxLyDfdCJs17EjnlKz5Et6EmZ3tOv90l+9/Avhn1zjGF
bqHAYix5unlqJ7TnRMIUx/ocsF2E/tv88fEJ5d2GQNLcX7+thrMj0e0CWMIxT56/Xh/RbrVtVMWS
kWXofqD03xdXxSBPWe3lwOg8+w0E3sY+Rm/sBCI8vJm9UT0Tl+DtfHyZdk1th/6DaDp99zOur0WJ
Xf7ngaupNgQGv9nGceNhz6Jt/blDhw4f/3+z6UK/uW8Cd66UUO9QQ0fpyPtgVgCbQ+VxXm1DNoSj
u3d4pBXkne0IeIYrrSLSZY6si7fWf8dUPjLOBqdrTyzokyFnmU4lr143X9BLlXMXsUYwb/4390E5
6ItH6hEre1TiMYMyphPnGVvEKxue63BMz+Q3I1HuSc0aYyuTb+IkN44yb2vHwpAgXein1tJ35MCN
iPt9XxSWb14n/S/BobANuWrcmebsNkhAPkM6ZihAoO9qvsPVeerEy53nSvGeXTC7q17NpI1PyF58
vHJWJstdfx7+XKilnXzAFEzAVdcklYC5RpukkBIdmu57CG/nbQzoranPVcMIpwkpR03GhYY7Lixw
MufxQeZMmTEW4JSu7Yil2BZZL6NY/jqNg7uW1zXNwqOEIouhCRjVXW5h1/duZyf2+6XHjthfX2Gy
sb18ta1RvlXXg72sHHQtMz+ZZi2fayoicb6gRphS4dpPGpJHsYYpz3wn6uPjsY2xrWOS98M620NZ
CSbNR2Wsjp5bUifYAW/SN5L7G4splK8+3cwCGCUUsO2op0RmP7GDrhkn+0iY3S2RK9ZlEvxpBv0J
BgZ1t/Y/JiZPgjje7VRRsYmlkzDNBEDWCYiyjG3VbzFWLMnU5GrQg/Qgfig54Du4VihKzMdcE7jK
J9bxqCxvvRy+kw7/P4yeAkfpH/NhPyNw6M5+JlEszmD2jVF4PhiEQYZ4Nkmb4fHFL0gcyffEkRJv
NS7fw0BBzMDiHTvpMX1qSxaSua+67tUQyTHydSZVNVYtgqpIfrGIBOgAZq0mFxZ1cBAeUhxeP8He
aRPJcpwIzjhzSL0/AEbLLVee8j29Jv+LxhDOkAIj0J0ymMmqV7SvvayjAlQmVd96MVvNKXiAmxO+
hwElpS2nEhHAceRgf+DCOseYwsDu6ojVCuQjjnesbyB6ICUL8w0LN0yyHTp2Rn0VKk+Lvga+AymV
D/PtQKuEYUngh7MtEomR6ds0Ptdtfp6kO6GoEnMuDtd2xgS2JV1JbVroGqS0RLsJ/GK4iDRD8jmI
FkI9Hel8+ooLTmsu6KJO4II3aPoBWXtxc+f+WNU8GBJYHFFbg1hxfiR+SCpoEanzKLbwoc+VaPBx
/i42/m/YNqHYSX2KkQGOr3bGpfmOloVEeUkJFvS7kUns/Ch51SIGw8mnErDyyzO0xT7Da4DKF1de
kDDVkLntdh9YlrVEf+/zdIXRpywI01zLHC3XBSFsd7ROqO6qffioCY/uPWkhaoujfANwAb2jXgCW
YJYhAsiMF8BbpZwoToh2yiRZKnwxPMIqq2pH+127DXb8LEHdWxZYL6Wc4clEF/RaobVg1IJiKIWH
kj5pxyH2g5Ax+mfW7r2LXNoYQCyw5r1TSzbhcBmDu5MrIYJycMFhiOa7EAQGKmI8i7IvOTEezetz
ed0V9bw288awM3j2BIvlP8t6PkMv/TvRlK23U/CwV5c39tnSNoni78l+6wlu1Nt6UeHxcR15AfHi
11c7a/1i52NBqDe4DF5WFXhX7EeO/mEwJnQZK0WX7WK8CE8ctzPFI/AZ2r/64dwF94jiFhTaS7IN
1u5XapIXfkvXwEa+pslexJWW3fRSZymPwwPLTTB4o3yFM2AGuiTgTbnqglyaNswdzYfnHzBDirz6
Qu8gCAM4htxkDKiKZ6Opm/3DsWwahoxSLPMH7rmGuivaCuOduAcvvhPvNRJM1Rfe99UEVTRne/01
N8V+/1o9x5c3P5n5npoemMoOYL7MLDrHwaMZ81KDrdMjGA16dECYZSu2ch4fDuefbsZt9DgulZ/m
aEJK1rwqwCDwDRetJ0doVMYcU43qdtJmM8qHwQJ9nl+B/vCYX/rsZ59eR8hFueughZYhXUu+O2S4
8qpiu/xFrsbLbRRiDWt3UlejkInqAj3KVYz8rnzHRmxRVKLxRg1F93k+kLDJs9hnevbUDzB9UuC4
rAzqmSg/j2fAKyjF8lhWyezI1K89q5u1W+9YBZ7gh2qoLiyEOBBQrXchHCm+aDCGMQWf4YsG96jT
zvMD6PNAjlz2zF/iM3VTV/oAWMNTZJAG7keHI8WHx+izMUdAEXr1dm2j48LJYVe1MilNA83HFCAh
1oKHFbGNxTciJ5bLKa6i1BpCKFya7x0N+SXP/NsVjafKAh4sBk6Tnr8R40j8BUwizs6v+WOm7KC4
ncGCkaQpVdEPo6nkzUlIC5OKiS2ucrMi/6ZkjUTkJe7Wckj6DlMcmPRYgEUdircl89zlGbiTK2mh
KYL9vi7U46jhOlLmu4di0IUhE0vsehEAlaXXkYlScUWEbXgpfIBKJgeCCsqOBwgZz3BoqnGg55Fh
mYiyrImHyDQ+WNBuWyXGYDBbaPklPegVTwzJpi7VpOZOujzycdGDCAui6+IgzuqVlGBuY3ChliRc
creiIn0EzTtEOK2pYjunTP/n/6NYhGQ16ZsKTlQOfOacPf0WP49j9g9/UK5EBf5l1QdzjJ1noSqX
fwNQcsXKlyrd8zNP1YCcAfFaFTRnZJpFmsp73bumn/5jjM/P4jk1tkNKDiNIviS322dkol01XF48
0CErI1bbUFvO7ZNFPVgJSN93KlQ6GILq1fFP892mmDSpyTHAoPZSx3sx/Qs9sGK09oImw/KqZMFy
7Bk2WBNew5DMksAUZneEHIG2zqukHtY3qBeXu2jaz/Zq0PxPHJphUjomKVzBsmQbfYVKGEZaRa1q
7aBriQIZ7pHsS4WMIvvw9OQtIQXmUG6b7xeeAalQvhWsl0TD/F8tNNcM93nEKFUivnjQE2VQu1ju
kTCUv9JN5t6SkWoENpitkvzPu3E6lGDHJn4YS/sC070B5f7bv4jKLm9mkQQ03hTSFrjyLu9Do5yM
tdqStdlQdsogWGzgPXHfFzqFpzznEkCDSUg6sqLl4hZA47MrGXiLNcbRM98K5sPt2aj2tqm7tvVe
RrogAv39F2biCLgoOHB7Equjx1AIBfKkDkON6/MKvJ3NCaf1U0kO7HgrgXns8jJ319NrMqY5w9lL
A6mcODZW3PZWItVR14RPtlr2cWPnaF9WTw7RtAexieqpXw5Zak2VN1Oy1It1ANk/nZ2LX9+zjG6f
XlRA/q3NJN6X8U7k6yBm5Fhbd9V/U86T6EjLWu4zUrx+tFqKuUfdJqLW/c114KEMfvXY3+3SN+jh
tNXhSdeIUe5PeOayLUwLWWcr4ShFdVPVWPHhXeKYeHW/nsDqDEQwnpviimC5EFpa1NTtqJerjkFA
lhmqFrnqofmeu+NU4BpO735gsjMy65UiBUM3CI3RP6m6IpD9Mx/2LUonew3wuBBtQCsvmPiZQzEn
Ar2JBLWW/sggxAj3ZCIBmTsL2OExtAZZ/JciDqrmHJEi3rFC4l5K64uSeCP0FjQkCOF7nI9nA2R5
V8UBYFEXtsQQKnn1cLjiHNV2Wf/C2KLrBCcvdvw4FkqR/vnPbIQQEbBbI7dHPg7Mm+Ou+dShWhZ9
3evzlKBN3lSiahyn7WLKjqcjHJ9Wi1nA51QJcjT/g62jb7lZiTG9nbSTvrZaT0DrIjDq1uCYf1xO
Wgc7SqzikLS0UTgSyo11o56NTVl+RuNKUPTGZOnKfJq0CzqHgLUzD27fg0NgBlR4jWjEOM0s97qX
vZzG8PNInSarG6hMc6+c/auATmKOG7fiP3wEBswlz055YoJjYBCK1eXYaSwLxG9SFY9SSTV/px8z
tPb0311DrelUdqPT1vcq9ZH0poTmN4T/8taYrpUxQkDHO8eKqPTZ2qxTL/q3NVKx/9H7KhIf5D+s
yAmzHraYWBq9YisvtGun9jvpwrZf5n/3ruUIIqpHuQkCk8O2ykYi7IbB5uMSu4t6arXOinGhRH8h
AJoAcnBmANBuH0X1Qxko9jnBn3+ecfu+i8J/yd93qDGdf0ZxdzZpQvtgS9LTWHoXIb6APIp3VmoT
OeKZAt9zhRIW4TiCbaZ1hWFuVpjW3l7vY7OqwPsDlZ+aNaslj4qV5eyV1AEaMtoZml1jQ3ySRkKl
eo2ryFWNDJWeVqnqQf0EuYcoIEIf0l6OcklfAyuK9094pnJzDCBk3pD5/jY+WbQ4hBzF5ynuELvm
BJrGfGKj/1I8iGoF2TpR+NsHDcb7eDEc9EPZr8OmceZNxj6xEwsfCGjC+ElmDbdCCMkA65kcRvGP
RwhzuZrCEZn8U9nFIZ3UK+AGBwJIJLzeVtGhSokdR2bfaFHbcvRFKhCwhcGDwU9udTiPfDSTPr48
2zfyZaxNbVKOcaIttAx+Id+UkNXBGHSDQ5mEIX8lG9ViXIfMIJs1nweb+SyfAlHakQDBEtttecJt
i1a8msuYh3zcztOivCcKoszhNs+7MFB55axV/aDTjUa+JEOYOXczXuTEHBkgSIQVej1jn5JaDEH0
VypDqPqUlT+tCWN5tWTdVKzhc7zrcfwD0k1IKmVyz1qCihrboeuMVzsa9vkKDPn7tUiK+J6kmlAG
pwmp9/M4hsDKKnV9wWIBTXj04l/GWqxJChPqAR0+073ve/kWNYmy7SUOQZ9AHWoPVL+0GvHxEpLH
RulQ/+hlpsC9HcWi2rUgEHksA7nBm+nNFXC0P5AFyLi7lYAFHXJxeRq1Kii2Qhobcojta/v+jrJu
/If4j0XNDYnR/7AUk9eReqaOfzvxIQshD1uQ5o8vqeQSLVk8yjk/VoI8zjupDpMcC07eYmxIC5Br
8b0/C0oGQa/lzQ/8xOJmKAj396KWdktjIFzNJlKMNDmfEdk+ZA3waQOAoaN6lQ2KNApE01yqpRZT
nX1F8zeLkWpllgCpkRhLpu7o3dZ27NWrhOahooRUT5T7t7E4EF/Nzci4E4byjPxLpQvblNAB+LSY
I5DfZXUQio5AjQoDjLMhxLsWpnSH0BXW7AYtr4ppqfG7tRBWHBhYPr22e+G3CL6Ejj/RQ3yL8TIp
NiZ78aG3MgEhBTbjHBcxJI0Fn8YLXQEFwucqyjngVIXZYAX7BidFOdEynRcqH9Gx1syLkyv4Asuj
U9czHxtApxMDvnSC1TX80RO5LPIJs/JODyIv5k0mJNEleq+KCu9cY0DrvrmhemwHopLe+l9NX6LM
UmSyPm8CwqeVVr+cGxH9zb/1NpgerOGRaBsFVDlZZsk+ovWzR7QMVpGTUtqsDWnByZXb/yoBCsNT
u67lZ2B/IiMtqor3kAWD2UV0+gJ1y9GCDTiKcri+EDcAggwEpoK1DwqkZfSvuUkFkhQsoVRYRGS1
KGfRjoqC6wUPwhwykg/vzGm0H/dCscCr8ai4asJodYusjFKz4SWrXbdPi+PlmqNZmYOuxI7Sh5PG
b1YT477gLZ2Dwt6gy9fP2yYpqr9AShRecsANj+t/ZKbozhaslk2XsZdkSavNVNdSxNOV2YHZt2s2
2xRtMvpESD76MZD+os3hYtFPIEkYlainsqJv1jZ47A/L3d7HlAv0AA6pjwjkEL6eOmC1DhTPQmKr
vWm8QM8F3Hv41iGc4cEzPD/fssbnvHDvw2eOI1irWigJQwLXTxsnROJzqx/v0TANBrd6eGNqopQk
yfnnAauQ6cDXFUbxq16jZ4IqtSlgfI6a0eTAuZ0C8tIqU1DvBTQf6MJ3zAz+E/ui7JcyBAJthLDc
vUVR/X2wKprmxIRmTUcj0aqWPeOJzaINvONNmS/l40wZyaT4hZZWai7xre2CZXvDGrEaRouSsnWI
UErbopWILj4UatiymVD7lLVX0PgitJPsuddthl/2+URAls96SevZz2+IdlPrrC8idN9ZPaC1RA1R
z/B/DVp7BBikQ2oDVdQ1jiztt2v20/0kC36wZbZ28ZE5Dr5FYsLfwYdceWf5uvJkaWExjtM2mmI8
ilMhrV8DYFhoj6u6xPYzjo2rpE+9F8ZVPFMVTRK/bdikeu3x0I6K4OiR5wf8koH8WOhF+mpd+cdq
5319bipCItcydbLuSfPqNBj2XkeqSGlWbW9tD9iY4HE5RJ9l51O6aZJpYR1ml0qvd1t4FndTD/2p
1J215xW+NDoU4rAeW7RxawEKvc7XV11IW24ZmHFTTyABOuoKzEUfMPOUr2CPf9O/FuBTQhUwbsEZ
4CtUurnTv7N4lzV1+vfn8JE4YQ+UTe1U5d9aqDIUg+hnThQsDxGca6kuYASLgeFvoi1mD4ll6l2H
vb/iExSv55eEhVR/W2+rv3iuZjD53dodHBiXAzRBktDfud7KgtoEGAfDm2ufsNVRHyIf7BSHFyLq
7Oxy87kccu/iXSV7m5cOjGSSzDnTRRtsGzAxxbIBqBxIASode+GGIKdxs89IadYvjJrUJcvty3KX
nra2m6GTPmjilR4cHw6Xsj4fm8kZBOciWtIb0O1OG6t9ntDwqcak94SHitmgzAhrsBvD4kVuBXYC
RGysb3LXOaVKxCuVhNk6IkT38W0br5+tDcTdte9DJs+T36mAV9uFbDBEGtLlhp6RTqKtgfnpAjrM
p4IMD7RBOOr9UpXENbypcMztY4eJt9RwNm85I939TctkkQ8FuGxcQYiPVU9DDCxtElfDzRprHjTA
fsyrVKF/1hf4CaORXdCx+SUZQ/7pu2HEJ3OcCIJdZ1uqdtEj31eyy6nCsIdhei5uKF2uPDV9ASmm
7uA3RzWteFBgbcfGsJSn4K1P85aK4+0DeD6KWlaSiNG9voRk/+oN6nFm/mqRxG/WAvfLQAAX9ht0
O1CvRQ8rspPU9YLkarUmsQNWTxRm1z+NnwZQ3sXrWLXJAjnyuRrWIz8EgdM0dNYnL2qVl+eRQkay
g0qIJqVk93P9mIxMc/j0x97KUKKiwkOsWbFgIxmvNZ/F//2w8H2khe0wZ8SQ5l0L7l4VmgO/nr+m
ItXEw/qlva+ds6exuQ5IJEH5Khis1yxTZCOqmwcVaNn+lPvtgNnHRWY586R7tc+nWVL7IV6jHXCf
f6XL1ydRMTRi7ItYeNPGJk3zJT2oyz6O4o8C4EnyHqoSr3+evdMkjL/XH9DL2hSI2xPWcTV6yvEb
i7r+QEoymhMHwZz+gw4REBQR2OiunI8DH5RInJqplBwd6IMi73ScodHozYar7nk5AX3QhqAd0vel
U1SqTYyZsc+MDvZnTgiX7udamANIEn0s2s3HbmcXRUAR9yLz2pHZqkJtrGHJAoes7d3g84t8H496
NInSXi0JycqNhYrksWvR1v1zlg55xxFUAoePYdss8RCWGVjCuuJ6yMuwQnIkLGbr8wBA1qHN2KW/
6HAt/GB25+/tjcP8ITYvUCE1ZUCRDi76woMXvpcRBT8R2AcwV26OFtJzk2zt+adyVpf8EnsZbQAx
FZXf1aK3rZPD6Ke9LL47j2W7e8MPHzDrs3CuVD2KfOqs13MSc0wCzbk2lvh2ozKydDHLwZUmgr4b
2r57JpU94kSIrcQCkwsU1SzekvwFKXpFSsBpHs4beZhSOAFLX6lYvnu88CbRVsJ1fdJzB6F+3pmm
tSBYKbo3Oz04OC2/oOFPgpv4wK9BH04VNRP7T7LzfDYZTMmkZeBl8Bb5D0xE/8jiAKAVIta39RIF
+ZApFWDa39dDlA5khDq2ryOUd4B1hJpLnUdTqmnVtXyz49dEaadFUDZNtngGdWOaHwBDXOr3lh3C
Vxms3jPvCioLwo0IXVCiyOSxWvQit/lEUvtqj3hVYDrjndPgQJhxe5r7nl96SLReIvCtV/7VVSZN
GGpB2AGpdUcFgizI62EfRARY7mwTbRvVYi3ie6CRt3uj0GBLAbIlogTfN7sHAhPyFW+DoFKlsMHv
aeMdS7qA2GQeu6BwSt0cLa9J4cbzN5wlUGGqDuEglGhWUuBMeLPIuJKHhPFNm/RyQ1VZNIa9kfmX
+FGrGMBGmyTcC9Tkq6ydcjqj9XWNip55p80ay2/JuuG5EWwxttgHrXtLycA40l54vNlXaT35e1Yq
Zkni6qguyfS0mQLL6PuTpUaV+4ILiw/1tif4IhcfNQFeIsispJkKEtm4R2Wdx1RaN8YixDQtZC6V
2QrcoolGIoAuBU5Q8Ix5fHNgfj+chVzA1EYZPIpvXWhwUxOgcdSz8asuxbODlv4kglCE9UYPgQw+
3IXmUEyIAEwwygvnvFSbTZ+X/HU7zTD4CGjwnTCotfxQbQluh5EIuLuYsUDNW9wNMosnfOU1hRA3
p36ULEu4pT1S3h51j/GNj/Uee7jyDTS3W7lXW+6Pr8Hc9T/dLtC4R4Ez+IZ23Y79jqOZa1D8xU+r
q3RwNEBNaF6EXpm73RfsqoOtaOXUZGdGGRNKU5KHmRW7K8619Hd+V8f1vyO1ZF1aIZDsyJfE/ksk
Twj0ZO97e3bDkEMlfkqXjdLj7Qwb/JwCHQhcWKCiEpncaOP3ZkA+gobuzYRmgOvJyEuwwgt0tg3d
h+x02BfMItMf8fydJOa8oegFaEzl1vSfyues4o22LqMlSLv/nCKTodbl8e0KOKwlYUz6dVManoOd
GpE4Hdtl15nm1IUZsCpbtTSKwJqMPpYXslI5Hcj7D+F3O7aJp1XcHRVGROr2BwcRSC/6o0Ts9TfI
HniIp7L+ttQ3NOUu9o+zWZkZxUN/4WjXCEHDi1ShdgsxGyDsILJki+nHHynDL83dFC9pW/KMVH91
STYtgVVuoRBu8ydUwC9FPw3SSH95WBXEzV+CBh+I3r/VlGbxAVSj4I+bh8jX9ofibpmJKoXCSM4m
GnYDeTv1UB5LU/2WpCNefjNvWDMAuwwePvLjiTsMJ+43VJrj4+2vOcOmNdsa/Dso2wFbfBra48E2
DsIgRXI6+qJ4JQkPfZyP/zneCUIfa5/Z9A+6dRQQpQ/FY17azS+DebWfJ7j0kZUx9NEis5l/iY+e
UjQJiMYb9moeinn4Y87+Bx5wQlyScjoTm+7CNDoNnGCOrlGO5RH2jS/mh3uRnzejg4isPnleyDIs
QL27/vuJXwupu8U6G9l3ztNJUB/A2WA2iTdesfZSenrlN33CORkCrQnwajU/+QYODxob/EejmCsP
dSwAebB9ui5Xe5ulKlU+KaAUh8rc0/1keWLSZWKtfrkTdX2v9pgbhHV0Te0PNbT9rh5b2id/V83W
R+A0VIqaQGJNf2z6GxQy8O510SEtgo7WFxLIM1tC92jNTUzM+4MNJyG/ZeyV5G0N6zkLX/Avpmyb
YCQRY5Rx9obwwWPyQzieltCooM88Ac8azk+w8cCAhqX2h31p51NvEHSZWbVoJLe0S6XQ6eZj7G1c
w936EfBmqXlYiNy8EaZMFl6gGquDwhI19XzN4PnX7pNHth80U6H4qa1a1zIcepWR3xqsMv/Ivdni
1qjiKUNA+yDSjUe0xPTdZKWt6PICemqpmOK9XieNosVHxC7CTwgI5m605i1FGjSZAoAFLGuUYgb5
6OlU3HOcPBdHsPXXjSLNVPsXrme9yF/xmSdz/354TEkq5u8WgCs5llKfnn8FmS3BbWr/jaNo8+uz
Q/pu+mtb+9DgSti0zfXfqO4ClBztzu4AgRq2FWxA3IUEqyoNg2Z+je6p8Y+yKjT7BZooZjH2ZXIl
oaPsCCndUWLRCz3GhIgqIv4pjUG9DPrWD9d/wcsng0ASw3rRGxH4jihntMSj+FmaM3f7x2S+pjTh
CR0U30/RyJO/HARjGedDLRN29CSa77s6F47GT5xdOJh7r1Uws24APfx4ObCc/RRPD4lKVl5azVkm
AokMj7wkDCM20zMnlpkiamyYkAEzEKPVxWrgiF1caNFScFgg3taqjYL2eHcFmVkl4tX49Hibl7oS
kXml2T7OIsCeJ2hl2PMD5+/wZX4FoCDR2fj30jNByzZWsaHuHg4k6JDj8epAjDYkp+U2uZnlIvIq
TIcvqA+1KQ7cHV0dyhiJPcvoRZYDxw3AcJdceli9NDGfyyeBVjNF73xqnPqfFntXZEnrJBz5QU3e
2SaNc011xuIxMJh98l+VtV1tFwIM58/h0Ux2rpM+/7dN/dVeyBSLqdsD2SdURwQRXbSJv7CrU5EQ
tQqXDVD4NLP2vQRPpEuv23M9RZZwoOMVohA3zcQkMqKkKOQGn4CKDbxSlNofnUvPItBY5vm22iYh
Spx4r07MEDNhBQCvL2ujRCXQUMcKNvqL4JCF8uTnrhFXGr+R7MstBgMraLDYEp170GsjIoWcXaUL
6shoY2nQfoNDj2WA/Eyfntmdk11CpeKpZ5eBLE4FE3tM34Ftf6hwQ7aPmgiD4CvYXKvF3YnYWig6
7qOEdtJpy8s+8M+LKKbrlJKQzziAVL3NOioZVmOAue1Htly3DJWsWbheyZXb9LnK5KSlG8x9xkOy
us1TtS5gTNiO9jun+mCrbrwb4NW/GvTmKnXis5zRtRokDG6KT31JZ/kP1DMAG7mgadd5eN33vXaP
Ab2RPAQc7xO/JIvx02aGtYm+QjYt3eLphbNT8tbuv5KNY6myKIxF0rkqR3CRQpHFZ2jsKhA3oeWi
rge/L32Js2alDnet0JfPset6JxHnc3pPeMjPD3wWs7hC1gJ4tQk6UirG8IHDGCE26mELuPeFYqMK
FVXbYhH0TPsvhT2m1MK/8uRCR4xuy+uOeEZ9TVkV2J+EtwwCljdPBUoZgVCupn29pD8MPjTtkLtd
NFGa5GSXWAinVzi7TK7EkB4QKFHS7wl5HmqUJjCMuTFRu3ciOyEDpx5vYjX8DcDtD5Nw2a9ON+Q0
jD408bFB5/KwLaKvAtheCB1vNw9pzjcQIL3C+Our9KwzNrJ0v4xu5uWib5QSJLBoqGKYWxf7qd62
30mVJ9L2E6qqYleiELuL48oQ607HD+pjmlIWPkwAoqP7SwyKD1bal0IuRdEIU8GpMZDvFSgkqgng
qal8Sso0FdALnpeOmfD7jrFVNY0wIJU9c0pbr+CGYrQ081D7kTDFSK5JxiKnhTyTq0sN/gQCKBO6
NkG7mB5DzWwkImcxDEJAn4LbEUJezntx0HzusmRyrP1KrRLC+IvRkn6Wv1/tYR0QTQMcwRClWcQF
1ihwGBuk1dlMBAqEi+ryQrhAFhBNlgUlC5O/YXjS6I/bfRJxLMmwKvpp++ywj6DG3yNTaP6PIDMv
Pp4zPlsk/uWdy7qD8isNp2JTezRgm5b+nrJzdzt/aT11nnq5ZOTL/pf8MdWXBC/7/x5eiT4hijMS
pAC60O4OBcwbMXTYwO2gdZdZATmNRoohho+w9x6UihglJvNtexPc5f/Tfp0lyg328zCnFttW4c2j
V67MaIhkZ2+WVI+oB2p7u4zhLvJqAsU6yrDlBzbsaMRpUeYxtlNl8o7yWZaDfCYCyLot+Ju3f5f9
ZJpz5s6Ew8ORw/aNbU3/6MD8eNH71R6pB2qN1tVo1NId1Hmzy/3qcNMkhk4imVGiGVoFkYQZKDcT
gnvJdLhKBfBUf+j7ZUKNP/2kDw3claDK3LZoZ49hb0iLfNiRbc0FdH4rSsxo0iABBxNK4B2n9AfG
xlQHSte6xGOLT3xLr0Vc/z/3WXLDW5zG2tXXz6Rc41lhY2N4l6zmo3pC3jk2F7LFxMVbGl341vxg
d18YoRxJyDou3r5qI4woPQgWzlmZlbqIyLpc3WGawi49IU1miCfivMgdD93BR+3LDNab3XBdC/Fv
TwuY35Yi1fx3ZX3hpAtEEptDkHgl6/3pcnNkC1NwJQRmL4slAV2OU6OEE3dNzkwdKxNZhvz5W0mX
vX0NpZsi0szO4CmgvNZwTroAYx9K0W3B1q/fTgYRAlkRAUfKNYluJhTsalz72n+w8kx44iZ91vR7
ZLWPtXjJhT++Rtsi2qEe9LI8W8aKOCdYR/Ei894ik7TPSqqaCJ+nNllul0Paygh5thhWxPnpgAhr
4bIf/iJQ4xUUtUqpF32TU24WrXDfQaKL7oazAenB6ZPVd25itKvrs3jFOmOvNBCU+gXtgULLZOTM
+qLLaw7Kyl3ARzFLbwk3nZur/HZxXjTtRCqUQiJX0naQroveq+dqHpMlevJuL4wNUQwGsM0XvtQf
/COZFaZqcNk13xqjrrfoQ7PzLl8SHeOlG+63w0chLm24YVY0KHiCBIS+ppUtMdjjG2HKNiM7Wm3o
hMBauot/mcarUZKL6cSp4bBUuxqIWXY1mR9FFeFXau0jGSaste7znNshzejJCyFtfqbxoBKD9asC
gfqPC/c+w04ngGjdqP8hem//71wy1YYZxVcCvjroCPZ07a4qCKiAspImpa4CjHo48z8RJGBq05Au
i2NBIPcbafB4D3pANX4YOFQCOYJGlaO2C9AM0BLt3QKApQLqACgj9xW0nSxbdUXGhwjhjTYuJx9c
i9QK3ZgRPQMniEw5ggkblAiFPhL68J93YJqxi6OKrWhbZhCIPRE09K0U65QIIrwcVWaTqGvaQdZb
Phd+oFQav3d6TXqpBOBMTcyZFps4RRvwccxF5XzXk2+4BeeWdaUiNYqpov74vdeZSs4dem5tgjSe
FMJDIATs67kFZFJ01m1TSf4lAj7SdRqNCYlKRAEjE7bUQsr49LE2aBxSthgxA6sPPG/AvWbw7VuE
kp76T7iAKW8QEP6TJMNocdtKno6c+j50Dhduh5kGWGJFpzcd51mBPxgu48rI4KPWilY8GLQQhGx4
XZCxYXcZz8jxckxOS4U30mTKtB5I4jrLpy8yGrHFOPl5VSEtkWEuiKdRIRCHLHnMs4aB9rmsbYoB
3/wWPiUkXJWDW59/YnVAIYpMOh+RZRXXJU2SODcki6sxYbzCfqNXoaoQt70tydMeRZyyM3tphvSr
lGsil2+Wdi1ClPO0prlg3M+C2ddK/WOuOtgHgg3f9K0UKPfRtjdBPMkSf4ICkdnbrYjfLyHe96YH
aW6yhtPwVNMrnlCDsrMPEXYgL4qSGod7JQl27Iovh2ktXr/k7zlypAVgcP9oU1j+vlZJzkxhIH/6
FOpA7aGehDPdxjk3NL2fJfm60hoF/3FqU4umkqMxOPGOn+ql9XdsneQ5f9kQ6cie8Jjt6afk16bm
vAXKCILp2RWDDQ3bYcXIM4ixnmd7ZhTBKt7uNwfoZmilrjOIrPItOVPuWG7k9hrrvtF3ovgNDBwT
To0Yx87P71dJ+VFG5ZTbqq1cSC/Y4aLY+8ntGgkoZPIk7sXiLCD00ucwH4UR2HAydpVzJhXYx7mC
/TJMvuFdXklzXhHTFv1jb5fmg3ZGhFYGn+hv266Q5oHaBdJe0+XguXWxnARUYwCuJZaqXSRgOfbF
ed/owgJgf1Ih4HB/7GmUvQixgwUudoCmN3YyUe/iaJoxen7tEO8buBH7+uoXW8nJJ/YGRf71A3JJ
yXSV+KqUcCyUbBrtbz9/xe5pP/lWfP32PTbVnk54RJe7GJk54Oy5KownUJn/BXpwGr6B7MMvdG0V
u7v0PvzzAhjm19MyzYpnITuwGaRgksS9HwWH5yOGCmM0+8F7lY54gkXgUj6H7p0myobZlOV/q9tt
zL9o8Z5+dbIPQnLstKjnMUUx4J+Kf1w0omSOplHzvo53ZmftdE0Nc2dOv9a0cjQHMzMWeYh4jPDi
I/q13ZbX+6/JxTiPVAto5D2fzL5K3X/biLOizKEnnuqWnWjXlEhk8b9ar79/G2xkIcmGuPj+8Er8
mEh+XItvwDuEoVQeO6VFs9DlMLMwEqV+SbQjVvMhNWkRcZ5y4D3YdAgoV8TnuMVB+YAu+JbjJupX
ES0DlIfK1vjmI57Skdcm/S7pa3I347PCjXejFMJwynP8QUui4UytFSB0sBicps/ob5GzuwmaYllK
sVCSJbYQh/VE5k7OkQp0SdmQrBauONiLcEAeUSTj4E3LvJIILXoH00S5AuNSl6HzNFcnbYP/3nej
L2f1gxEgFOnihl9Zkvyk1f4fLWBiv6pg/UNJd0POHvYSBdxKHsn5taQkhQ/3LSbp+9un8uSVIIh1
T0qGFu20fz5BeUXlhecX4NhtP9FVGdVR+vlIJCeylO4zkTL7bZ1Gt+VLF/mp3uao3iG6ltzPCsvd
zAW615qpuXcdyNLzltsVdmOcFf5RysrHRas0QNxU+cwDwpA+0uYpuPktfn9jNHjVSm9HoFTHeTDz
Up52e2dP0WdjDJ9maBQUyvjzeEVBfu0ALX/eYmmjdbdUT/hH91cLRCxGyRyAxCsNLDBJmT4rAVdV
Kr/ja8V2jO1MJ1XVzhUxzdrkrF70dJFNrh2VvMxRtiFAYbEy4AAn7u/0pJmKsUvyilxWVmCkTTW+
d8yxSGdHP0jUG3CPdua2pTx82icvO7xwqcEH3d42kJr02OD4Zk9/MkXAQq/N8p8vW8nV/FHd8Iq/
W/J0N7ohYReXp1I1NP1ajZzPxY93eA69vGhisW97Df87yHRHIV/IHMFmNz1LkmhMTT7I/OYYA5mz
KnwlxC5F9YehnjbTD52196B0L4EwAxG1KnjFYMxlNt3E8q9znuDm72BmbRfIeuEeqFWjed3f1YC8
cRCa5TSBB3A4wKjE7Y4SJmtn9qSliVv5fHiMBcU9FTvTdjJ5wRTlT343AHwP9L61cq5De1aYCql0
EhJE2S/cTLHmhkh3NCTSVPZf7gb6orbiR3ApijRIRyslUBRu2yEl1u0yxq7hGmYVARNOCMOlJxUj
PvC4/cbKyaODegHGoxSSHPtf+KoONjR/Hx9+WnSsPXNt6J/llyUY6GDiB1uh98PEfcqC2HMty5su
Loqn1puBf0wTcSFRdY9O0glbY1aTUBRd3DcIs6Q1W5mCZe/EtIqU7yjnjZ7+/GbJs97H34KtDD2q
upZBLXkgQjorOSnWT6oPrIRqo/pZSCDvFpFSLCVmzDU3xlPkCPfMPz3XYLiG7je7cWPTV76ubecF
+oU9Vrib2mTJe95Rkc5rPBLk/VWMACAhC35pyLeipc9h+CGdjfaK37N9UJXMO7uHrP26OOSUM/0j
MEz6Luj6TM+sTNZJHwW4oS/zmVtD4tK4vhlgi7aTS3efbRndAMMhx9IrVXSqIKEDqXFbBRz39uIH
LLVj5rZFcJoGbjZ5XlKTI1NdRGWGYspdl7ku0yASrs6NKMAlQ6+q5Bb3ib8L9nTUbWS4c71//ARo
hIgg69sukonNxrX8lrNHIdKbHgoI9HZkSWkKxJAH5BEalGgtmAeTInjkdw7kpkGoW8wXQxsSeFv1
D5sThUkr8gvOlDHcv6y+78I4nmkXvHIOm0TLc6Mq7e0Pii/DHdcUf7tK/LB9GKobsrXbHPqrTInl
wCjkblgp/I/dvAYPSXFFqgw4HfQbYV2E1H3kroeVDoiFb4HTw7RQ2joZ/mvUmFTz7QW76pwINwmy
2dF7PMruF/tX2wcKzz5womqnTdTvfnfxSd0f0zsybDoJCNwrbu12Oik1LutzaeN8bXGJcsy98y/M
QtWWlHr9Hkg8MrV9l/IYtID6Kj2p7HPf8m1mIrYpNXdpFhsOTDocwZJLD1pmv4kfcvZHkvWW+0p1
lhEpyFp9xk46EODm97/E0phJYVAILo9Jfl7slzgrJoH310aiEgGit/bCD6OqwOReFI5FZ+oghAGu
uud1/5s1cjTjSrHRewyd7o01HfgLfOiskksyjr4OI1cIV5aSxbMq/IVqTUFf4EDjQvkghd4zEbND
+hcspXkwrkIOi/IxlIvlWte8u2Sfd4mhtfivG/9fO8jCfF3Z883CBAyy0NMCoVQRXBujlkYVZ1FH
5lje/FZZtu2T14FWaNnCfEM8OYqsnXxlZYIgeRRd5Dvw5p4lR1tdXezaMoxUiwTG2GRugKuWXhK9
V23nI+lS8a0+RGk+1fcY7pLhoh127lhHmUwRIczBB/KNOppWgSjZN2yiqYjLe1NfvbeGhIDUoLH4
FY6tqR8Cd8rL2Po/7dLcXCG8KxAS+UGeWIO0+xqqBAXhFJe2TFzUvaTA1Zdkq/pwPJL69otXnMYV
hxdGywzw6qZqSDwrj6VzZuu2p+ZP4JBiAWng24jnd9bxoUauoiUh5euNERnl0rIjZcUBSwTA882H
tyuDXmW7a7sCphMTWhTPEYhvz8N8ZqrMif/h6F5vCBoaLGE9EtdfZgcxg6XO4a7fqx2NTjnlYkdi
9vV0SSeT1rESQZ9mEVv5WsLg/dgkTcE9I019Lm4a5PQ6rE0LZwujC7qkpNPN34PXiOEyO4Crm1zj
77EOGOuq9ZAlaZ5qKpIB+7J+MOljsFUqjEQLUbrIIQCVxH/y2ckOl2xBBJsgsowISNwV9oBXj+T2
RB2HFGsu2gCJ1mnCICN2iYWWmNrCs89fcdvpN1QCRC8k0C0f2nrSVuryv/Vo7QTBzwQ7ddA/tqPI
CtPgx9oGogRRO0SGF0lz5rSGvYnCAOBbWe/onIsgcbHYlJbHMk5Stm2y4DoP3ND+i081Ncqoecw1
CG+6fc3H77fcJ9egI6y2/GqyLBy9AuP4JuygmfecFD4iqe1EusvmDmm2QS2Bzhvn+KEM625fDcnl
0eTdlYFuRXQtsyz892ws/nesNhPDJcrrPw+FH0/uySnYx76FiGP7F7rAKJmX981ZbMTRp3BFpoXn
jM/007hK66QQIQPFDRpbqAGR3qlld0FuQtR372gqvzWihK6VbyJGuD1pG0cXc0aWXxxedPhy0T/w
taQDdwKpQSgJv2j4Z3fHPuV342HgSVKQsUpkY6RR3ZCvYbgEfMDhwg24sDb9RVv56OOxBs7oR1Ex
XjIU4DvFLm1ny4dAFdxadJ8BasIoNI1XeZpHvdfJxkmaTC9+RsD1aMBAyZfPc4EJ3E4KLFqlV05E
azN/r7lh76/4lwOhUnoBIRqo+uHLM0H/5zXpYtUtMwdn7ir5I2CzoD0DQS/2Kv7cJIuLtSHaQ0HO
V+UXprTRk8f7GEkwlZAfY9b/sQpJtwW3ZGUH8tZBrMi4tzBdvpLC7lv0r/oEplnWyNZMG2F7Rmki
DhkwiL5G59kbmabJ1hdRn6QoJtNj8uDHFruqt9koloaP0fDkJ6upFr5j8Rte+qSPamdW1tCGgpcB
gItDjckGdshEawUre5AuNndkD83z+omOWoqLJrF8CrXjrFKzhAjymLrv1zio7NNRAqjCXp2XlAfs
++2/6qncea7W+X7eCrlJAGmT7IoqRDhKhoZhVm3T/MZRwLxwy/oLM0HBzR/omugojjZpky9ZuGwj
+K0Daj4qiNZvg5lF3c6pRoaE3GkU/o5AjeGZG6lxHVq5VoHp97kbxwQ6Il9FwIykXK7+vx2M2Llm
Cj2I45e4ipq+GYc0aPzjk6a2Z1NAdhFD9gOJPozrLFlBnhK7hEVe2FPFK68sJW1XSyzV5cbZO8Cw
kJ1XrB1vnsh81P+T0+XDm6yYsn4ZE+yWhpMjqL340LcRKqxGM0Wzi7osmvv/ywfestqoeEjserc7
IKQKLeLGQXe2ABRVMLcds+RTfWxt5JP3wUxNV/DfXoCUS/eyktAX7Bzo/5+FTDKvT5nWRemI1Oo3
3s6pAd2kx3BdwbamdRIRtUAeIDhIRoCQWddUkLqIaJfLIyqKzlOlcgYXtAKk4dewTcjSzzFCB6rn
LZ9cb/p46b1yab4ACuShhDDAJBLrzAmTcARn4C6ePCjpr4qkuWR6/8qjLqDiIhLaa5GF8KLQgvsS
QRR3YNbRHJjK1/wvrO+obeIM4em4SSfrPwl2XQiXX5YyArwkq6fqzzZYb30Slijko3fb2FaaIPxl
sPLpr+UXWON4sUuQp+ZQNTBN0jc0Q6fCJ01WBUG/mZcwKFcpl4fh46i6Qn2aShOc7Q94BlbWZEvz
M6NUvZx4PphA/l2g14oBRXPHW23CK9+wKsTOStYbGaLHJ1HkCliqCXluh2FmF5X8Dr0bXZX/akJn
aVXLB8prSR91jhAccO9VipALe1gJOQjVWrDKop7Uh7zYuYyKnNsvHaeoIj8dubzw+AJ0sb4Gh+0x
UzXN6IgNyt+HAHSCBzdVgImItkaJ+SCxeoe9E1TPpDXDZOYFbnZ+Zu2taRzmFMveTjFN/hGF0Dhe
hXYDskX6gWyV+6gK0ouVvWxHmUzMCHb6C+PQEKtG7kf01EGm2HwpQ1tyrkwEWk/4uKoAaDNmi1k9
QJoENK9kGH8yKeJqEGTiVsHG5YQp9T8mJEnouxfcyqE18bs0aNjBGxyG66VEVnL3OETHpLRUQVu7
ZYfPIt23Hws2k5YcH2Zue6jhOp7g1XQbxznlRS6I0JNi7X1CU6gppud6k//+/BO9GRPM6V+TGezR
XG1AH7aiQ8QTCwbgfbtjMHKugWftQ4wd3SNl9CEaCb9F+6PUqLRcF8Ptk1UG2VcvIXmBmU/3ojXt
qcABtmI6mXWhmW5ts3tPgSAkQupWGfX+ww1tqIOcfZYw8EzKjeeNsLFsB0dJogFGbmkJvr7GY3TW
MjQeYGft0pTCIyHmK7ie02f9xaqhuoACUMJHDkWyBclhcMBC1kYCO/FbxSxQeic7YhXpkOiCLzXl
oFKy71d3jWySIQMCgUKxLWXx5hiqM18UvCl7a4n87fJu6we+5OXZCOmrbpqFyMgNYO637vXtcmNA
jHf6yEE855MKACAR8G7KNbH/ekZLwoZU3304D5yst4qqI3iv6cTVDK551IzvKpd8N/fDhJ8Q2oMP
FntFCSprxECVF2+6AKp7Yu4eHoKubPB7PFa9HQZf5i0l/yLjiCv+jgULYxU9gMUGKeTfF1reXPjX
B7swH/v58zow0huejtAwDgztQvEcVWZjPTCiAa7TYgCqGWNsUZchg8f2WcWQC3AOTROej/uLukK9
BvW8R3QO3aGt3dD3TbCQ3YKdG/IBTqx73Vjivh3rIMHe+zf9YEgQ4QUg7WCKnB5COYYhk5XSdDSc
X5TkQYOAVQLnKWVYVqkzunXcJ2by9xT54j6vuY6WNBEcNfWzK1aiygKBLCiy+1A28uFS6lZkXI2w
0Kh4LuA18aA9/wPoXL/3QO9yGMiV7QUBwc9BNLCfOtTOUQw2AAGclnMmbUyiDmnsD7VopYs0izs1
bJT7set7oiQIa2275j86desnbLZ90UIshUB6Zp6yGfkcdRnenxOd/k7R7PqBuJMsLHcMuJ5krhqg
2SBNjIfG2PdiG0zxajqTI+mb+QQvZZdj/K7TQ0hG48A6IOChOSyEf3JynquUSjvfGaJln8HUE8TP
gKLYYqvsJb9rxu/OYXxsk5J/XXW7wO92FSv6IeQHi1wHEjwcIUK3ie0NK9BuUtWocykp/Fq5KIT6
0Hk42FjzPsktLoJUwd0V0Dn8A10F4et2KZsogk4lZr+sRIaLFwPpEWkWgYx7dyO4EKanMlfUkh9b
ec8404ial9OBmYzZlwRpPxFNWzuqj90DnCQnhQ8y+7oiPi5mhCMS8R9I720jFUNJdGMSlZsunckW
OXV9F8/CN2v3sfulAH5iduPwYynhl1Uyei+t7SaJKgVpp7GpH/bPgb6FlPvb+vKzylwaeMiIm3FZ
CVQbsOzQz5BLCjbl/piWE1YPtt5sq2QFcOTJHHQQQXxQLERTb7cLymmoA3A+lpsYr2g8n95sI4i6
qLieJ6ZEX1bdB5StfoqO1eOU3FxaWeUisV9+PdudT+JvTT2mnHoLcU0nj64sZ712Xz9s31KxEFg2
52ohE1W6z0MxIvw9eAcJQQlMJMiH5NxM1Q1S2GaHFzgIGiqOnOfDcVo2Gq7odypD3siY8n4UxUpf
ZRGX5tNuE0Qo4aQCb/7e2v5936682pl92185qBmN7dIjP9SXMsfZOsYb2sQgbAyWgxqXOv6ElHuc
dlUzC424Eddoml1eveNQKMz8TZaVATJF6Lhd62fPR4g3ldaLjXHs1qe6WyuqEL6MHxfs5dgGbMSt
ECnW5h59aAzzs9OO+mf5QjkiS0Emg71tTAt3bpCRhKNvuzjy1YSSV4UCtqVgno0vGTXLzfdN8Se0
/eLbGHQpDJeaY2sNWiXEWGn2ArPPo5Z92G3egR7F4LWOjgC59b2ylZK55exXayvW2Xt/lv9LbSBP
2OhDFx/Doy1oxK/ES8Deil7jfCRe+3zRsMMHeznbvqyrzlgS0G8T5P8CKNxB6EL5XWUidw+c79Y7
WLQDY+RXdkDb0/Kmfu0hzkdix3HYcnmM1xPwi+0xUVVhbF33DvUr+hfjbgs7YuucVZ1ni0DvMqiD
Amog5HCKZOb6XrzDNsCUIpSR+i1g5IeqlWrm+m8GUWWh6ufDt1bCkMawLJM7SU4Xxv6BjTBOJ05k
Yy9t1HQcf8UqWuKBqp/JK6BTguRmUEKJ7fSwSY8SuUTfocPZo9PUsjQ9GsSPxYNKSi/TaWagxu7K
XVxXHWxo/TLVJ2t6zXFnJcV4ZNds4D6S+XyT8bdLRRV/3+FnNnWdG1HkvkFB/OLFaWz5R/2+9ke7
dLTtPWJ5ocua5Ebr786Uv3hVQ9DbuugSwtuv8Q0vWH0YkowSyt/f6d4q4DvSgP0W9c3lipXMyccH
dWehH1HDgdWcS3kuKbsr692bCc3DPOL45Paq6ImBN+9RLA0EBWf2izamI5h1Qwan4lm2Hl9jd40o
/5K7ykpwfZqcEt1ODKVma8Dx0LizaaVFskIspYv17P48FVhZXBocikciYsQ7ctxDpgXVBF0U6poA
5GA/jwFjRjmdCW3BMT40fGxuA+PbQ9K4GQ4nLJ/DF3mRv4VgW56Q6JdAfy2ZGIeN1eiEymMMfsRV
DNcAZOj6ZOQOljVVsIl7Hk3NKAOzGhtqyXHAMvWJxBYU1xgF2xYoB9dEAXb2xvldWa1oFbeQozEo
zdoKdYfPVaOjKjv5uRjvjyE592qgCI7VwYAs3xw5bggT+n7RnyJArQhiHFTst3B5QYNWnHEeyG+c
SPvIMTXQOj6J+ol2eqjjYidAa0ivxSFbxWhVrRMR5k0DUCOFuqbVYxZWpI3X347c1MEOhADT7QyT
nOxarf5jbriYTA+76XUEMHSzG1Dh+9ZJFg6JCEC7pIlJNxIaBP8OxxZYn1W2IUQJyGmH16SC0OEs
cdV60r+SEsocjJkKVTdKUBOc82Lve3ojcF3FbRBamaKmC0VdKpIJ4XK0FarMZWTisGHjcQvwj8+j
jm1tpauvloeexRdWIwB7CpSoxEDZiykg2WRVO4S5+TqHjkILsj6sSWPqCZDenMsmhbF+usJPrAX+
Kw+fnDjjk77Gk1MURgcgxeIGUah7gEeCPNDI/Nv1Aq6hylHyAZaQ3ZVutUjZXxwsKXLLCJaOz5LI
n5O8gioj2NxfmBztkqq56x7zhx4469Vvg9frjQfxGS+HdnoCKlblRqlm1q08BJfx5HZ4FCh20Xzl
QYbts7NB/bh6c+RaLYBu42T0vK1KiazYh5UmmXtV8RIID44sEL7maxHfI9Q7rJiS1YhDWh2sbMkW
54XooV46SglKAMf5z8tEoK4KijFs88dx+cHu5LzH8Vwo8OTEHkqkIvOfGA7c3++7jMA7smt6Hkcx
gVdBx4iCGH74ZmSGZ1iKQxokTpaq6F9FM660aW9rTS5R3lJ8wNBgLweGn1TCHmdFwMqR2EMs1Da6
1F8kBD/iXVoTUiMFOX9C0DRQubMycJan9io/pW83bx7a6zNLUDo7A+pEIoPiVBmbJQJ3jwcQ8VJ3
aAgsgkzFx+BK9VRojVUugQJDiG5NskOf7LrM7NS3QnecNhtKunwsucKxjxkYRTPGkeL4douyFttP
ARz1qs2SWLvQUcK94+kpDI/2HA/wDau3MFfCloCmneGne9ODxWawACNYMnGA5UV+IpPBELn+wrrJ
rGO2ktpuLDk8HyZU+sHIHNxkFZzyaeJDzy7ULpPHYt5RUjwP4Ej5mxosJdr3pG07Dk6z2kkNF4aB
F6SYXB8T5ZF0qlUYoccIerWpHA3j3X2Z38rmDgBnCh8nlnjC+33Y2eufdpAO+j+PziO+AvD7rOEV
60hCNZc7cEGrVXQ+5sAIk2qwh0zjH56FdeY2Rul46cWNXfOpciez1xSavXjK4ZjPeP7+1/cc2vnv
hfb5xKTZcutKXZ+d5cCZVuLWp6ggz+V3dD0xDMpoSXJ4NXI+fFvxpwZfnYYbggZlEfWKIo/Wwf94
esHn9H5sgVpZj71vJF6HDdEnQHm0jLqEG/sZ3sIJVnPD7LWxcfRPGqKRpJtaO/vSSFDjDslCfZul
w6Yje/49XMyEwgv4IsZdmC/Z9PmW0DYmNcwctdzeTdyoLoWIZFW5PKq+Kjt2b7Og30JRANkgxdQY
vwSkghl2j66kIMPuwvkBlURJyXY0PmrcqVDgcc6MfsU7JelsIMXscXlTlVYk1s7IH0FJOa2QEBxo
YpDpzSgRB4orasIrNU1T6lA6Xpu3J1vvDsuNafMR/Khhk5m/oK9880zXdk2NDgWl/d79JsSbW6si
cf89MTdyfvoa6Gsfi+yYzQRWlHZRFJEDbmhL6sKmHxtaryP15xt44WFQ4rhy8rHPyUnBkopt+iL4
rRfkIipVa0yMGGdWfMWJOdHMFrrX2s2k/3QfhrBifHS2jX19/lE25iGqYidXhfZMmvD2Mi58JjZx
FuvbygVXQjcz7BcoB9h8ISkqun7jpiN2k9Z79PnxK0Sa2BTSbTA1+02ns0JDC6hmceSa6egT1YcS
ScHdJdjgHVk9dCGq/HFVh+VRdGOqL+x+5rFnaijk2mx45KO7gYWaT5YxRqDwlTof5W9OS2ipWTUf
bki1e1rshTED1EBZLnSGjviaNerpZ9U157NzVDpUbVVvaahTD41c4rJqF3vw13o6LqZ0NV6iNQyZ
oLaGbqjkoxmLdunqLcYHmV3SVISodWcOm/zI4+BdcU/7zNcnbs96JONJKbNXXPdtzyDHxNt6u9g+
FYrHvtMOeIkSarH7lnDYNhC7rJDzC5rYHBe4GjXXaOHPFdNXgORy3Ep/t4hdhdhCjolslDQGYuoo
6ze1ioNnAt8IpGtYrkP7Feex6tN1ySJakJboFR6M6msIH2CrEYWFWwY4hri5ppBXm2TlYQTTAWu9
OMUmd/tzzMr/pUKq67QfsUq4YvBOfs5O4wkOGH1F161+IIvFbHHgA4luvpK7aE21lVLZFZzoXc/Y
5nSxjYslc/2vYD3MJ2TEEPm+7LDuyu9D/XdDFPKiZLoQRA3eLH86/eT8Bsj4L5D4FXP7ILYo8VsL
dNti4S5qWKfnTlPE92nJLCExgzznjLT16fvVHNDTeiffwX5ZcwR8MSDo+a/DNgotDvT0VLODke4k
bah8mro0gjNPL/vYUlvBYa4Nubud/x3xQmY+q2BLf5MzsGCmN9b0cbI05Xovp64iqDeyhDAbHIhr
wpYlTDeaaV3I2ItwteCqimplSPpqQnekwSZ0jBq+Kc3vB8B6x3Q+TWUNoamgh8ufISN+yYjOEguz
cwaCxAq6wGC0JKs/xJzL8EGQqch6fyryJX9UxdQi67PWNAe9HVGNYJDg4sGyJC49ZaqYZaEq2Ots
D44TNoWBHnJIQVqYG+RsKz3ccaHpf+zAb2B9ZKf7kav9MjoYhJiUb1Cx5198SrOQe1/s/IKwCtnm
Io0O471gs6ickQGghgFmXEPKx4UV5v+rrJCv+R4EE9VgsIr+pNR8SpEJcNf1C7KeClHIa2CAaQwh
KNHBALO/wuVKZxt8RUptYHQk6mXZEO8ENIdpRSKD8R3NQjhgtuRyxMnEfTAjbyLpqDZ0vxy7KY66
CMhyVE9D8Aazemu+JR+4yemXM78+19RLgiHDAG4c1bTBzk5FzLuGs16b6LJeapIECi55p1poqPpS
6lTBgJoWjmwO1mHsAijs+afkEAJWtO/YxoFQTu0vwQiE+74rnZq6nQ8zILuBgroCPhPHd7RBTlCc
66+wkGFL+x26MxV5krrfUz/KTFJOXQjUyTrY7cNEKjrrwPSL7EyLTxo/ZO0x4yY28DhuWvZ660HA
EDg1aA9xUJIhX0mcB3PFPim/151INQ2QJSXlZ+1u7wKCoFuwKNxtIg6y+tB+s6VluiCY9Zl3wfoi
zn6OLmKH4PXvetTsuR5PJEsPnJICBDQPeKYzoZUWUiDzJRkMyMVWXp07a2XAkd3YXEwZGA/A5GuU
anYHvFznl/UZvWPdOJf3atfCaItLpHHM4NS2ytrY0L/yWMhBeZOJ7GiTJolE+n+87OC4KB+41/pE
xk3zl8n1+9JEef6tqcqiU29osvof3rTZwQoHnLQNA1vLt/aO5wMqbtQ4LMWYn/h4JOkBXBWlPBmu
7ve4wR39D4olUiDuwH8oySHe1H5OV4/jvh8LRBuY4lVveQhey79e4taGIcVDn8AFBPsUVVmwppj0
8N0D4pQAfuJt6zN3eE4ai9pfaHBOJKle8fqnLFw9mLIrMndwOUoq7NelV3qpzWZLOqlqQceNVF/J
796lznqY9F27hPeZ1EprsP4VJTkpTpgmTcFuiVI2WKIwxzTCxyWlfgi/qD9sEYbxjbauDuIv4d8E
+SQ801aCuusiNQdEvsU7Vy18/1RTSy+EWCRAAZAxFHrGXoqf4XeNN7fm77qdU8prMIoMl0g7ELgp
+EKk9bj2u4qnHRI3lL+cZxJ4AqAzLORMIPJYzA/TkWzihSa0FNI40CewMwlDjJwmMLvHZkPaE0Tx
8cASdKYaCLaYO/45cSOkUb4dHLnjAjlLtBx/8yQ2OICe2FnTceb+y2hKc5CNejysp9U4qzUggqXZ
dVqoJ/AhZWMXOF7BJg/P/AX+3j90tovkXIvYNr9kpw1PV0CcOfeKoQy5YDtp5xHvpB/lrGzqzCqR
2IM94T5B0DPXv4kj8DLfwd8WoaPLRw8DJ/pGZ4AnQJ8t228OOvMTVX+ye/R6BmZzeexIjnO+7swy
VaGPbMlO79st44cGhZt1eh7SUlkqxnPYQzkyuUccy90GJiBKHpxzcVFz10zo9JFd2veKL57K+vG4
o62JPyfv2DKrGj1CBna2FAWciJGLUvGjt9OIIo2KlicGwYekr3Su3IdE69+LJNWuoXu+4m/Y+oQq
Z6oK4yr5N70kCH6EagliE63/uFrTwlxaJtUAn1M6gRAYiqDZ7GMPFuW+iBm5KZ9yH1bKyMNgdgT0
XP9nbtMtjVcuFkmQ9kV1ikmjHIXiRzL/1tdqqodBW6ex+pMIfaxvdKHxYb0iQU85LEbE/4WsuUNP
nPaqtZmY6a83VdN4rdLtUeqzop8XdDT93ZXTsbI6ZbV2LNzOLoGIBbpQbEzyrI+AOP8iHkFuKEcy
vWZIgMsPOGKPdICqsuR1ILzoO3D0h2pFJOYktgdzixsf9Ti/LAMO1bkqh8cK6Vi/mcFmLMTiJWfU
qgbV2wgs+OBvt1Wk8lWt1l3j7QV7ngLiWtghcU+X+l+QsZUguyonKoDY++u9jWqmu/nRyM9xeRUD
q472wvQnlk+0HuABb18JXkLC09mDVwDA2RuylpJd+uHBF9aj/Evqub+YFe2HR5GGY7pAAFBpHZCB
gf9oLXsaJDaZAkPR9wU3Q5bn8S3WdgfuSJ5EKNazFPjbPtZu5m5Rs3WTHtBFXOgPyRwfBlrHLqMD
2w76EMfR2yxGrYBw5e+pBOEpjVSP5Dvw6P1skb0xXu87tosnLc7BItAK1rUyZXlntNH2mCNXBC0U
ZMEw8x/65T5uQTuJv5jcSmORmmJnUa0bZRhOZWesU3XFUFATMWtPo6xse45VEeCAdcpccthWVa23
AnY3hJkelhpUFurT+eHP1i/7WOv2VVTtMe6k9LWaSdcqFPNQ73mBqYbwNBx83j+33rYut2KcClbE
tzFbtMe/ftjUAA3RqAUpc8H4yAdnBgPo3Kkij7DkDmXkbc3hECEbp1ViM9xv2F2dFL/q/fkMsoKw
6WGKEKERGQHq3X1CjnMEzggImTtJV4yB/4QmgbJa/TGesEDY0B/OfrTnPfd/sKKQ/GuDAv6huIg4
J7tDAK/IL8g4Xx0lJsITXKPMAIDAARwI6aCuy/J8p3VuUCuYgrKjl9Z3+pMIWJ8EFC9yKXHLjDer
xjcjXfxThu/OVoeI84N2Kil0NF5kLq0mpx4xl1CwZbBbNic0JYAvNJtrdG14Q1i+ktiMsrCzwbMs
m7Y/S/rdQXWIp9veOAyPfcDL2twjX/aAr7ecpkqU2PvVaN8vx4NAkK8tY/qg8isUR7yKZyBgjDwb
J8X8pz3fLGNuiSokFzTIINXZIMmUPpCyWvxgJo+o8tfktzN6ukNyOJ6a2qGc+8MAV1W7dGplyEob
A2JcvrM7IzescmMSWWcVcMjdB5RVRBrIR/xx1CmuoxSpMenuf3M7je1VOoopkG88WRbWY8PXNhGQ
7usrfao84ZLazh6FPOyon/knTgo20HXAnhGLxCVxeOlxBUD0Zfog5S2GAQ5bMo/ZvHTH+w7IUsRm
p+Ush3xc5FsjWc3t9WvcbcYqbww6sNjZhT6d/H7YoxRbCgfR/0muIRRYauYvSJV5XMX0DzFmo5qd
0EfthcIC+ObK6tmml/2nfXxd8JyeNDJx71koGuUL/BKB5RNet5dbjFi3umG/oNVSvq+Gq5X7iimz
DIVLGDkHj0lnwG7oyaBun6Ldrh/8yZrqRILdD4laiFHdhwobG8b69z4FjyDQZFOINlcQbUSF2D69
LPJknUqJa1HAH6eKvuUb7ioZv5OchyA6N8VuapwNSKKNsg07Hh81fow464xn0Kdduq0uvMujknVA
c/6w2vmIhBB5MWaWPYeRdysS1Hbi+st3GZp+1UNkuE23myrtadsF/TJBE6bOHYGYzBMHLWQ6ruTu
G2xPYayee6ck4Yo2E5LT6eFqiHAHpl7JUju84y9hhs2z0s5t3RQyUAkQdr9oHZTRNxnNFaP83qFj
B13ByT4xiXcDl4qGE4vsx+1tsK1cmK6tEC8aVXxEAAs/r6SrpxdsoGAPvgURKhIJckmiBZgCqDFb
Vhe3Jf0jzamqTPeDm+otBJsvVKqNcUKwUPwWjEBPcpo+5jcZxEuNfLS/THdq8p1JgplIp/qmX9Oz
m40xw9vz480Qtfv566WbThEsNRTG8FH7ptlLH1Jv6I2bCmqISgRndw0me8nE+RplYwka8Tf6ACGj
luOCGRnnZ0gxEKpX9DqLAGlYtLPjnAbZxHozsXZNsem5HgyVhtNmfSFQ3e2T3tTA5UpiKzZC9gAQ
/Gla3SbMl5+Bezs+pAxxG1pNHqbMN5Nv6My+JDIpRdm5imcyB3Pc7r8B2aeO+XRtkvcKQEFvKObo
X9SJ5FrewkX7vry3XUBKHsvVjnEbyT3GROmeXxLmE8HoUTBAJ1bSn4cHmr0PrwGOpZqQ+S73onke
2heF10jtGCANo8CxhgXGxvqig3iT6uwmU3JEXAw4aFmRUidoO2wrTOFVLoQv3yFQu+ZWHrQBdvxY
7MkODJjFS0ufRr9Kw8eJ1a7iNDB9yue3zsnxRshsklqVSzrf4b8B5VDLzdZ2/mxQ2esitW6IcjMt
xmvLkz/S62fKjvn0PnWIEgbXK2TSydrgHh/EQsKNCrZ4Wjqxw5GCBFZy1yCJdgrM8wiY/Bdx9ROd
gv+usSBrFvk7i3RLjTsZNSH6cXToIJTmDA+uAn3OCSbsCnNK+sn13qH/Lvb+imZekZXzNKYemS/+
SeYmC8LPtvg7cyEFK8Zc+OtUEAN+uSciwbssNB4UKHQISJRvQTARH2bP6TZ8l7enBK2ShW4+rusR
i2YTUHTQ+0sptZZg0GBxPNyMhWSQi07MKLApilUWb4RQWDWfi2PypaLOdy3/7YpE+yuWdE+7DLso
RM75nKfgH006rzAxvYcPZjTmztRGIDUtKAEYrikmntO1nE4JrWd/CaYKVXcLv1HRbPXL1DLn8UJB
sXp7Uzc2Z1v4k7D3CIi4nfCZE2kWcnJebRKG+4kR2nCSYNntHOob90LBOWXm0oArLWH2kDwStGsu
hYRKAtVzh2v/PBU6v4X9e6BSrI8SFGxZq1wNUgDKa5FBorJdSY0CwE3JfEHkU7a5EVW4H9jfndJT
Huw2Mv2Qp0AT31R+HnR2biKKUB1CSMrCX/cYdTlNhpkTK/3N1x+YEynATlfw6QBrhkWMtMWrqlj5
i3L2Mg0dDyJU1p1I9BNJH0tNRkraJ5XywYCMbyzSvOUXBMHaqDGgMb7lbDQyxsW9FKyaFtWUouaq
8KQ3U9Y3XLz36CSrs1ul4vqmBABn938IyYVrApYL5rBNV7bupBd60Cq5QeARtf5wXJF0a8gBInYF
2/H2Vk+EBzlGXfd8cgNaidrRBzmkmmuxfvS/FaYp+azt8bZa9cs72QxPwFO/4KRo9ptx3lewojYE
BWJ9bgu4pdxASOF0JVyIYq+68vbe0MDpHcKWvm58sjE+/63cd/7SBnObBAzk31NYqRQUdYRmtz7d
ELeoJxgjw26A4JIWUterdXKGSluhkAiFCjfRLBprfVyvulCbW6q1e7Mfgma5MUUN4KVRUeWFWvP0
KZIf8BRYsU+CxcT2Ry7a59/TIHuS5FhdhRhcWiB6lShC9aCKBLlNf1rCW2CReuD8RYjy2q/r+XD3
kna48VhF/FyKI9cpsC1PUTb9QP6BqPoa+ARACGwPBRaLq58peaPbGqbH18RXIopCdDK3RBx1yk0s
87Mel0jP05UyXgFi+tZ+utGUFzaQEMWeV4fzwtODOg9HT2nw/ojEhpWD8TYFox0VBIgzNCX9o0U1
0U9Hhj3q8YxX8iz/DJhR3XJNfimNwlnufnqYIc8Pvu9Wy6uX+0fRX6+f82m3ZVkm/hlldCDwaAzx
1pM1Y+G9z7SB1faUnXngXfnubVgs5CsnAY5N8PeegubMaq6gPytUusI1xDWl6XbWq9AaC9MQV8t1
5BIyhj3uUdaUV72wIRSdC7CbxX8sguPJyLsGL9QpkjQJedkNGXmAKO7mpd0ml+wtXjJJ0yjdHwAC
zhErKTQ6iRUR66WzVYs05AC7qigyw08NMWivOIBt5wsqmAJehjNCAt9DNkLsPOdNAbmGXWbnrlX8
IVc3vcmDKC/p1uXEBBYLwEjQO5GlreLgbKA94xv034RozhOsmA+McgscjLhJTUgnASMO8gJfpDYi
XvPMrM/wLngbqeQvBl1oofWDGAVTD/gPf/oWs2iiH5WXY0jbJhkBxqxIeHp5wu+EmU3AzuzKF3m+
fJSOapKHL6Sr+P5ZeSVkc+dhVq4cjehjeldMhgdEehsXN0QrG2ceOdCG2eo/Oah225RP0Sn0clqR
er+R9Cb/trUEwNlS1OFHm43kuc0Ge+7xQ12xhzMw38ipO0rxrCw3rERAhUiX1VqQ5zlaBheNmDub
OM1nSkevwaqfVJT5HU52NccnR0oQGU6CKjxtn99J5mulfCmuSwl6ytnxdWsAW32eNnJLTkcVnynm
mgL9Wi7lYrUMlo9zfUkO5NIQaJm9RCLkQBGQJnJ+roOrEB6Tpbc18yvpFwfKYdmMJ1DeFBqiGc3+
F9ZtQpI1MeRnE0yITMqbfkr2DUSqLX/obtxMnyE+0awWdQXqQiMkdyCIZu2Ve2kzuxRMVjZeHQ0l
6iEOIUNKMYNf8QL6o8Yc1p14MGEkhGFC0MVrABX1Ouy5zWpPZB33Z8uMYbO7Gub1nWq+EW4K8bUs
qLzWwFR62qNWwiyVauKboSc7E0vPLuMaNEEdxExfhBkz5MJwlg6vxOgm2E0KFQk8Q88EFbhDId63
aH7rMxRnEacu4k0u/w2CM4si76RFNqI44LmRgFWeSKx0zIY0V4W28z1c+WcOCkMgfsAgaqaW+UFu
SqxqQVXRLxMnlA0/Qk0NySeWxTLyez40LyV/AWtDbeTee5Jdee/Rcg1yPST4xeeNPFTjc6kx1/KR
ybDWSqSOuQ3EO6ObFBPmcKIHd/NlAigJAbOcwTrBNBZ/6Eq3/lQDekQvDKjmqBGBwud5yLSokndx
pzor8kzTKpgy5b2BW1NN569V3QuVIqmyRakhjU/dJJXRExQ7BbazgOVxod+b3z59XxGFNoQqx0XM
ZkJKMkblorTi2Gy5UmaDTIoH0SA0V5yOe4roVxaD18MV/dTBs9rMrnRMcMFTRpWQNGCiSlyJjI7V
mRvp3fbex29z3pvfJYPjtxR95tcrZJPm9pJSTtjUNA9QPQQMGxXpVswAHLEUvAe1arvSft2vQnAX
2Hz0MnLHf8cAsQMPcbyqJayXMsGH0NUJu3nDVtwRJYd1wtNB/zr9pU3xqtuIMSEfTacHyQjHXvvm
sBF9IS/s1W4PyB5uJ6nWJoit7tpWd1ZKS7mmGPxb8KIVPIbRfr8d4R/NkXbvpGQAm+jc1Vm7IFln
oSj3Qt8LnHmvU1Q41zlLBh5Y+p8EBvQ70Aw68nbBjhKHncxYfcMOpu2Yz7DPZHixnRlj0rNney0z
JFfrwsmr/B45DzBXn6uWCgGpaT+vDKb+IYkWlMnnf5AfNIPPjajrk8jnGXUU5m0pe+WPlrzFtEVU
JvGg/IAYYAcMlE6NC4ukU2d/q5slJZMtB5E/QjvLICurw1MiUp2OC6OXvriKltriI/Lw8p0omr0w
6wJjxtSEQYrJIDzaS+mGu+x3ulHO0iniUOKt4fPeWE0M2LtQJxrVQvYPznXW04636GvOhzbPDtSG
ydW1Pz5hd5Oz9wr3dm8TVh1ml5iDT7FYNxHwlvM9LKgE4NlFgZm1uF25psVcuFYKew5WLgt0KZqa
ZWJc35D/VhG9YjSHZRiTEcFVwOZQcdHNQJncpinoIDfAN0PEfWTvGJ9JetbNBBobNiCNPziFN5jL
TwnLuN/uJ2PFFiJ/V2WK3mg3hjo0VlSodoNtLlqH/p8/51XFNwjKkLGLhnnQketFWu4jqqNDfeuC
qTcHmLux+8zp58+bPBbwP40VrJIDkbgO2e4bJkJu09IvWP71qY7lg83OdDqkx3PakVtr9ji1lI/5
AvXEGq0GEbuX0Ws+STEZp3YQKTuvK6fcoOQ2lh3F0As8rUlHGTmUnVZZIXsWk4yB3WPoNNmhKhc8
Ma3EeApUl5ZjndpWypCtSCUn+zxk4oVZz4BpVDmc1iN3DxoqcgTyeshH7ekfdnYJ8ZI8phKnZd3N
6Y2HhXW1Fn8fvhg4AKyfJ+3iyELkqg4MiVp/ZxbLMuVJsh9A6VCYRQG/OsNfCh0gXFnj+ZpJFtE2
iBw75lygO97JsD7Vq4BsNsZGFqlfWJPw0Tw4TuOEh2HlEb3SZw7o9N+NBvcpVMi/QovDs7S84T0F
IGiBUXeTsjXFQWvVMkNO7wjQMThd4Sva3UiLWSN96muNbnkVzFFE+Q8rxHDcwP5QjWbNzrIXUc8n
BBOjAIzoz26P+Be44L3FTOlrDT1m1uPvllnUnrytQl8PQd6C3ucbctwk2n+mMChWirjQvKHYvMky
gWkpL7yQ7BoMpFdSs+jU2H3jecqoj+W1Jk1dDbhbnvYhd41EBf+EFI5x2vLBaHopl3wBx0fZmbfl
VCNrh53BYgaa+KKWlFsP/4pxqzR5zes2xE1KlbuaQeNaeNLxOPO9b4ikmit3GeooeelHmicRfypj
riSH+/JDClyo5I6qDNkiaBNwa+vtnsUiI/X10QNZKKBC28WAzHejpZiYM3Szyy7K2vdwcrzIEYvK
0AhmLAGWBkcB26QGETCEWUXxmXk6A6SiwarK0ItRZ7/JbOuWApio/1Z5QFI6lBmbYnBCub5N8gdD
jCNfQPoiRJ0dX70hqSiue3OOw/DYUGo63gSDD5AlpW5ldRVtZkXN/nsAePYYhAsJBBv71JXJk9lu
HqlvWJdhLwvX4jGZ5HeXd55XG5pgXtLiyRsYHsf3lIz3tzd1Kew4ZmjLlQ8TgmJePHgLV7e55jrX
mbJm29zAlNLEsFUFUvo6ukNd+Wj1uFQshMgT8Sch/+m3QD+oihpY2wMnA9jRGv0XCdxDDS76VFfn
f82c4sBbHdtyKQohwe3Dms1f9eSccJW+YitJQTcvXplJHtx/BrZey8swVVgR/Ymtp7RAktVPXsML
FWGabhM3wzOv1g5yofrSjxGEKQHHjUJV+FeWJTUF/I7rIDBW2XILnxjQqSECefx16UnlD5Gm2Eqw
3+xzYtVWdrX0ydd/OT5z4qw2CMwAZpP+1vsHByql/eZOq3Amb81oql3pZe5pitUeqauVers3giBL
1C4EiX9IHlYkTMLb7FCpDwGl+TpzFamfbif/3rJjoDQ/1VV/GvSLy7cRoG0fHNs1NBfAjBj3Ri25
LocPjXpbJCXwcu3lfPC/EOpa98VD9MEciri92o7AHJ3Ig+M89tKhTMCL2wcCCuDeQ2g/kcEk0XlY
mHsq81XX+88mWcXgAjrbBt7UZNu2sXYUGhOWNRqBqT1gV8xx73oNcg91Z/tF+rRySU4HnMHLiyV0
IXk3oLXB9GI/Ify3bgBoDP2NZfElNpEGVdMpOnS8+D5mJmiHCQPg2vXyLUKA6ZxNawQG9L4wcQpF
kukAy+AJXM7F9GE0oDljFfUnkScjs713MwPm/jObkn+BjTSVXGKDGgvGzOAl4FsYxD/Uzibx8JoZ
UA8TfUeMOueNxoiKeoRvUAHzvEHc2jL1U8ancb1S4/MIftx2sD9Pr4pWYvtOHH2dT/FPmCB6In+3
CdmT2zK6LWa22CpZEVK/2exe7O3pLv1nqYWMy6gfCkfGpeR20IgOCPjiYh4cPLV8rvKnMeCtkWtn
R0XktYXPOjIkLdLqHjRatOgqLCSHm/hR0Mpu4OHKxon+sbvgRYt/7MkMoD6Ki28R0POSaho0Zggz
Ceqnx+ZrR9ymC+n+uBCXoYc4O5Lhaap6tFRp7qar6NnY9wSewuAWXJklxiwUmwG9HxHTbYwr9bY0
rp5Bmh01AjrVTyxMVP/mIPdz7hSO5hKewiQtqkk1g9u2GVR3UIm18qV9q7SWPSDlb+yjFVAC3nqR
a7gvptC9RvyaBAsPudABdVcVGGD5JdsFwevbwM9wWpIoMAX9bv/ge/5GpKUnT7Czx/FHh3+fIiD6
ZrGbZnSSNORQYCvhGNfDD5iETz/OlVz1H8xdyyTiIL4VW1hn75DlYOSrxAERrx3KAZlZHhaobh/K
rYxue2vrD8SyZ29vYazzqfPgOAxHlDpxEtxiA+XurD1CgIySAFQou4qdjzocw4n2JWHMCW7yoyR6
OZM2fS0uH5Xkl4LkrKTH2+HGLObG7v64U2yhBYX0YJG/H71GpAaN/tZ2c6cYuiql/mN6gfjaNlIf
+8wES1SGXBzqerdptGk9QNBnpC6sShR8QnnYz5YARzoE9WJ3mO7k/TrmjudG1HGSU3Tb3KtjiV+Q
z/CIl/545JODVf2+G+SdBi/hs4Mx8Uc+kra7ZpeSUQsq5qbSDjTJISqZKSkCgxwiOoZvWXKz/xZt
eNrbYEMWdsMVtI3Q2/zUmn4wWLDJiQn8f5BzBgtK+l/JU3ulW4oPkCXXtsVcluvPumN4EYdEzl89
2zhqDWdvmlxHCA6mhdH4CzcLgbQraee5rRqbee8y+VZF8OsSlgQjyOadtpHNIeEG/sluKe6MeDYC
+2sv5rpSiwrbY9ldjq7X97ZdbR7KI5gx+47GOKuk7F7Cvs3A2Fik0ZJxP0O/+vJVnPhp9KsdEjpc
SUbJKC00vygPpxMw2zVJW7pK5fs0it5T8iZ8Xl2O/nVR30mGRJkHb3LxsCDYxlSg4dpdUyjneVU2
R1ZKdbb1EAxmXPUrvrBj1T8H50kKLhs/mRJsCrZiR5Ouk0bGTnMfYGJHVyvN/pD+xXF1ss3ktYOx
C2PJR/5Th6eerKcs7nYvSDxy8Z1+Fffoi9uLFkGWxYDEHMa/CO/xch/lBlH4fje85UuqLkHwijRZ
f5odSjAzTWkuUDG8XDGuEoUvT+8XygiCY4lLMjv4GSqBMcvCtXF9FAtsjHgHAQ2tiYQzERaIVZVr
27KPK75gO4JVzAMSnFEKI6r/HxH8HWEO7Bio3CTZlMNddX2ZqLuvRApIbj+af5VBuBmuQmlln2qj
g42VAyawnGYrnPyWCQoWAx7NnQVzuGzOzBNn/KRwre7ig4UtM5Jj/eoasZDYaHeBVJpPcrX79GxT
WPqECJs2m+EYsdReliiSFcJbpO4kN1r0nUKr2RlfURtU2d4qKX4JIzmxthBJQBg4qmpPoTqXB8X7
vQ00pCWCJbp5GCd0cuX4JUst1SAK3DDgGRiID9ACAn7+1STZGJx1Z+wI1aaX7/fQyv2NGPaApDcG
DTwXIJC6voi3MdX2aG83bH4n4PBbmR+I8KM+98wC1P8l7sB4kyLcZgz6HoPDk2GMNLAcN5fvXO1Q
U17idYOX8RKKUs+QkRlqkCNhRKn+NsRSXTMOUvUAZkdqodNmMO+x4C7gAy2MLwLhVZ3YHk/8fVtd
Cy3IZQ+TJ/50NofBkDGJMZJBHdyFOGQn6MIwWLRjVZScNWXVNthXPSP9QF5X2Pe2CP0K2CnfnSaP
nDNKJSaw+SWugTrsE5Yu3kdbIpTMiYfF6aRFslrWysmRnMToj08GqEPFGHoBk+LWu7JiOYGlUdIt
yIMNrAwSfnLyGS8yT6YNBwBO2EiKd+Q6yfGYTKfwLgUcUnXMFqZY5eABmFWcYVb82YoeQQY+XAz9
oq50yxEGfotsUjgzAFrfPn37vk0i8DiWTob6Fv5vJh2UtiwWmq2q+GbnnTSsBiU+Z3zpifyEy1bc
i3CGv6YyWC55kYtW2MdpugRvIMgDnG6IqodgT9XPrcLeqBrsLuvHH89Dx6yY5caquVLKBDhQjg3g
Ed61yp1plYp2bNFf0FsDYuYJe1yMIP22WxhNHvwQNFJFeaTrCLpjAb0n6ev/cMK6CRoLn/AVRCgh
bxJNlOlHsbCGjB1Pvg4Bp5gxxMbcTEXG+aIip+Oi18c7B+qsQ70d77wq2XM1zXEplywGf0U3GibF
Gkfv8l8kUQh1E8kj0tWUGlibNj7DxLIsZ6JKgxbSPPcSQgaM6tVP5rRag2XFyrVMU8DsAS+UJnnN
yKAVs5XQ5RLq3ibQzxiAKtsFRMk+TIJIxtd2gAVAvOmgAu2rSdfhQeffMaOd+jamvP23Lf+E1FkE
RbmMnoXBQGyroSNL85QpwSNuE+lHtsSrv76NTLPwJV324disG8PlokmEjtW24GkjMjfnI7jZnXvT
1E6AoI4CM5M4IMTv41z3PBlMji9ri923tck+Mt6ero/9YfTP8F0kQiQgb4oxiUDNf3vxjkMCRBze
e3vrFpAZUYAnnK8MCd/2yHT5emj/kTofYmmO8GlodEulEArmFZMJXQx0GvOY+m7KW60xPdS+mrKq
9ol3SjBQ08vsyQR2SdiOVWg1wRFw/trJFAW7+PTKKZgHV1aiWIVDNqnMSbdDkWECN3F/e3rhWjH1
yy0efqetMXmFtcdMDmuVBhSySvSUH9lb4LSsQPFy00ZjL7+b/NJJLaqFJBvoyd/0Yk0rGP0HyFNm
/TS7RfB/iWY+9niZdeOfAys3VpXoFTHeBVR+GizVqGTZ9vbGIeeJRSrHFEuOkSuRtRtuWBmfnn/Z
ySqUhORsQ+icpWRYAaqt/KExhZfK4s5tZf/oB+j2E8PBNSFh8WvkPNh7UOe5QYXR/+ZnILZ3XbjB
ppnNd0esK9PtyBZlVerxK9Q4W34NvRAcHawmxQNEV9VQNbc5MbK/eXC/d4vPVIs7r7WuPJNeh3gq
fBh/Rr+NhFVLiANprJ5cCg7L/XpG9BL8HEtZcJRMHonxWqhpWaJExFfU9ml4WKDa36cnBVDnqVK0
SQgTpeuoPW053rtuQrtXeBpPD5/M88qXZMfRenTK1rKkPiVflTTDYPtodXwlFk+jTS3tvTjDJ1hk
8HdCryxgW1mCcwkk8ewir+vCeFricL5kLg6mogM9MdRDGjf2OCFJoUxRarwlYIV0+sVq/kvmB093
atK/zaSRO3lJ134O6v6quS9fhbePegCq0qmTF0su/qMhJDGhuoZfi8IZwWx4CbeyuoF6RO6O+H5j
LGIt4SWRX0s8yJw2esg9XDks/IdsBA9W9xU8XVnnrRI8KeMbMTMD+5r4kkAoCfhp3ze60qz1GD+K
jStv3zmqnysNYRlD6FDjmegcrGtKo3d4/3IERZU9sKG6ItDPlnpireC9fjA8qd8uZV6YmO9uMnlK
5sj52ItQQkhOCD7RYe0insxrNyADMQJL/D4vCNkh3BJ0EE30XuSY8cmO+s+ti4TP3KD88ywmshOF
DObVn7I0f7Pr3uctwlOP73C1NcWJrjO16HJ2nGPSl0UxMOM26zheF/2WpeRJRIHcEZ1SBfJ9H3En
1zyGDmEcbQtl/5HZ2a7O4A5deGPWuINlozTT0GkzoIsL27rXr6luO7krlEwfpaVL4l1dQ4brOTLS
Ir7URpQJLMy+IjoZ+27rMeKWBHiU+hRPWTC2oRkqilZuBcIIlLDbW/5rsH+KkxHaURYQI6533cvL
0ChR1i11QMEbZrDPnF6WNc3dUQNhFpbnRGKIXxM9B4477/Qg0JvQv/HsnhiyYvg+M2ocirDG1+wD
hZjyZjIhaeIaPJWF6Gq3taQ6YEnm/fvjIj7vjfjMhRpx60692CBD6NdjvRBmjeznK3JY94KY0MFE
I/pSV+CMGUcOyNZkshQFjPjfe5dOTVpNWnSDxtDZQDAyc9NRTRon7CPQ7NvGaREyn5Kr7/+0pnYv
8Gu/k6YvRb4RstFixudvSZoNVViBxRi+YfzsTJ3sKzFEWApdZODUlXv9Q0912D9n2aLESmsHIgUJ
YUSk2T1O+Z0Bmyt9+iTHA+BGwcl5bw/sN9h3spBEHSOyMlLWfkkm2RbeK45dgPU4E8Klwf1n5pIS
HX+kHzuhG9VHdR8xKFkac6bqYY2BjyLU8+PamB+Sa0QLflSYGRFnP+D5kgUOquXfAf1jSnZI4vTG
ep69NrcpZ3tyx6pG92IwtyYJPhxGUdbiNBAqWyHY75JgGs3bejPeKdNM9G6T352T50gDlEUfP8n6
0jxwNquGLPFPP5cfFMEGwZcESUgBWiQZIGlFqfBEn9enDUSc0R3KG8SZutO0jrnX9nGY9lcZeJC0
qAIUzGEjnejH0jC3n4j3lvsBdkGjCrPg3RXCaPuNkEt0JBJ+tkoCt9QFn0xH6mP+KzOnRJfuv4Nw
Dp8mX+IF+z33+sMlSY8X9Idj6CSfD/+uzt9ze4wDN6G9KLmQpn6/Hx4DeIJE2BiNddJukfiAR3bx
241ItoYHQm1OTD1t1hAJpKDLyEWTliD42jQIqQMj0djsFhreZRtXXbjs7elYVoadJlGESjLqx2sX
kc7IfKE66urdIgZZRzBNiQmwmFet/ruOd+mxQ8mN+zjOBRVEIELXtxEbL7HZueJioSYR2tH3cMve
Mytf/GzRNQYOsDVbHx20zxiNL9ImAVl96mTCDWghMbzcHSVizkcAqpHy4AvkXU64a8TOEBvnpn8B
3fWF/up2sX4CruRR0OJJ/nfjv6HnYGFwRgBtdJk0x7ZI8jU82dNBpoKQ9F0PVx7Og3OmtfTM1pfd
cWXMCElfGpLjUchBz/3rIJE37Chilz6Af3RaOgLKPUOuWlkEoXicNYRxV5Q5MzvlafvZexRuGGsz
qP8STyR5WJyR3wog0glT0J8ibGhazxeS4HXl57grutwk7r9+eR5nkPQLbnHCQlKcq9vmJEYDYpw7
3pYKRAsRWhPJw1fT4EgNWmfRZNSmYv65ynO/Vwy5OcC0cAgnilN47wNhJdbOGZgL+I04tT5l0BVS
NYQ3qNiIE8UQPy/cWuF/XbuG21AccrS4ztpvLj+2d2ayzSRoNS7tnaHyNRX41CYm8dDGvMpch5Kp
niLLGPuBiMySy4epkkdyuauEYkognNYcXnR7amdML9XEYf1rVeKkSZiBMpviytR81NCBZw1WD93x
8BZoAJw7Wq/x1HQgAEY0pTtDNvsNA58vF+u2QUcBOIP3ToOR6aALedaAhGrlAT2QZMTUPRuDBoVn
GQOPcCjnHpJxoeCDfzPA05WpFvOE2E/lirdOF78QdauvbVr+dAoXx9ag9IWbLsG0oUs73wgHTT0z
dQUUlVPyTNyTsot+KcI04BsVMlK2M+QWuJfYohYiX9MKYNhkGXcQUoKXX0WxN5xCZ91LRJdq8T6x
NFVWUAJAPL37bEpUh2J9TwQFD1QhBBwKtLz1qR721y0DD4AgmBvlWZoLv2k9biyYcXn0nvfg5uW+
gsKjCb2ooeSOqLxHQOH93dTTuBlirz32gQW/TcwMB9uvYJ11O9LvN6pNZXn9X2/TiCZ6TTvjGuiY
HySyciJDs/t+Ey9KsFN7uae8b4R7ySkPZaZk1SaZrUoL5p+UptL1kcBQNLPT7vGbhbTl+xCSqwT6
USHntK5N1MT5ROioochgx6gi4hBm5ngYeP+09FLGWeA0XRuY/ccsKA7y92cl5z9Tiyhn7zIo3/3h
JC+nyBjNLYIdFZm/Av7e5WcwCbFmBk3tq4UKtVjhRzcCufHcbvyUKsFIpqO7jgitkBGJ7r2qbtQD
ZyoepIxnjSY4DvB4YeUk2NHdMRmftSclQVDjnq+y/jr0DKkbm6tYkKTpmbYdUJoc7PwGcZVl/E+E
p8jfkWmB9RtjQeFDuRwFiY3xVAOHrpbcHF2XX3eJXsJivkSmpbctGLMzGLRe76m3yrNk/BpKjipa
4/LZ/VDIH0v5WP/fD2+NVP1eDGEvrjvHiV1daWQKzHykZtqN+BCQepOZi25sIRhZPci7RQF1zTJC
/XFIqXXBwxqRw9/DifUGajkbZVOO2LO5PseOxKFJZDrDn38jGsGnLLLqEk4/2DLT2qLpLc7dvv0Z
3y50LbSIGtl/UODgEU19fhL1s9n/rZjgmDA4H6gSKles2+NlT3LuSsITCcK+JPwUul4uz9sfvSt9
94Vqh+4IYsSynOjZoRLIlAf/8dBelvItEZmNEEzg4yJvg/7Ww5bImQG9gPMvmOnPfssOtdBCuR6v
ItwYAe5sU1zNFzc543p7R66X8ag+T1yi8cDQo22sA+RzNY78way+X1R7gyo5fHaRhW6u9UAujJoD
lYeFy2vgQhf80M7E2e205S/EdurA2+oCyhCSyy3TtTPICHZwNB34eB3yIlJg5gNzXzbY3eR7Nu9A
ZJZkuRhZ5iyxyNeCwXTvvJEhMRnJ/5vaKu1HUdsn5L6DSVhOX7paXjvUx0oK2+a45PIVVcziyidG
1rfs5E0kGhtNgBOwZWndZgk8my0LQxaLl+j3LgiLpRavxCcN5nb4h+LwoByOcj8PW+1G4Q9qbsvc
/iOC2yXp1EPtSexyFPDO79m+5IrxW5ZfiZFaO6sao3XlFkCj/aciMURnG+4+W+f21uqMwbyIaEQj
mZuU+xj+fSLjGebdBFlwnZOzvFA9OPmZkL3Jd6r9CJdx4H0dqSfIcwR1We/ekRjMfh6gnKwSAm42
K6rlbO2XqNsvfd/mX+qQ2xZMwEQL7+i+lXRtKMnLTdTjCErE9mPhBIAXsyxL4+1UDaqlLYvgqcmm
IcPr1q4vxW40zDuWDhvy0O00Xui1VMz2z0wv3WLQ/SFyP3cW8UBImG38n4BCDfgTR/ztlGdLRTE8
gTibL0TXh2owLEg0fBC0RV+vIK19+YFHfi5GMKcGBheEJuRJY++/rnY/K2VS5zyT3DWesC87B0Ix
oEkS+LvUL96pFNEIUD55FxixgWXbTu/6WFV9OHnZqJapnRwaGH6Te+6NCEVPwdslLUwM0lsyI8Bu
pt+waGl1ilKheiF6ZaPi2r7kVT0iASmY5MDhscxrqDP2QrIOWpesYWIEVkJlcQlvbw4goj0YezPV
H2xd9yzoP0sMZZlrWTT2mJvZ6+IECvPaHASJ309Se5V49YFtA+icsbYhovd6Emq91hP2T9RhXG0o
deATkgQ0QL2DxaxaSvkdMN6dHKoCKTDFN4eKe8SvJ6+91xBaA4rz1A0F98zMncWnySZcRQIMAVd+
h66Ny6Du9UwR1AgBhxWNWIMjE4qoiNM2ZZDiUUHH8SomMDEzgAxVKUYMT5kKfMubFZpgbP5sqLiC
ZlUrxhjWPD3tyI2Qz8NTzGCV31qdwvW0LAWDVHa+ng9/3tFzcg7Axvy/O+AqdsXjkgm/g7JabDZs
VHMxG8KyjxkmPmWy1r3KLXlrlo162oAMtoCVQ67v2vsWQnKCJtzroz5dpLUH6jpMHyMowYttKX3X
JrPfSuU9RpP9LQfqIwITgVJpuYPuWTgDiFfm5DANjTrIF7maGIWqTzBAPPkxaRfvaQUfngw5GlR4
NTSPWa67lbzyPIU8DE2FtyV3pj7Z4cYY0qWReQgNNkvJ5CaYnXJ02nlBP/FTS9PFkRmiqooGtUM1
mnJRqwmqooczxNNVHuwDvsr/ViH4zEkyj98AGhb865ypeBLap1LNjDzY7ZvS+lEUjN0FQIZFtmCY
59EgybN3WXYKawCNVkT+x5mvGhNXHlgDG9fWk4lJ/SXozfulu9/3Xt0iheulPlaPYxIA79vjN42K
nUigvCvVvyW+cUfyHF07IVtX1nHz9Yvz4Jh30oi2OPOsDQFQLbLT3q+gzAW4ncXvQUw8YikmhEq6
2maC8iDtBMwJkd3dAj4JluHMYzUml8BEAjg7YILJEte9qSfMXAbzpdJPLh6EEw3BJ/u22vKYeb20
zlxPmrs7qV9pILqvSOn/JvQNU7yxufx0M0FR2mJw56kSfpKt5Ig2ThcIaUuclSY1PbmulW/g4H7q
BuviH4nFw5sanOdRE/eGxp8w6S6bo+7TKIXk1EHxFp2nQkBGotgzRdvSl3Nr/QQDaT4+3dSgb0UH
CHuFojYaSfivOju/MZePWwZOFa7PP4/XPQO7BTORSr4N2ru08FCV/qZ6lKEY9wbW5u+XzJVa/Pra
7iKUYq2n2ViECv2YH3gMbfizCOsj6z5Ko8DK8K1vkpp4cMeHQ1zU084ZkgV70mCG0yGldTH4Ive3
9CWF7i3gGx0ntoTVVqxX3MQCqLcTMFWnSWeZ+yz21FYDZY1TS+zjeZJF/Yd7emTmbEHXICpNgwtF
BzPvWa+VrzKJtFhAkc50w9c1hw3QEi0gxnvPm8A1lvZWZHDiZuB2zhUaIfg4l8wl5ZtRiGCHn8Xk
GEDHcYSiLpX1b5uXo+u+H9xAcEzbE3FwVDVTmKD/M440sLTaobeGMkImkmz+XBKhNSv90n1eA9zA
lbR6i9DsCOx+2k+OOfmcSe8+anqG3YWkZtQDwM2Z5wIfAI07nizTlLluIJfLHmO193e25uPeXmw/
GD7LqPLuq97RNycLnOh8ZkNbfDzO5cq+PsTkY6toyEwj0ml/Ja/6wccR8oF/vUwldvi083u7tETz
5MP65byO4Sd2Mw3e0swmJJhsmQjMkMLWLpIME8/mwcXxwqI1UTj7I6UGgcZYQD+JaI5msew+WcFi
eqhM4Bi8AEbiRhPhWDJc85aKC73su4cr4DwZoToBuKrzKIIKuGrMvJZt316mOaBBMzP+DKqkOGvf
9MtjIpIG6MDuduxAyfUEDXLFwQIqfnf7e+SPKKFahCWsZWMHIHdZR5xK45M5i6h4sxex3UMLQHgB
wT/NUysY3PxXFBGqt56C0+z16TT2eR4T+C5ZPecyQnQ208jwWZ6Vy1I4xg5LlZ103N8j28X/32QW
06N+riP/azd9tyJqWRmUcG3sOdAtdu1bC4lbz3y/RXOXCx5YOga1EjfmUYKBOs1n17CvhPQTMfRe
5lxjErw8MQQvClRAtgEIft0nQOqikVFgdaefzv8jHN+hcX7/53COr4zS46yEDU2JV9LVXR54rrjl
oLOifqB9pNOfEOXhFeC/+jEUv98+4dUTRpiCAxvZniuoGav38IofVNYvmw402bhvzxG+lQeD3CkE
hQxX2kpMgUFeO3CZpFjiNnQKM8F095bUPEDYInXxnDs1kZkfb0ZxtD/ZT9yln52//UtZmdr+l9jU
yJHiQjTRpG3W4QvfJeNfkeC1XqBOLqGqeg2HCqpBkKHn17ocmoIPu010CRfZJQGbNNfgSG4gjtiQ
MNNLjgutQvtpn7kts0iCcY+O/vnpMNDkX0axW31eRQzjwTKFtSKlYkU8HGdv1XW+yAaRg1kp7xsj
YqnJsl6hEJFey5Fu6t7KArOwuVqY/T7lYvImTzLHZ2R+S/bFnmdtfmyjA9JDsfkkipOHSZlJVvN6
dKEjQItH1NiY8t52yoN/jgv1sx+dntZZ3lK5a/noBIHtwuZgA7Gsj6Bj1dV4QXtbotd7/1xnwYji
mlC37VmvVBiX//jF1U/9Eld9wAkBPRsamLUhhDviDahdtU2J5CjBaOyBQDO8bnuhqImJatBoqqCD
d6ZyN6S6srqbL1pRitub5Z+DEDE0Kg01SnDhXchtikVBWiK2QmFCPvN+sSlWTxIxR5HWjFrdcwXv
Lhm0jWUykBKEZAGMvjtlTyAvyx3CeyWjw3TKStjuJjOWigf+atCXEL2lblbcvPNstXYJJeXALCp2
KSQm45TxZSN71dQ5RnpHjVfmusIGZw4uvLX7FvqSJYi1Y8a44NGbns8YU5XytY1sdVCBPGogYFBO
ksI30xkmP6KtY4JGoA5jZElSkjAl8IXSB3juIoF4UQkuLsQwgmxcTVaPwzEqLouyT7x/0tPhBHSG
eFgcOGuQ2L8+FmdwUJEVlgtuJnt75totnXcQqa8n0fb92XsT07B/4j/zEbOCZPsFsYxlZ5pzSmdw
6ICwo2z48SuBNKWVgo/MFIHaOu4m8wvRA/10LCz7IKaaoQaBe7oj9zArJMwguA4JDm9WCgh85ION
N0Bybfl+cR1yjCngZ4ITeUbuJhh5cxrf6g6d3G9c+IvDmy/sEfmR0lnyGXokUvM5PJvM/NJGmluD
6WJqiXCjXvNUqYF7g/WIL0Ck8ydxyOLUVAdSoRks7KwVUel1nH6lyH6yi1MyByziPLrVGV9EqZYV
sKbgvm3vS1bwFjVD1YQZzpVe7bnmjarfPF4KpGo8vpEbvRkQVlnSyToKdGKCcRHnu4xtlUcCOZRt
Hoo+t0PgC23OVcTGDXo/+i6yYXQAfg19CZm1GWbSdhS96LMACOA2b4LQCpcjOAMpAGcWYdulrgmb
8RUagweJsZp3Ieo4167rUW1FRpZGIwCHvUpYDqnk5KS/7JCT4/N5A2Xj8zzjYkAJXXGlzsXhiLoK
KXt5YRnfgyzslhQHDAD8KJ3MK+MMmKk/puJPzxJ7/opXY62kmTuLtfALInP9sKRIaNK9iP5+Kg8g
4xlEA4Db1hJMa7/GjYx6oCmvYesNEvmcU6SbkLSruVgoIaAFlESD4Xds/ODabtTlW8r48qJCoBdz
oVIXqoqAz3XXrGQU8iy01nRuNb085XjpOBU7taf2KxxygD89MBAXh9a+eWx17AZ2CPSP1sfQf9AE
yL+1MINE8yGVdUQLoY65sgthggaG477UdL1H7kVUF6VJhcRQx6mj5LVfkynxvSuUTmrCfY2EaCbh
yUID/Ev/0pzIFGoaTmw5RGGQoStwkP8QMESmaj86VHmK1hu3pvHVGp+f5/+oHW/MceLOMM3mSSgI
U/f8laO92HtInT73PyD1tycE6NQYo9Bq+wEeigzbaM6AfFA0d46OX3Il3JICtokoqYZ135jaIRB2
kC35vr3pMrRbFRVjc+fcHgM3EdEf3XOH9HScQ5naHHFT2x9gdh0XgUlWd40563SIFf/hvQMjXYsx
9INZv937gzoUUe6yhEKp2iM37ywdga3bV2uzPxHQ2AdHa4xAEmJU1zQ3f4JObQ35VUoK5ekSwVd2
eEEpUjywTwIrP5iQO2kDKKQHX8Cngy+ImyhM0LjHJZJIaZBnf/Fi7aBl0MVjzAIMGrH+/MREQBvW
wAPDGAibo/S5fFsOFHP2mL6sbsLzb4rIjSmNOsVAJbiiV3Wv9vwC6cfdvieamYUDBdsQyxZK1AB8
N9M031S76gTuFZTiPelsG7wLZlCmTE5vDCEBz2nLTyPbv8qEx+tiUzmTbHz/fL5ReSTJXWaxYk9m
DJqJy+OOYmuCyz1rwkRlYBaliA68eJMKBun6feydrIcG3yVKkBO+/hxK0Dd4gTuFLhTr4Znvjp+d
s3yfpZ9K5+Ttwc72gAkPrPybJkdYHDm+4xCXCpjW6t+NJ8BTqh8zcpdzvkjc7lXks2mJRAshTC0N
tkX4uywTapKIz08piTQIw+lYLLxztsPAeFLMJ14U0INdQQ8ONhIISxXCzxDOlKqO2HAy6K6VhlWn
yZfQ+I8qgiUEC8zXlCevs+4phy+AHLWZEiF0hpKdMAIkTPbHPK3mUGlnZdMbep4vyTTVEZK6Uhcx
OJsiPEk3w6HVINLDG8vnsmvtN9GlHIK4RTjDJ4MHy1sOnXbboiCS3uZNfeFpfKZuGHVfkQ14kDYX
aQLWOo+dSUOFCAqI8QzkzoY/qeUWDEBoBOGFeXASQA0lpKy/gwY9so70+rN0cUwjw/GTXH2I8rsL
IZFp7TkTZJUrJ5JoM2S4muCPqqVVI/VYJ9nnjHqev+q0aTNb2UUbQc1ECkowAqSF7LpHogdb5TJi
PMaBJIxJD2qmwBldQgknSjuxlXch/nu/ogP2+mr0Yd0Nukoq0ubdqNL4qWEgdChcTUbXTt0CNaop
W1FB/bpmEqvLWOUr5oNZ257DZtEsQ4PoD+ddId2PnI3hAmx0x9xXvLNVMX2VVnTX1cgWfJNEvkeo
4J6U9lcqNGVApXve1Zytga/kPLwdNyIgrwv9jBG4eAHXvOk8jWrLGVmBmgXROenota/FX3yZT3Cp
/gt0UoWhdw22gY/3EnSvo1NKHqo/Zj2QQLse03GTBQk8UAp9jAvv9hCUC6P9/5YIbvTMiLz3sqSM
n6Pu+ofI0W+uw00r5CwG/eN48qeNgOZl22jDOPV8wcBbD5ewRZkO74XgeZ7LtALh7fRqF0kouUwr
APtrFQbr2rhuBg2zfd5OaFjMASvt7zKVpbbznb8q0FY3MAINW+7dfAF1L1wWdu41QOgfBxB153Mz
s9pJSbBPX/rxpwFuMv+RAZPZ7WI2pOmawEctlqoCEDEZth0wy9Ya/MKcjfjykkLIzWdo4UBVfCRC
gBtlsxTGqDC0z4gZPPeWj26UPb1vk47k4dOt61pO5DtD+qI9vPZbGzlwiaYMrw8cPO+8yvR8WhB8
IA+fsLNHg5Ha2xP6ujJjTK32uY3pFpyUoazZAqnv5B/CfN3joB9Pcp3XWmsIG+oICmd17xBfBDg/
MCZd30hj94GAOceq1z61xSD54XsMRZAxYwAaxs7S8e8EysfOoUFBxR5GFw/es9Jx5nDO9xVq50IN
f0Naw6L0cPRkhhWFIrwTfqQn9Tzlm1KwPr/wjPaozLDlpzj6GbtaS48Wx3p0b2jXQsYxZyN3crfB
Oa2d0fx+wlu+WmgviIkKIhe6T0WQL1vjt1eoN9J1/EvIu0VKqFY7r3u1qB9/RgSLIIvTXDw8SVx7
ZCIRyJhnpYht4jllaxFIXvdsI3YoxcTJ6Id5Atl41lOidtMjDAg2qDI5uIDZQsOx4BK8iBQxG6m9
DAbjEuRdvpumYYRs1k48jIRNewWHxwAx/A0+3BKIkTqNWx7XyRf7hOfen367cBlzlTBRGrXcRe7G
7sO4Z/bpX9uruuTrZVkZkHiJGEWPMGig5lQzvtxNeKeFjcIyS7Y41yOf7vY55u+Y7pHGiqh4HMLl
InNU6MsBWJDU9/cZCUoBn6n4tO6q1mCKMu8pySThwSDu+DFwSdF4vXTVCVSwrXkXN2M620tTvTCF
uOU/AFZhzfjS4k/MRrTfNjS44YzNJYDchfwfOPh3VVtU3hq4ClHFikTx9ry6jfCuhs6w4zimIrnO
3BwbFW9QW1oGQ4UW5Yw29MsYGhdOqKc7uvlpN2VW8vD7npct0Qmk/bIFOazjvh/4XFx/23a7eheW
Fw6Gw7falQndpA8KIWkWRD3jRfabYgiUmsjHY5LF1xyq1VlyIfOrYNF4aeSgQFzYvM+ITGr7ZJ+T
S92swGTqodR5Rf7UU3POXQoswqRtTGgL7tOFrgFUnRIWQtqHRG/iXB2KlNeIqkB1a3di5iz2rJL7
KdZhTqEZOYPsQ3hrKfzDfLY9/oloSYxn/8rJlu6fbMuQXhU2hR6AdyPJoPb7HpPvx5uDVJf/kYEe
2uvRwiqOEbfCkTCBH3Uz9sAoDdSgYdXhxYF4qTnqHNH7TTvJwXDZGiuu5mPXpLZBw6/zW2jXz0ee
gFYtuEM51qsCxNQm6k1OIa4DRgJpvyHDUjxVtcIr3AoWjVWtc8Lin5buzJrtae8UR74sk8UNCoV0
dhMn6+pZB79w0nkmkZmFMRgQcVJZ8ndWMozxcSFXCuTaVy5f7dyxwPYibBYNb8aqLdVAG66f1WzT
0hSFW0up3NnJRtAb6Mr4sdvylxMuZ24HWBp2zRULLWgwRQropwFwC0bTChKsVkcltsqUZ3rkaS+C
K19mtw/JevB9vdNo7oGvNERm+QSNXCOnEe07dUd3GADjvCCTnvna3nWN/CtG5ecz8IclaD5+KJjl
fSJ5BbCZx87EOLdOFxUSAsbnOQnM5LhGT+kqiOP9HJAeic4do/+EKa5f6xpq1eJ41vFbXpsjqOuo
r2xLJ45fYD6ljPtmVGG5G+de6FO0QGDkILbcvNmjsvpGUU4Xtm9QPcQcfkXhvX4k/j+Xe7+ivJZ6
wZpnMHJ41GBmdNQDCkDWDNMQrzVWgh5+DngQvXaMOfjtFKMFNPulZOzgI9ClSmYlET4UjkT7BPwL
wGSaF+WoE/GlksYosBC/cwgOivMKgKytxKg0sThpMbSpVb+l0n3B8sCWOh3Z2q8Mqg81T7auULGV
Ntt7HL1tkNAJAOT5Uyn8CnaP1v4eDLy8J1bARmx/ZNLOslLu6PZ5B2M6ArgBeckesHSeCwJvvuOu
0L5mii3JhF3e5TMFQmRkT3+YIJCjPZTfYSBKzlQXMqF38V55BMWDlembxiMjquL8pnhRXXjY/Fd2
E3sPzpbDDSLAqMZgmJN2EHJM9BGR1XdsG2riQd9SDf2jWg0GpguAi6U0cQflBd/lc7naD3yyDC5A
FxIZMmiDxLqz2jee2R1B9+Zn0S1Bc3+QeRMCJVoUximTjhk53cpsJSQP7wFzsCTOyquJr0179Iu9
knYDiE7mkdJx4THSaN5kCDtuNMvX33Sd+Gj5KRo95n4DENbghKOjyi/N9aRov+YY3fGKPdGxVWgo
PxSZsfumj047AewYG5GLYEpLcNn3BwCxTbqs/neGvD9VjkO0s7ToQqEIk75dyXKepMsB7F0XL0+d
4zCeopv9CfDL9DS43o8jsHKx5fy+nZ8D3MoP0dfRgda4NOqTh4O2L6ZzqCeURwPBnw0KcrIHWo+i
m58mUeUoQoCcyj9tdbASWThaRlUryOJOyE7QsnF5YQGtsNIIjjWWVKJfO5aWd9fk+uyczbcI3oq4
6sIeJZU8t/Il64ECVL5Jt46ftHDsESYxxUS+tOFKd1iWtsMR3WBzLGkSinjrd0KyKm8ex5KDXiUL
IrRwBVw8EaylUuL3YE/jvyA3KpC3SSo/kt481L6eL7JNRuZc9bP8wjfjGL9I1i8G0rTy93B3W0H4
qWlyPcE+07Lr7slZ+vtZ50zai0/7C7DOliwD8/FSX9KRcfK9MuQT15OfsVWdo5MROl2bNPYSQcNY
9Xpr6SkYTRWAGEnQit8FKr+2hIHR4IwKHkYPd+v8lq8gFBKphnWDiY8Ps3mIWrRGpupQkpiV+EbK
8+riIkSgqVnnKlUBzAc4BWfUIOv3mRgKLYkFPCJX38r9oFL5HAs9oidRJMtOSZ4Zt6xg825+dEsc
5+0ZHw+GQDihU+5elN0e6yS2sYx5pusuILr/32QNQAni84Zhm5mF0BKkxwWljDex1pQ0I5cHzoxY
nu2Kpf9JC4P0oYK8f+Z+suqRbVA/XsPgErwpblUL/VIQqdJqiQF2tL4N64bLBFh31FGnH+2hwOnI
v+NdbtGzBJQdKEyDrXQ/FqNA2pCm6uYB52RdYWjDa907rzMa0bnHFkOft3RjasjvVNbBCumbH7FP
xn7f/8zjSmlhY6EW6xZhROAYXoatxVAdAwK9GNWRq1XFxzlgkKUzn8AHc3LLyDUnH98ePsxOZ0Ry
fZ60ni1ez8DtbJowu2VHyHzushegvvXnFp5IUHSz/PxMY2tysMNKnQ3GTFm96LSi/q0rVf0gJPlT
98axIUypZZGEc8+xpT3fdVk3DQhW8Bp1FGM19awsVEBLf149UAum7Vtwq3epiCxncNPSZ2ymWUFD
hnxqCaK8pmuulxv9UWB+BTmj7alerD4ZIzotJNGDUo1Cr92hYGx9hAyUv+FT1EQW61Bmh6OrHX3E
DWtxy7Z1J0kbAACvUqVlyhovBBEWPz9RUPfc+XLE61LI8oceyY7jVG/Y20Arj7sJy5iePKymjf+B
j8IUemnwN8ffxNeZOJv3K5cbG26SL+N/oz9PbEm/Loo1AtSHEPs95HH9WJAxMRIZkLEfxbqNCuDo
ANz11bvSSjzoed/YlEejx4HWMrXItpFdTzBTPFY2fltT9hZLrFEDgFaBf8XcQzNq9rPWJLKQUYTE
iw4kIFpeB7LR6bOUqvelOpuBy2Z1Av0n92rsyBNN0QUgsioQ+VNnlaXRHZ0GFO3DvcXb1Kb3Mon7
B1O9G2WzSOgHON1KzBknXDf+PWYeNG6KqfUbO8au9bZiYwZUF4TOdrr26ng2/kh5uqYiM2DTOLNu
3YdPq59WHWA7A3GybN8QdwWOzfZE3rZtCnEaRn6wETMTv6YT5ZkuTjv+4iq06AH/HuL7oagONN6i
uxPwd3p1l1Ad3hvUNTef5xiwIKg2OZfz2Jcp0bp52lUjtAt1HQg5MPmVn/ye+zwdo7cgy4amgWBK
+Lahut9EksZTm843m+st0StfoQ77dfBQau8ZeaCZ27khcUyCEtmp4YR4V9PabyvnlVUEGFZQ5FAb
D2h/NbTPeHmMfnlDH3FDuoqj97LogGox2TGdDBFn1sqLl1j1vOGo5MnpcSA05q4ecqxp6hGPxABl
Gj9eung1dW6HM8fwuNMOSPk+JA+G37q5R40GIhsT1/9McHd9hXfPEzf4uYwB+HDSPHQGCd1OkYjX
dyIzw4g9iP9/hdjL1l7Akn0ZKJpmaEDyAmBWrdXQBz9ikRhZ7ddqpZCF35vePZ2pgSphTCEeK39y
3wN0dbz4oJgDn+UT8cUupo5AbdAoWtqXnzVHfAuUy2F5eyfiGhmUoM+zxVOu8Se05FeSdrAFNslu
iFBnxn6fzbjGc+ttd3O5l4q4S6fXlTAMnzfqQ96sgP+HWnMGUYwRMVOfen5AXirOw9CRWsGlM3Oy
GCRNZncFTC893WgXerFCtQepA+1mUeDYg4U7v/a1goCDWPH70PhWfK95iO8DK7su0JOVuRZND0cZ
neRJUFXV+UWHPnEsRJ0zhFtPIgAx9gWHqZKGpYTZCSW2epomF0LT3OWZTQL3NzndkDHF44lNbcCg
zePDoHCiROTsHME98mrJ3HKqCSMvcxgUmqPXRQRaOPC8bnm2bjdO6+/gx3unpuLhj+mQA4j6Hq4G
Mp9rEsyFA+6M63xOLfFwXajUM1uktKhjzQ6XWh7G1P7yvc7rWSQAs+c8g1tPtoA3c3URmgIZaHZP
+K4Wuozh15BlNnjYBqk3ZdN4HHVWRrH+ku/suz0VbojD7oZNjfeK11XW5Z/4O9GhEtWr+9WcyqI/
OfrsgDzyBHPnkXfsfxnPfj2FO8K4aBUwpLkKqLW05AFwERB4+Z5xobZsWSsCuMGIv+cWufdzb/5i
12Z7Q5F6TVWcB3Ue+21mXVg6L3Zo+fSI7OIS6K66tXEaIr+8jnIrz15iEbqaBapivh6NIrOleCA6
LCNf8KsMhKf9ldExTbqXnCmMBqsWb+RjVhyWnYpXCfwUEifIG1YPe4l3X3FYaZdNba1UaGkB1s8M
hn1hSBhQElWuRnMgkFSMuFqjLojyik1rE8B8UyT7GhHrOzKLGeufmsaCHGyurbO3JFH2Sie1gnbB
ghBrEBmoLC+BemvNx3F1pQk9NUJIgZZZ8mRlLpui6Xhg++v0t6CvQajG5s68Oz/mTQuufOXhZn+6
XrpVlMdh3CZIZjB2NVITvXwR9SwG33cNfmOTVBLOKHMYgmCYgRCddgR72dPqLMKElsYZgmBVtg8I
X1nw0xvioUso2vBZyoEL6OEl+0NGiBnaYKV/xYYZYMHyY337bh15V3OpzcJUgt2t43FOmsVRUCJb
3Cwkpq3p5pSEFS5kXudjGZZUhr2WLd48YY2U9O4uCggxX8IWEwgbOq3MeyMebf4tptn0rqqh4P//
AKylr0vXm6vOJu8zr0ezYzMoBS2cjdy9X2+VQrkOBCd9H5wQZ+zr6Mz65j57B81YaMPjpGP3zTJw
Dh5ijfqpyHVSbNFjoWm3j7S/pKLHBaR6m85nZbLlSNU4u9o9S6JFldY1sKgdTZAn/hj3az0Hq2kV
7vQ9/BRp421XT0YovB8Uf17KiPTxkKm6yakrmDgHxHz7+lccLThZlrhiQAEcipwL7cq50p4awpdV
iU09is4frAc153lOmrcuo4DEU72Z8q76j7AnpYLryhSK6zHyu6FapCzVFM0d1pydI5RiCUYQhaBK
apUDnBG7VF6pVYnyXRN5J3ISbPyPTYtKCVIMWtrx2F0UM4jp09mnIR6oE7nd88J8psRd7HWfDaM6
kTChrxQ6PiBTqO3SpKaOvI0NzFg6YgjQsXTSFZsWzlLFnBauMezhN+56xCr9yyAW9puXxOfK77hb
54DkMx75q/W7Chfzu4fkJyf5HMNr93MJZMng+AJopr67Rl9gPwORA8ZBu6Ph4aAymrL0l8tMNl/q
fUqgfKWV3GNh8cVuUztU1+I8iykmW/jIuB6CIeZXkE8kKma3dcuIBs9rxRD7Pgp1evN7QA094EmS
Pw+RBEuHwcH/KwveVCFDkusp187pkjVDwhB4bCyFphdI+uNAYm7wpmKWvojt4adlKVd+T2c7T4Zj
kbFaGXvD3mHyBRnDEz0azT4/Y/UAhXTatkosMS4LHDbG7aF/y4cxPte0RtcH79kbJCbLlDDjSbZ6
CjOg661abFthLxFXchyJea+EYXKLAZrbDTjz9y9AID27pVz7vk9AxrOd2/fKV2Tbp1jN6b/uP2Ad
gBFShJSTKXME70Z+vcRoXHceS/4q1pWJOD0aIhELF2QYsRckOxnOXmii6TrVfFAAghL/EnwjbmIz
yWwCqBQRVBVfj/1Kyj501XKyJmTZb/DKSMMQnQ8XKJAVr3RXHF9m1G1fcdWIeAex/VT7g7ctcvE8
7lO6lhRAuOJJWsimRRfLkQ1hARL3dbZPnNK0Ng5uoj5P2HeiuXKIFx6OemK7j/7KpEdkuwXSpdGf
u2EyVZxeSqZ8tm+3xbZMUd5fYVdOfg6RkbmRMPd0TbthI8zLDloFWqtw2gJgq3ONFg7dxP3/W1GY
zuTw6RfnE4O9iYeDauK3JI3/Ymmnr320mONKdl3Vd5k/6jvs+hGhpzuYZx/JnaNI8I9hdPeqafLS
YP0qOabHt8j5bAVTXNDYtluinWxMHg7+jdMhjxtFqoqIc1Wrt6JYOI+hWN2L2De7/6eEekZ9j46C
brw5j9yIcJ4VCUFD9AUOXoSDSk2ZzYiS4xLXswm7JcM/cpuKGM2ErUclsRxvfb6zFN3/ttBIiaZV
43hAV48+VJnmF7OwZMwbnNRePwkAXdC8TLE4eXN63K9waqTs6obkjqpaVIaPfd9cjHuxXRSFn7Kh
3lSvJigiap3SPk4aXeOZ1Y3eNIe91Agm1ulykq3yD4+KRHPcSidw4mtHsS2Rt58IIHwdVCYBv6BF
nuabUQY5Kc+wX0y2100U77iR1F6EUqXSnTWZVV8X9e8bc4cU1yydBFTra97gUoZsvd+bB9EX8OPA
pUFWDbXIwMmmeaWoGzjQEEyBF6UUrQdn6F6hogVevQh+lSamr/8gH4+XyAOsy0nwice0IhQ5EX9j
d8kwDp8vmNQHTPEFrRZVS/AW/u/mEA8Xh1vJHRnhyXosKAEtdxSdT6OPOAwIfyQ+f1mFyIVCx5y5
/H36lJJtPcMwcmiknwk0WXd3BSLg0U3C8/7P3Ke0WheTj7PZRQXbCTmU1qfuqtnG42V56WI5pljM
aOrPZBiVfpn9yop6mng+mbGKbIpbDWDF/x24jy1mS2qV8Kjug4j14cV7hxlWDLaGgWl1xWl8RjJd
EHRbuedjr4OuV4KiRrRQ3ELSrBQs1tpdBoXrcyzr7brehygHMmlAN4gcUPIERD/fYaqekDYAXgpP
fLgCCO/0awSDlFNDoQdWVy3ybIyq4c1Z/Ryx30ioRNyKrcv5LL/qABFoIWyhEa6I2EbhlqtBMein
f3X3jhrBwDLYN8rJyXOg1IZjV43r1NY6GAwu7Rqyjv2RiNlsBWzuiFoyCd4q+h8eTLd+rCrdq3eT
DWep5ccIeSVl+mZVl9A02I5X0Uv8E7APVKwjlTL4YquZypkrf30fRZza/8LPvINTNOmgHnExNz0V
JHVoGouk4czFRh8YZPAISD5jWds5LVXBWoRAP2XMuK5qTxfiji/Xgb03tXGvrWqN/e7izd852Mgp
8pn5wHFk475+qfQ2yjcWn9+NWLRtIXnCfrvWDdTpqVUBbMBQyKDXdq8xNdoEyo7UF5M4gebHojfE
zSNMA5veAbtddU/+F8h9S9tOZiNAMnr5T9M8of4JYOwKIBilEeWNxiLqPM7Mk/2bMcKEiOIgXPx3
4S5OqrFPG7GKROOqjAydYDXin10B6xXoarJ8dZNK0U7QaVVsPFkr2j+7gq6hLqJVgsVDPxCpV6bn
Ij2QUKEhJufa8jOdNyQhTG7lJRX2uh6uHuBpifl/LFdeYR5TZbHsB5lDizMBiAxCfvdSLtgSCd6S
nnvqL70ALh3bROtkJGpCxYe917te5xFkbFlzNdxytK4vKbF4yN0QhqQAmasPMoHFCxKmTMuaeKRC
mgQc1/iMoxu8C50w6lCmEh6iA+GhV4PX1xgdeg+GsXoWY/U7Bdd6KVoZC65ZyKSDLxQuWwGFyGpK
QdaQAZdgD1Zxti/sZifwZCHXVx2F0PUhkvQsECHzobF1543Aa8NLjYM1svGH1RTPlU7lsfQZ5DY+
rVR5iNXZsojdfPdys0l4osw2ZFJaJbEl30SDfFv5E1d/7/57VsMr6/+Qi3o5tE4EIoPa4z4uXINa
3hZuS0aI1kHHjn5jAdPLxaZFTfWxl3FIbXO6FauKYDqrwO3/wxQdM/f//cEzyVGodxaPnLt3GLFd
cH6wwGPV5hVbfIUhTCDuYNMYUv64NqRwhR0dNw25Pg4Ias/2G662YdkY1XXe6kL65sBJpDw4C/LH
N2pvTApypin5bZBHW8lbBERc2IKsxnf7fWl+flRd3778bgGwJ4NUoF3wUUpPS0kX9fsUeZGlC/CE
YAEyJOuU6BURT0k9Ut5GoVHlH8V41OUANti6sYHeueQxg6PWsQotwL2z4RIHr0sWD6FPxliLGWaA
vPcOqtITA79TE3oYuPqVtI+FK1/RFqajyuWxUXwe9sTmZr+dbfwshb3C8tm57YC2hwcmrUYr1aey
v9wK7HwKA0R+zT/US1EWFH5MfYZBf7PBKO0fvJDzj9O6QoEM7bc082WfbBkejHeF1H3lgVUAngAI
P/zp3lQQ4rZJe6NiPGEBi88rpJI1vOtfS9QUjyVmmkm5rxl6kpU7+7HMfG4kbQmOZZiuuevsYQ2v
6i/ZVeUwffVV0xtnepbUtg+LiKwHqE9R28G+D0gtzEihrXDMPq0sjjQMmXzdjXRtiUJg2FLCf2GM
8trN8Nyh+NBOj1Y76WbTsrESqWa7fBnKqfnRyUC47oPNAKBQhEgZi61bHV4u7EfaxGAHA9iLsaWn
wsPCn2+XL8TE3Nb+p6q/cHmH+/0zOmW8cIQ21jW+gjR8kftVy18oyBtFs5H/ScObJcYfPXJykvpE
bBbjA9Se8qU261XR/djFSjikpZ5nva0Bz5Z6T5xqx2kh67nZrylfUJojirvIScI4KL82OIw7yqus
hZKSGJzZopn2h8rWZOQPwTIcow/YMrp784iht8IBvi1jnus3uHPNRNqUsef6gKG7cUUt2VXLT4sF
1uPUsCTGNURQ/ovumD8kUvPCu7jS8sETqn4LKuYN1zrm9wpZx5bZ2wJVkyn9tnDwtpkLaPUAXSxr
nXo4sD/4Z4hUqvBn1v4X7RZgAFg1p8MjnU247AEl8H+ejthI+fSAqa+Lzm/g/es5k8e0agtXivmw
/3jEBui5UZkA3TeVUmlohUKt9fiW7vJsI0hJij5ovuEJYEOodiiI3FF8dZUiaujlybFmM4kdEy3z
BT52k/IdzKRyrI9r/k5dP+liTXyABb7bzLqJExAmfZ8BrSiti6XW2RaBhyfkDftqLApADBipCEA+
S4uSWgZ9LNc3+p8EDXDfQD9+Z4cxvE7qm5e7LtpEnMZ+smORa1/fpjCU249DotSLxM5tsnNWApGx
ugHTWUn3YmpFmIvpmIwqqA4xXvMMyZLGBYsXiXYta45jf9PGdT32Dh/ezdX9anKLsvjolInLbIWn
vPun3IyLhZRPgU+HTvFgpnj2J6s2FEZ4p2KXa2Gt9BPLvdH4R5y0ImFnOLxDngWZYk22myjtaqHC
XF9XN1KH9bGCX9C6PBotGwIMydMaongF3c8PPdSf5ySxhFQOKF90Q6/STuEEFRPOWkUeNyRY6zRW
pRGhh3esG88NvBk/o0EErl+OYyZ24m+V6wtCXmF1zjccuoEmZKoplytsMJz6LR1DC1ejgGm9DaMn
dL1tOYgAJS+CDkDsLdD/N7Mn9Q631tcCm58AS1TGITbBdU8p8klIDTQsJAw5VUx0JfOu6+rgkpTp
Q76U9eC6cXicEGINM46WhV9RnYXpeI9mkCoh39HadOQrpxZRBSAZyY1zOmv1zGZ9XCc9oPFD8Iuk
LQVuy8I6ktCFjxd9xyZHLx4NRk/FAMW82uZ3v3lISSKavvz7pTnvmYXXOm+6VQdzPKIS/B9A09RY
O3NNVW/H0R6iF0TrtoNXIRRotUiopkwm/d+wWbaJdP1jesfWQuJahN7+YOjVLcnP6Y2e+wGOX+aZ
dRGU14gr7OlzcOUccEf+lpBHUE9IuhRCXrjw1WS/ICL4rNOlloc44eb0hfwEy+9bdbNHsIHs3QN+
ZqaCB19hNNWHsYXWbBYjjAA0tyjYXt0xxyAXKrd44atydji7twkqFvnaOXg00s/91WIdddC13RA2
tmbBW305kWfseHOdt/AzIvxrpHtVnKap04dtGtij68IIZHhlkMn17LpuKNU46NHqMudIyPlVAQHj
c5+GVdqWzrk4eD0hcwnIwsi45wMzU/4ZuIO1UGHCIkAWHfwM3rR0Wub8mc4tSO+72/l1xHQ6SgAX
4jRiXJzNWaRk3CN6wjE6Q44ur8Gp0Uky5KrUwQ6ccTT7fAo8/DGui9a8r3MBi84ZshMC7lkaLwAu
yIuMmyYtrVIE4hVa0lg+xpi/8t90UxvaL+NQP5N0q6jMy/HDIn48mc9s4QRH1N6GZ11Hi9X11ETU
kBp4f2exnARQPeBhgVifskqR0HXrNMlyjTwVL+TDASbqqv4jIFypguOoK6P0JpNcingziIvQJsvK
sbNJZSYvjDi7gwWSptN6wfzNenNWqNN6TOx85Delrh4GC6VeVZ9vLgPr8a6Xn7lwziapTqjWqSHs
p2y8tKkc9p6ECZo5FZQFKY8lW4umw+j6gPRM2WcEERJorCFvfYmTIgxk7Yhjg9pyZBebgt4zGNiL
+7niAa6zjvPknNKsLJlG6GbTgNGfl9wf42j2G09vGLTQxwwQ10cdob7NcnaqQAtvRVCxwS9Y2ZxM
1/LZlwGpMQBj+gkpO9g6bRDsbmTRH44hiuL6drgAhLWRMeEr9LeHqj4bA9XboHifW/pIv9AUDg7i
W2h5hkkSXjOFu1JCMCGhZxEU8ZtFdXOjr3XeNi6jhi+B5GkhWUMg3gjvrGEYZqpzVqiqW46zeoRy
MOBu0XREtCmfCZQOmE7zlgZBodApheqLLMpnCeOCn0UxJ560VwczIwfrEVa9n8lvByu/1EzVegGI
S6YIAyu6AtdxdIzON8T4uFwJPSB7HRSji9PZKMWDJY9qHl8N0TgcRvE3XDQS4+altQvUdquLNak7
L6utPtvo/dMVSS8zMq1BbdjpQ2iCyCG0qlyKT4H5zDJ8k2sVOrIqLV0LLgv+cae9GONIdtvKjZwU
/Jbta0gvMbu/wB+aRYQQr8J6CjeKBW2sviCWXU0Vf664LLsZRDYaWA+kgkt3Fn9ED0CG9f00GLjE
vPvRxouDavHeDCKoL6Etr/KgVzq7YTHJ5tec3y0TAaAI2hk6Iq9k6y+iwnTKQ8nxh60NWT3cRYYM
8liynWQu1NggWp0DxsFDp9rsWFphIpi8n3Qb8niPMZ1NrptrWzH3O5NA7vkjnhAFO1jYk7nz1uKq
DoYaYxAO2RROUfbSmi7OlTeaCIdws1/tkewfmlnUes0ToiFiaIu7vqfT7p2nGXMHYs2IjXDy2vF/
s2new44uKPORcYwbb8YFHsDspwGuWKqOirzO+nhuzatgopF9RH+UHv9w0iMH3j5/vHPi7Fs3HT9a
9JLrmsz4FkzWVtlSs13XoosGtQYcWIFA/A3PwXp7VM1aKkmtOjvrHkpEA0dCkvR6Vv6sxbsid3Bn
fgzflGhCV+RUA4qkJ1NNoWRopB4hP2IzGoI87dVTo+JWApKoYmTUgEoiNAsARXvqZn/v47llpHIx
HNCMpCU2M2s/NpGKo5HPaohe5V6R1suc6bIHoULNHM+0UMtpplI8n9qUzfVU4ho5YrSFlb6zuS1W
Oz4yfCIO0D/Oe3Lzs5Lt9p/VTaRe58vbDCt1mZOaJRd3yLcN/8jQ5B3egJCk5aOsNKZurEn4RAVt
wrxDQwOthSA6IZlLby+qstuUoVqt7hBFeAO44K2ucOmm56TrIoxW4TXNMVgBZ8JD6FhO0gwnFulW
14UPrE8X6UGZ7OM1mCcKGHmcRfhO3+kKkqe4sEA1ct7DZSKnqBt2hLF0Ostxim5vQInc3BVN+q85
4ROGvoJmdo930SUqzItwmuGrpRIXVpWzZ3Z5goPM45tchiUlI3IQuxgxwdDakuqeFdm0zOhL3vO3
wLbo8b7lPqHsRPuEGueqRW0jyHR3GMZvTVDSUIkLrZ8POZOW+kyy8S5orAl8NjXS+AwAAFcq10x5
4uKnh7LaAGLA67FTsZ0vDUN2E1Sw0evHJsWnYVSaa0JaWIH05YxuY5Hx9TdbMh7JFlcMoNk70CqT
buWK3qmeuuHmw7tPufCZBSfO8knRBDl3KtXQF2BIDa3HTeVCi3pdjxF/NqEQw2Khu4L+8au0ch2t
eFQeZnsXtu+YF4PjSp4k548mWOwjXdQmFNzaUceFraMuwL9U+2CN6Y3WGyyE/XtLMsquzrrOsY1k
EOxZge/eOMVKtSUOS6rBmiA+T41LE3IOrXZH1QVnQtK0bPA3lWiA1176h11gaokUgi7vjjq+q599
WDCmWLbuP5qBLFC5bMCRzqhWdIlqpOYhYDTmOBPdJBX6yTv0Yprwp65y/iaKDiNlq2LvEJtGzkrW
xDlWEAMwRO5wSc9jmRYSrzt93xKgQwQgu87qzORaXVjFdk0jy7Y9t1oOmqXzIfuBUA+nS4hDkUe9
GSHhXArvy9b71jbBnmsxbtr7qnqWrp6GeomsjXnJJN+GrU7hmSUQMSil7ZXzO8YGdNzSwZsATwFL
Ck30T+ZUkrc7om2VwoBb1XF9eMhM0HzxOy+jP12msioNhc5p86cBJrePwTWnku1mfh0bAIq5a11m
Xm4CsmN+Pd8Kr8vdHZwaf7G0Xk4envYl22FYl8SioxZ/0WRJXM6a9h16ndna45zEcOrUESysuXa/
d7fVuHFpPXlw/VLLdOtEbD4FhaXoyfQS042K8P4VQVWVerfYF++0YZJbP9Di17rBifxPtgskHhz9
vWc4qro33XEv4p0VyIbibasiLvMgyRYQQwvjjUKMcLrS+uaXJORgEMn0uUnXLkbQfT7iCr67VjG9
txs29pZupNV/ikMdaP4YPh2zhkwN4rN/jgvUi29JC9x/tCnXxxNUgXuB2lJChC0EiyfvkqHKXico
yVvuYOU97phV3xKYkoNZKyFvZmY5PmbW+GUAv97ZceaOIaDpWWzlGO1ucmv2Z/Elz86kvqDWTvLn
kFxHnnEGEOOL7/C7VyuAz9Z0QDAVddac1RKYGccULuQKFymPj7iI4kgbVE9w2XPJLHsqvZgqS7YW
hQX1jUkl40CDdDw24mXmCn6igHMWmaSMv9Rcwz+OnOawvWCQpcK6rO2xi+JiTtcGZ2HlAO9ciW2c
anxJT1Zv/7RePUhGz+tgiBacIDBsjCf6V/BHbyG0K/9LWSqXbU7PecQbn9R719vRJmnTP57yXCUP
5MB4VAdCaHvxpsgtnfhq3trlRHpa8XneeWsPu2OzzQV7mdMszNPpXzw2smqvRD5OfVZubxOctnj4
OB2HNjK+FuZRLjBnJ4hfBhP7SjRkrf0nO1AVZUMiLdhFUci+znFZ/i2QoxWxX+kS6vb5tOjD4knI
yABgtp7Rw9Gyd4yjZkVnwPj2daQC872pEtF7Xx73Y8DKt+hShwHWcHAkwNysMMoCmGbYjnxKeZnl
J+moyylbLShw9yOQTerF75evc62HLLFyAa05/Hr4L19Gz/+iPHCZ5HahWvw9XS81JZuIS9NoM0Ep
71VBzax55od5MZ7oM81J5DTKDY3hpuNQIQuDY+Zqp12m5r6BJdnxOQpMm3Hl90TatPxcKluVA1dT
MX0Z2oxxCe9jyKcV+KX38wzJXz0EJGVb/9aJ/FplemDUNIBU+S72ZV6GEsghQ39nQZsZMpGPRSX2
K/zS8Z4yHHnWPpTO6Dj2ylL6/lFdfK1/io+sj3sR/S3Y+ivqwJAmK19qMdJWfTN21dVccgdSA1s7
EbW0KcbUGbIZd75L62MgkpjvteFYQ2be91SHXyqAlJ/sB66gOTr/4BZOL8OrqaLsEx8J8f78KNT/
GzSZ7E7y2VfCW9VXj8i3lkp7vF6Q4xfxJ+ptwr/ZY8ODOqiJVH2rOJckU+gONPsmbhZsubmGFlRj
jlHvoaz6dEBgWh2bN06gOZVHKE5EXs39Gt6o5+MURDXaYT18DPv+KGlxBu8J8XKZr27I8DfT6uGN
wxQZ71tUPhQZbhpKcO58uEVg4sCjg4vBcJ62wNul8vpiQeQXMZaEjuwN0W64n1S6xUNUFyXSV461
+80Tku1LX2QJsKLTYoWQewTX4UnOAAwsWK0GHB3ACGluy3875IL2bi52eV+ev27qtGxglHNyBGBe
+SgzzZ94Dk8Z+u7rTj8PZTFTVBRggFXLITuU63Qrm2ciRB1DZLx11r0AR1htRRoTPoXChk3NfrwA
rK/vS9NAL7lNh0X/jIib3iEJbJyU88Vym51s+qu9ej2GN/V8gv5a8KuS2mHSM8gdEqxapn7NRF+C
HqFG7fpYOJCVpLK9wzeUpnEglwxinh7cZgi2paWV6rvcoCIirc0uUyxMOItY5rvOOPIIrNPuCbBz
upMn7CBcvYYy0nzFxOj1qr1grI4G/Ul1cdtVKRtCqHHnNomKqX5L5Aas17n5PpPXI73x1GyHwclE
o4yWjbYJGPeD3EZsIBARPxJ+arAODch4R0DC0SSAmqC5xHIPf0tgentzLHNx2qtm5C49oloaPnzw
OqloVWXeJXEHQWoyv0jukQaH/mWWG9S7JwTwpRP0N4WoTPebdIGHgwUz3WLlNdWxGnRWylMbgW4m
0MrZ2PxdDAQvUb1mF32aH/+7gd676uVduEgcK9dJlVizmFZEmiFjVSKNVJwBOwjCakPcl87OcUsq
5qHb9BnOfkffCKLUxph+AupmFTfW1+nCnsVcp1fvoDRTS8QlrrFoyitYvUvkhqDFZjC4cvsMG4wl
3hlhiI+5WNX1XPRq6TzeQ6/bo1UYGatc4Gb8UdrAGDsx0bYnez3QtabnJXmkRWMCfSxEdn+OVgDr
x2PHiQQQbK6MeS83rLah5d6MdbF2mgVqekIMKn2KOvSJAJOz2JfsafEVsb30CqeKOCjhLoJO6XTL
RioGg04xOhgdptiMUDkzlwGATgABCj2pbXA49sV2yg1iirXauFYsNklx5bc2wtyG8JwkLbehRrMi
Xxjy8yyI9dFGpdxjNIyae/rbR+Qw/QmrGFjHbaQ7m1vOJbzfFsF+E5drr8CHYFl+r51P5ydwvvYd
spgWNiHno7QwvDZYKmLCD8VN6tFcgZInIUlM37UOBxPLq1tFkvwEMKAuT615klrJ0Qva3hLGGB3h
CDu0KZm4fBWxfbF9PjUWfIiYA4j/Kx9fDUd4Y0R3DTd2owMUCoJD1vYrKzC7PsYpc+oQM2m+DEhb
pzIFfKMwW42BrsZE9I5vLdvNUDTo3iqHYpQtnULEk2A53GIsemeajHNm1E9Aiqy4nDZZym9Lc5SD
itx7l2+rOeTbI1c7y0vmYqSPlThbkFAnIyg607HJpexFiQWwA/VwOmbAJM4Ly39adSrvHRKCZu8o
WLkQfoojCAICuNmpBUwy1iq8V2Z/DBJcOHOMaDhDhK/taO7S5YPdXNTvO2vyh+8cZQr2bg+zpgNM
7tQsBvpXeYx41lJXwR2smGtk9MmP9fxpMe6eNJf3swI/GcSXYka5I5c4YwT3y1FOMrF+Utl2JUcf
jK+wCujqLn/0DpK9ITYbJRkWew4kmsgiav90DhFUQyjjUIVLl78t/KelxH+hDHDIRTqogNH6XpzV
wnzMRezOQeRILinzCzIn2jF0pxH/GGPtZe/lYFC66VjXbCCG8u7DO7Z+8M9c7yP5O8mLYN+Q6cBr
Yww1WgdO+4evOsZXw2NjfURi2vLaYlCbP/6ETmYjZAzhkrAxqFxUFWlVws8laqDXhxWNtiIE1jVY
kTD+t/3uLyKvbqDWQNn5qVyGq9PxC16kIjcrf2bciCCntoN5uMxE/4ia+NzfVCJYKbzOBqdU6dye
dY9uv5mEhPFUthtMWVTzhvzczYrbnDjlRD1gMbcheUlrdS2D1Uee1zCgRCa+PHrJAiSSPcqaBjWW
FrnVPwy9Eth1xoFffVEWGTvXFPMRhA+Iv2hyWoiM57NEX3Dn51OG5ACDGO0+aBr9kQ7Zx2oGpoTV
NvHjjDxT2bSMh7BOkQ8dBdNGODSUPQfn/KwiMT+rN3pSkrTOZ1TWtAzt0dlzx2PkMP375CMqEsKV
rad9tFjN0M3X8x4ox7bxOAcOVjrhrs+pB9k8IGwgwoaDpR38ytuBZO44IMR/1yww6su9BnbCstWj
jdfziGk8vZivaZsy29JIwiLdQzHZQuJdlPdSThTHjD9WyuvAf61sFV5g5lwE157bG6718QRkeiLA
Te/9C7abq+gNlVxYeYVUs9vBmx5sGrU21m2f2gRRXyHEbUgcmjOUkF9KATTL4V1H7YWyKGYdELb2
ClPQ3HLdCObi+PJsVhEM0yDuRyAmjcjMaKpWCXl8oflZCeHPt0dMzk3gqc8/C956Yj76zdBNZnj0
8fhgm0uZhQs5G6IguQ/fpePSNJM3GzAzCGR6iIUl2E7V8qbGTVEwMSox6zdAyPegwXQdcUx2iZaa
/zQv9gRkiucleOE6awCMSO+6KHkR8XJiSwtTepoxDBHmjzrWMX2sfdY0Ajq2lSdC0EyY5Dt/3Agy
IX873cjl8X7YKKBvEGdY2ZpfCsD+w4dFSY5L6FN9KWjvQvEDgfPEqzEz17JaIV3pJW5mVFioKnAE
EXOZ7Sfq5mMReM0oYi02NzY0UHjDuu0Nh8VRIvdg00MgyrFhW+jslLAvraGgI1xf3xqLY40emBes
Nw/BwqJPTevT4E3/+4vbX4ZlMYQOi8GMLH4eyM7Dxnw0t+0XMeCkefUCLmJDdGnIb7sg5d35OH1/
YiBOPclf03LOa+xyeBw9Y0rB6oZHboU8I/9nRthTrptd0/+D7e6Ws63M2QTNYpc3h6V8Fqt/npmo
wjuumQF6LwhU/zZL1tZogsgNjJTVJROhKhGOEEmyC8o9Gs41p8/NLzrBnoYWbStxwL9DS/CpUhV5
eWDZiLd271cZ5qgcqbx8gfJOAxyT8XvGahW/k5KkiOGyvHIzU8DYc3mkHI7h8Jcx6Qe+cUwE9bSj
3SM6bJIsUMNDKZG91oPUNEDGUkCtRxPMChlLLTPoFeyt4BGi2vxXq/7ItpgvrBSQvShKx/ggP2DS
u2wH8Xlr2sMvKG9hjnnCyCXp3hY6sq9k5YtvxmMnus/tlRw5bZFdlJaPtL5Rw8LIPSKnZOSc7Bd0
2P69aWPg1kQJfw45ECoKVfPNl7hvCNzMsEBP/CfygpGV3Tseya26UdJHLeWRStHxOk2y1FbUacX7
W23hTes4RCqiBcAaKQUHwFx+FlT2aDGn2AmCOYaCxalrN1LAya6YhZ342N9yOCic3TNH4rfXvk+g
whQzB743sm2rhCykXtk2wtXPRLImmSl5JHap3kOV65kciDXQCfBO3oTA2TcsUJWCwTfqmSJXpMsA
UWMdFGFpb3O+pUxBua0m8nBCuIic3lAHAiN8VQcOiznUWLQ41D+Wo/AxINEeqP6OqH30XwPIWVGc
zyBOlrgOmlihvfmLgHDvu9mzcFxw/c7Cse6uI05n4run5b1ZCm39opvO4KYBhygGbdlhbbQJ8FqA
Ym04ZpMGbvRENnxtJaxHTdwPe56wCt+YSOC+PIxVgH8/S5BsKVG/J83oqPAeNjT0N23E4OoH3/Xf
76KMVflEsys8m00Ku1t3Cm9iInVJqgZotlR4ir6mIGcKu8Aw+7oXH5TBprVybFaf1zFe9wKc3JO2
Wlfoy1zK7fBIRfEL9wPk81f6C98DhSLpxOtHdUXIBgjqotcgwWQm22o639znVMw5K4HEmeYukhfL
EnuA0xolzNoKsteAEnLtkALhEIZBOap+9Ks9SY0+xZfSGunQ8V/pJL2oAiN0deCDxohuSzcD0nt9
b00yQiwyvxelU46mo9mTC1hC+mzNnz8YEDMY4si8qrxsYydVD5gUd2X0Uu16LhFVJzQ126LUv91/
Tz0TKYEsgAyzQ1pc4LDQ2YZpiXuLRPGj+EmQvAL5RTeQHYeLCn+cwawLEpFONYnqdR+jaMqbvVoV
LUFWG2lDIDJSCokKFEcnzVN4ZEWVbX48sjArFCf3R/E7QkKvKnEpxdrCsq7YuNPKy7GE5z3YrlMg
3LSzcooNcNsnTxHFcgd/B+E5kcQNWFP8gVVN/RAYeInfL2VxxgPlnqc/f/nquhMWrgLtlQbVvUiD
ApDdoZOe0nxbCM6eO+h/+m0O6I1nsSwSPYM7NsJ9RLPJ3877NByREOriJImaXDrjkjZgsDHe9vXl
qJ5eqFErF5ciI7kPSGCc77+pHoMzyINymOR3ljMjIW1Zi9GVLhoZqaTdmOWgPICZ1hrJbaVl4JGU
181fBzA4ea9KJZtXvbWQDyxz5E6JDLgyGF2B4HVpsEmSMrTsClyN6oO/0Nankc2FcF+a/ZWN0qqw
r32I1VfvPyphlSB+pdNkVtlHlj1YLEfhiAgJoBujmJyd8ovO76CZ0Da/maN6e3v2M7i7fuZftOKW
50tvUPboXYVbgn8vPEUF6BvvxTqAY1alHFL+Ry0eQH7Kpl1CcnMtUcah2O+lk4pHX0y71FCOvQ+I
dsygmYHgHZwuP/RG7+Mb0md0Pu9Di0c6FMPY+KsDQnOOJhpE6G5NSImKZrUFUGf0qkzXszhTyx7R
7ZR/zWjjy/uGjoWJ1iI/WrMWRsdLKbEbVkpVk2/yv/Kbuf2fJI/ebLDjWR6rr39SsOhaDL0uQwpy
pg/y+SBocU+tsp2nhwRC7DbtoexpSERtoPdN6c/peekolPgmPCLc6f4lsiLlPK+nL0+J80mvaMWA
gaVL/pSt04+DqIPS8XbqVKxCAByVsxkYjwUwwA3rILOiWZCqcQsru3+wvoQBDQVqWFERXcoCTjx8
MvoT0zYklLtavF3a92noxKIVWimHQg03+epncTzG07cfmDkavhldWPrqSz6t6uamuWWPhMLhF+YY
D2ftZj/tI6maOOImR4gD+SeBpkWNxEQeL07AEAhPfj9vuZ7safwSa+FQzJl2MRyUlSnqMFbsSCfY
KgJcyogIWEeZACIKPz04iioCDpMS9cXtMYQTqIdwvBkGnPPa5ZhZBDIvud+nAhZ8dgoLRI9vdY2h
zHj1e59o0sWZPUz+a08a4fXN6I7hAGhwxCHZ5kwOsWiRLvC2yZ8q/8+k3BQs6/mFy7Pf0+C9wNiB
XQhgpjnANyR1Teqi6p3Ic+LGrqnkDdcUYGgtOgSADQkjsSF94LGUBaS5SpAewK88yrvucfORUYen
cap9KY81ZxSnO0DlWHdi1+mfoN6+hKvR3yG/h+ls0ol31JyKiLlyM0bDXXEOiVHpA9FGOHXGjebm
W+t84mfwOP0B9Keobu3E9giRUjLpke9DyKqVJuv9l2m8PC8rgn648084sviRwXHg/qupJ5B0rZnw
TeUo6ANETERqwzSZS8qIM3DaAvbsbXYlZMzFgCBPLENoOF6XmkHGtQ+X6MCLni+VETctgdEWgr9h
NFFt02h6VSowYrh1p4kVobMxACne08/eG7srlEkgy9LaQAIlE7jO3RqJgIo4vy1dptymujBxMgGJ
Ix2CImtXzGQ7DAlA0l5CRQA9lc/C/e6TMnqv0XpRqZHxzLHxf2h3QtElCerlCuGTPXYP7b/YC16n
XVuMIgBJMzsStvG4lb60qYpZ4EeISML06y29tr8b3PFOUZJb2LMlHuWFUOUbAKIHOetc2nmotYKG
QqNXr/rMpDsw66oezy1FSeLvthwrsrxMzUH+TLhSywXoNC3vK8RvRbkwW+RDuS4tOuKjcmCS0m2U
/1iQqPxBffVeDAuFZrPMSCN8f1xUTQPl5vmT+TXfiBl6uLYtpYXsX/Bgp9HKMeu+jrFscPufLPSR
keLwdw1BweNOSDgMz1i4ylhAx4KZdGgLPTmIjd2IWXIRObQjbPmh8CJxQCOnjMWLZjDtinI0lBW2
1tVHdryfHz33tbbZ+2Zng7jYsms25wPWsdbkp8UBvCIKQqUBfvUDaeyE/zbvNvAOD+vU2xqmgQUM
MJe2A4WPvMMDPl8MnC0Yq1ca2ncwWMdVg/P0jQHQ5ZJPwfpQsFmlNAtcqmG3EqIKahXZkWr1Vqlx
WlgDyJ3t3HEt7V7y8rZ3DeIGFz6UUpXWt1mGr92XpTvDz3a2STTVZXeLzQaBqcJuyxVmZHTNwiE3
4LgvDHGRT/INdiepqz8h+2xVgJMZvi76Wilmfzeq7YJdiB+n53Tjj14VUYm+Wf8xcVYMW2KAVLaT
i8DWiyCLJfKbEhfg7Ytjanq4J7yxY9DaAlMgTaFtJkWsJwME6TRRe5Hhy9fcULZXwYkYVTnpoAwa
4Q3wBd1OuEHEaN+BmT4r6Hz0TEq9p4gBdfYUnkbt+gjRlG7abXKNmNmRAdFQjIK/Y870ZjeN0/w9
5yU++ahtc7UVMHMpqenoghEpeg5FLfqblbeJ46f0xX2HFtrh//TYHskFKqV0ZI0VFRYuG602Ia+8
dJ3p5Eag4txjPGZGTInFe6/GWNhP44QUjJ/HcRqaoTX8z093so/P/sdXjHoLEo/gu6c82UmF6vVh
gK4RAmL/uJqo/xNeryEp6Znv1p/hZO/sqx/ReNo0cZomf+IEdNwIpiqQiLaANT/ox1uyzvX1LWis
TMIyPAEXu0DmSufyCXG6cGf59m/kJhIhONfYfXiisB8ksQM1tT1hvUbQYte/eTsPu/FtdSN9ctUu
GKYd98tP4ia0dek+7SHK0vMM706H+kBOiSz3LOD8sWILfqJFecC+EZx8CHKG9wtDaW2ql0ZdJ933
DXQjzX0obgrEU/1tR9KoemHPa3RIpmcNCVwmF5tt9yNWIx9Vw/au7vNEoDY4m9u1ijf3wuSp03C9
NH+wferHa7mehlXMwbnYR+6fdzRUKdjZ7kGwvxL86spnQmUOFjbVrKMKdQj/HxScuMnos5XIwH72
ZIRvnLK9h34lkXaGt2wkHtpz6hD24U/RzdIwLWQoMDstkT1Hr9lYgcwMAunU9ATZjCM0kh0CcOmv
W3ZjW5wexvmThQKiR9HbM7kLBFSXywoHATnXtWV69ZZ+Rgx/I+hkXPzl0AdlBzX61ePOXaNLWbKe
BFri/Ymrhtc7hFYrESPhw2CWp+t+kP9A9jN9m2e8PmeETtudF6hWuwZv/vWqgoIb/bYrv1s0JTSv
FvRhbomnNWbe5m+80DQjvW3xhjNOux/A5q5kzDi7Fu+3CHobzgcMUMWPAkePFktaqeq7or+Xb+uM
aypJjJRpEcPgU0lnYSrtXixR1x9Ir9ojai8rYznwnBwT2O6wVXnbffK4rZgNUqDYhCf77uqN7j5k
RHgJ66h7XfjJmcWfYNrILm0NAXL3IwK0BzYGo5j7f1RuNLraQ2HasSVSRMYeSfvzsXftafj5pqBa
j1HHeO/oSaq6TIijqAyD4sGboLcAlqZYnEkgS8jhSs/SFU2DjTce/CVNqdzzwz+MQBTxYTSM1Ars
zNcfwDtiRHDS9R4PB18ffJ5CuzHCzpG8TJtFuL+2vEWIPBSHUSGnRHI2kNd5nbQguUw2rLOiwkGa
VbZqmPkNchR/uNYKHfsobLuBGXUOfi+Yb6TDT7uPUTu4dg2FBhFz8QR+7+T4Z4l54ac8ahW14gQL
eCcpOK66PckB0JED3QVIvaAmGAvaeQnXejL1FL3XaE2VW2X9CFluxGmDqKfxnGA741Z8UdDk++TO
ne05M5obIo/RGLbC19Yyb3/eUgac/ZIqd6Zw/+nBCPIFcZw+4qKJTEgw05mOkPGJV59Z1CADQ485
cTKYwt5Ugr12QWAPD+Qt9CNqSL31bTOM68m/kcGN1lTaUQn0Rgkd3Ai22658Fu3HsAY21JR+D6GC
PhAW6e/UVRVXCQePr5Ytto/XypeBjgzBqcaXrSGVqPTCpODt3o8icawRZBHbvLJ1+KnsMjIbCCvi
zpsrhQJ3zxiY2kSGNFrR5IGDBZJXUSesKCJhU+eSpRbvQQwymBSZo+7a+sEZCYPd/tZCBpA/g0Zc
W1490JYx9Uv+t4wBgiZxXP1ij8/vc/N6JZREaXcc+g6IT3wsl6efFXOKB/8wvyVmRVNqh3pKudvC
rLRbANB8gAMtaokJnkIVuk50Ml5VdU9OJqtAgCLfTbmZlX2SWRvKnx6INwLzJJmJLGcmGqVgjWnF
t+XAtNhylKbRqnkUr7oyNQDk3W01gZf8jGg0SH1JCxh5PYRtw+mNxQUf1jdkox/npCEcQhE83aou
mdJ9jzRMcRy/oSJehnJMB26i5oEC8QOw5hcX362GmFgRCsY9Wlr+KH0EYDqXhL8xOMu+dj3SYY4C
ykTWkpZ9l/NFWr7OA8BhS0jkx0eyBuGwM0Kgvz5f4T+Ek4TzUQhKxKs2h2jYfF4NXqBSKx/jSfO5
V4wt3TSH5319AlhH361++gAUtwXTXTXinym/x/UjUjrtl9fjVFRF6WZWNGdZyjC6RNPINL0YfzTs
AX5xvwk5EBPKwYlsyIdHYiNtbU/5BLVhH/7Ue5iG/10ke62NaiPVENSodpkGWHRFKJIASEXhm6Ft
tXkrS4jB/Ch+OGZHE5ScmGiuPVq0QFwLFDx0HXrBNUgPv++YhBxcVzhipAijDfzbTWJJbqHORKCw
uf0F6qjDVGZOvSVxZ5DRa755NuiI8BPqOgM9r0x9isi4kknVRM++jbxSCSGh9YaxstJpVzNjrVK/
Pu3XGht5fvXyl1DSTehYQIC0kGzJg6UwmtUDQZHLucf6RIvzX98levbJo7vVP3LoOY2rE20DcTYP
lyQdAfljQt4HkT3sxS45c2eRhlKmjCwAPHlImCGqb+lx8Wz46YzNAblsPku3pORcu6q5jdxqz9zU
OqhALPzjkSGeueYeAVtwpnUkT6mslBkvllVgA3oxwCJBj1xW9HhVHgtScXv0TVr3K+RQ2rdGtulo
tKfoIhG70ihnwqTDFTP6x4QYnuyhi3HCh+jPAGFsNG50NZrcqfGuz1nuSRTlhPO+spjUmFW9LWtK
0ZOFkj29ip7lIXul/MvCY/99zWVMYSvkOYBwzEj2QOaeAl8ENJEzdfFeGTAF/MEKRLtRWEFbG4vA
f4dYCOFEQluUxowL7tvIjK+AX0m0zYVYUrzHQ09tkz8TSGrZWQftWNsRZYRnShlHOuSd1Cf0KZqJ
Y/qg5wXcXCIN1hn5dz+Sddjc1t9UIsWiO4Wh8YJRXm0XrrzP3af2livdauJf6W4JNtu15fWvIQsx
7jgBz4kPpw8jzalSfMpWsKBYYd4yzUQdyFKmH3/seHbE4iBzHhOnlSYrlYtUQw8hcHVQZHKqsat/
5AhgYnIhc/k6Nk1dflm3xbiFaGZXaG0vArue5PHwb8a7ryMYk1EB+CS2pMr1rD7sJvSCvWYJUjBC
0TFWWhHcfRH6/MZNP5Qgn/XQqIxEUDno1g4Et+QyB3GyKm8kTyZzu6XGyVvs8BylJ/cUIbq2pudy
KtsKDQnhw9FwmLkVpC8o8TphsSK0qY0BmKYPnHwZLt94n4NebxKLw5DZikt5r4ZvByTr5POwhDVS
Zh6JBT0QYrUSr6r0BENnZ/nT6Dk6Sf56AZlWUEIieNKMNIIungN95GarExc/prUO7ITUolbLssmf
TPa5mwHX7mszlRCXO40b20odl+fRAavcV/hIH+oW4YZ26wUOhGymVTW1LxE9qG5JgVQOm6eTXys4
n6KEYu+8MJZzf0w028kryyg9GsmJZduIL7p0aSZ9t1b4EXBVi4eb7pZ/fgnhuIvEnNGkoAnO/rWO
5G6uTfszOGKB7jNTV/o6kailLv35TwGCBg/KwRk3z9GXojfGYdyEXYd7/Q2g/P2jEsh32zauRIkY
dI6xAJe1SORnY/lSGfNJd+C2oY3b0+4tmUYWbnqjCty3zT2qNDMEpNxggVL+iWlV+FbJ6/ys68C6
OliO38KPX5WdJvh/Xn0c5ObPjT1VvzUO2SEWF+aMeHFoiYIvqp1Q571GqTTuV/Efp/iU6Y54Uetm
pVe9tr/CqFnbNG+DbkFdSVON6eVSizKnDegJDmIYPXABVXIL7oYR97S0mxvcE3FsdzH1PZ1uwZHq
P0Wivyp0QMjT57CgBRqzUKYyGGCkve8hecJ8IinMIQDLZVebaZtyIM0+qlAZv8RNFDXHj+nw0Kxw
y6ULgNmWsnKgyjK5amBiJfT36zBujaql3MAdbWHiPtxYDlI3GMQm4KEBm07fxpKLyOA9Kn2phy2m
YH4BV5KGz+KbhX1mRUHJcFJ0dimfR8WPq/YeDNZMfIT6Ou/v3m2N+slQGogMuMTFDhqGrcwUKXtk
UyV9UNRZ5Ye9UVWGxqKMh4Y8TALNxzA80HENe1ah8xkJNmx+WoV8EBvlax7hvrxDr/AhVB9Oxy+Z
EDG2nuhqnerWoM+kROP6lek7TeqBNxnQO3j3YgunBK5/u9U0eg/Kgh1IPnhc96RrtEzHsva5hnR4
ekxL43wvH8LvS8k7P06+DWOmDE50zyAHAEryu3V8WStoa0t1BO5MXQpajjvgaSz4MWRZNMt4iO4F
wfF3oylLQig6XE/M4Zhsky0AuXmaLpbsHRBPzlbwL/hrwOXEX107WRlymVJShTP7J4X3pD/K1coG
oAvcV4gPPUmgrY1VmNTBYVX1QFqcoitVdju1GTUsz+ltFZ8Al+44/UBSQTgk/cXHNoY1iEp+/0Qf
IbDNO1vlFU/6aH+0eXtknI/Kvx8sHHK3kwQJ9AWFeP3nZdpguqy0PUEzfPMfkifRnVH4NqjZZeQL
ofP6raFnn/ALWpSlF4D6Dj7MPAVeF6FWBluMRyoug5n3zTG2MFrOY5ZxF8R71rv90IE4m+Z810Sn
w+NUf3kX6Gt2G3WGKWvER7oYBpQSTeJlGNTOgUzA8Uz36VFOEzWY/X9csd4YhY+a/Lb4fwDx2BLj
/sGwaqfvnmVjMt4giYVWityjg/LBRjLqat5ftB72N+r5sOlCRzz5WUwMM+6X669+eCGzdrrG4sEA
vOAGExvpRGm3NqtbI3G0S2aI+67FjZgI5zHDjZ4n6ttIGWfV6LaJebY+0rt5Xh3rFOcugn50v+LI
z6Y5PA81doXYnTmuJ6HjTsEhtgTZa2Qboh9m4yYcJ+5K3PlfJCe2l9toAexDC5W1PDm9ZyYKkEgm
cleY1UPGVnEqwaXI7JyPQ7LBObOpgdhsHTHwrq1FUFt/wtGZgsEF+QrEbY3dS96pVJ2Ysr9NF1iR
XpqcnTo2J4RdYXN0QWTepInWQcERt+GTXFyaAFH96Bj+oFX5egPXi/P4QJIX9ERcUaw6mm/H9d3F
6bk9GCITzqmxhRa9Zij1FFje/ViZq/H2c2E+r76JWOHsRF/j35VCm7YbESoGT5BRuAmDABiTLxyA
5Rfzw0nlJo/e82FSmf6OyWteozua/C+ws8eU1QxotK8Ys+v28JhHMb7oMFx6ErisGVzCVAFcyW1n
/M9S+/h9nkyz5qJmQkEteuOUPXZJukZuu7Iq4/CRZkAvaSiZR70yhZ4EhTJEtms5ZpVRtNfTPlgN
cIVyJwDzbhZbrII7d6izkvmS+x/h2BBHe+fIGE1TrHW9G/I4Km23EVGW49VqIOMl+oaLt+QBXBne
7DCaKDGJ5LBIzEq8hpOFYiyUnev8QaIH5NgOz62S8uTBgy+X0Blt/RA8U+84724btZyY5capFqPa
VR8SEFXlzDIKZoyCVIsK2JmC6TdrUMFtKDXYzyX8cgtfhBcANw2v69Zzp4vgRpHzEkhmJno/FCuT
3t70b4iiBJUy1GHDulC3x91khXuJJEAzc88v0u/kvwipgsbhyxqVnxGoHk2TwM+SNNgTvmB+/8t9
aWe7iiPktrpg65Vv5x4dr1nxsG625WZcB5GQbYPz6e5Ldz1hKDwobTHrb0nYqZ2aiN2wrej9lWRp
QhCDLgBSbJIb76SApdrJLY1O4KsnXEvGYGbveX/lbBcnW0JwuUCcz41NtOUL2gDrBc0I45FzlDmf
V7epvydph8m09Wo0vItqXe8ZbBCB1lt2snp252fHQcxFYFnF0AhWYecH82nB1JfHKThOQoLAuBwr
zLeCxTxinPJqywiBFPxl7QIz5JuMCz/5Z5Vy5cjDi8yeclvD+6VwOhTm6pOpueN2B5BeCkQ8r+we
YT/mSukjrur3y/3h/uIli0auCZl8gFe7oQyfPZWs5sp2GZ+4D+a4DvB0+8H/fBzaubmBLlvcHc2z
U5AMNkNRyEwYVkfXHddMySq6yTw/eRIf7fG9a3xUQUhKd4zmxK0UH0Y8nVqogCWx0wbod2g+4SL8
LB6Wcbsf60tM+crEfbRp5SvsVEW7ZzdlIw6C+18Z8UJ3VwYT6GKcwg3R3I4MppVzKg6mxMgjQxr0
SktP0XtpReZ3C2W1D7ZBljjBGXAdJuljfcSRVBVpoHNYaKqyhwlvDyxwq0rulcNgNExUG0x5Qv5Z
WhPNMmSYM/dyrjE8tIHLiExlvIbgUu/hX2Wx3CTcNNoeHRw50tyJP+nbVRAQ8ft55HWeAC4GlxNL
oDRa6c5SO0CsEFcv7CxZvw1/OQjWAzdLJXvZsg6TUM2Sa0ekXPFkDEVileZYijBYWYAr0ZB3Z5Ut
HiKYLhWFS2JKbj68bJvLNYsIVP9ieSDAXBKFAMSUeVULxXFuFumYKLlgpKZ06sBy8rU8uuG/AlEV
CEOdR71XLS0fV54wgWjagj0Lyp2umpWT+RV7lEAa7V/Ruo1BR4Ix9oQ6jjvAC4OLQBksrnu6/ljg
ADup89JSG7OK6KMhr1WcU0vfH5EU1ZuuO/hHyNisll+xlnmNY9eAhzexC4ZxnptGtRzakT0a5AdW
C8pJ04ImV4HE+qY5Q+DAQfYilPjboPRAHoVXoepamH1i2WZ7+Q8tJcZjyp7RllBm7UGH+8DrCfPR
kfku0P977/v/f1RwGDYdflE8ET2Dt5J+0unnMZLtF4T4csXKfbQ3N7EOtCNIYGp+FP3VWbNxIn58
dyXWnhy3vv+TFlC0yhay5rDi0FGFMxQm1xvBcmJYBAOKZepGQlXhEj+EWen+rOx5HBTKeccw7gMc
hoP6KvBmJlBVgBMjgtHXztPOl0KhSGSTpu0ukE8/xq5gSfJmNJvOJ40jXHCDyH0sNW/B4UCDIQa1
RT01Agf8s0gljKs2Q4LO/+BcGOHThLoUhL7u8hSQ1P8TWu3Et5U4ay1tCxMrKGROOGjz7FT6mz2q
YebqC8UgIPdLMd/iMJJptJPjq9Dg3sYTR3uP26+GwygagxB+uH4KomvjZaILYxlmBqHsUHyBCkK2
01mn2UNHvd2sHS+GhjLjlgM8tGO1i7FsScaCnAhmlplF1ptBzzuLbE49zZIQIh0BdHrxYL/fYg/N
94em35VDqdmOONCysWW/Eoke5HilsgMvLxpXlbFe7mSx0TNJ6yru2OFx/pQUOyEwakSteZvo8n3k
7UPNbXFzrNdXp4Rabm3VkXSg7636guElU2FThyDLx4K8sJ9gUlOru+QZe1y1GJk+v2BVJLss3M5R
buZwCm2b4MD8F0mm8r1HlBcF7Ljk9JfuuBPOW1OrOKlhJUU1RqqGnwTyru41644/uYnXUEtkuKjv
dctfJAu2gbhdEvkqF3v7a+XXXGtSr3MukBqTGXbAHr3AvMpm4xc8P9O4o8m6uJTGEZY041ohdZFy
yw8asZOktLw724ce5RJU8NKi4KhUBm45taKL9b/1UGSOeRa9UC9v9xwX9GxRIWqmtqWhQ3Ms84iK
EQbJQcKeGiJNi+fPfc04psBY7S04dubmxybgnqNKTWgqs4LYueSefVuejcRwuuqFYO5y7XF2beMr
XGHDMWbYAED7W5+HKr8ZKXWYnKWMZjFmsRiyDIG52pntcgrwGWQxA3vsmTzJzzPIMbgJ25I6nu7k
LFcm4olqzzAQnDL5/wkfLum3iV5sjfRnfqw+qgo6lD0l1MeHHIQR2hcWDURmrVskVXD/mKPF7wh5
LedwhPRuPyXPqApakrpAhQpvlONqZhrxRMRC5QyX+N4ieRQhfoHtV+TtJeDwmwhuuwhpaqZiUJk7
SfhiOM1rfBldIJpUnetNt3USKH74aDJUHmEF/8SOrcOI2Kabd68/YP8pOl6HVAgulfu3dAfYy0IJ
DBTCiAzW0txjrrHBV8orgFd2tHTF/o0JS6O3d4/tfkQ2e2MEDpogHkbtnHDtIA4iJ2fuJCFxR1vg
7V/ZYOqf9MFJdJbviixsY3ZmXEkggEM9llEmi4OkuCiZPVgjMl5cvJXgrdjV2iU4dGBAOI1HJQ2e
WRxIhq8yKFPVrlnfLlwnd6JjBbZhmfvG5bsUDmqlGK3/6wSGLP/rfsR6wtLksDq+E1dbDoZh7d8b
bUyVCbnHL8QUOB0qGIRyEQjQh+cG72ITsk5XRxObPeCACVnzoRsCfxiL3x9B+t0U4mQOjuHR67tv
0o9lD6SeXuxSHv9282LpWwFaD+8lT1ppn9LHtJnXWL5MI0YmvSAFBp+H93YdVlgkGthFnmYaMUFi
4UIOiawDlsNVRtoGMJKyP+1K4SGoAYo4olkGt2VPx5urN/a06Zlu1yPZ9rMMt2Q5fX9o5bZw17tg
Hu1eF1nHIGFwLm26VQxMLRivy9cf+gs5e+3+4WCWrzk2QCxo0Pq+Yc5aeZMNJfMTaEkxRcAc/wah
bWDdNl8qc5jJy8HrAM5cNtE22WIAN8L8mVzwYQbM+h/QObMQqOxv1Vdi9Jp7HFr+6boBlQ4Cw789
VtJINVCCU9scwomAy3CI7HUOFUxIe5go8/Z3FNeJ/F+EhYdA/E7+PdTqyf+SgkeCU6WAo1m+alBm
Xnz6CDbLl3BowjsXWkdSjzkWiC57s/1p7EQdXDT7MwVmk/pt/WfwDQD36bQSp5SkVkAQo1izBPie
/XoJ+NcG32RUZEtzJGMYM26Y+17EAvdXQqapagXZPQ1n9NHsXpxiq6cOiQoYkDOnqhwyyJyX/cij
ZmoU1rNd6xSv6nxD32wjSbfJmMZN8aISSEys9smiPDmVW66oJPrS4tDsa4tiqvA+ldnnS6G4nho9
ttFtmoudOaMuvpukUwFB4kom7Qm7B2WuAkCdE3+XsdrmsNuS9mMqEccm8BvTelEqrchJFpRZjPsV
mnhN8c81lVYvYY6UN3BYbWZdfOUWBKuhhrhRwSFhimJ1BlUyLZMSjI2mu27AsOiQL2BXybLnMe/H
KFcAodClXpTf6/UyOaDyoCHN5BUazzfmR1Rhiu28o3i1z+1eckvFrhv7EgzNIRFzyo9t4TB8zLWN
vRtUMXqxjYBMs6Wc6pxcASyrN0YJSmk+gf+HOBi+hJNVGisHGKyAfiO3w+fULxeDC1rssW2509bj
Y3I+ptwnQ8daA9T/aF+Eel2kpFCgBn1XP7IJ7fAT0PsI8XQtc8LEmUhPH6qXI+EnJnZEn/Gh+jr8
K5BU8pfccFTKAXtFk8S0yYB8nUtwH9JwDGZFQtR2uMK5BIsdM2h37ULJSgJ9P9ndXtRmYHt5OWoN
S+xW932w8j56IH/IozARaraS3JLh0mFOsk7LdCLlmmMyfVrgFUYNFwQ5e2f/rfiT4ZFrxEaMSEYx
zDJ5fjbQjysu98WZmjFJn3zhZjinhCsg5OzRi2XWP2CDrGcADntwly/Fm/nU2853CgZ90PTONwRV
K1UGyZGnVLptxsL02dLYk73Q2a3Z1EuiFKU9BfO8R+qYeeGet6BF46sql74bpwygQE31UG4gO/kp
ys0Ljj16Uk+8QMSefvCHRjhHtTbFrCFKqKaTBsBHqH4kiwphqAq5qXXEm52Pj3iObmQf9NAWKNDj
nxLnt4OyFxA+B8Fd9lcxP3bWVBSC5wI/zmElzqeWJjg7siuppH3Jc9BKf8bNg0fSvXH8PtQlqbr0
19hqhFu0dlXBNiJSW+Xp5pGZZPjO87DqHmnWIbsYus9refT//z7Ho1YVS+6kAIYDGsTWAd7zXpvR
dpFXMJMuHm50+jTUOcvqWdHrZT4obib5SdXSwBlUTjKUWgEKUUcBJgI+aiz8F8EiH0nenebfbHaN
/uQ4lZZjsh2bcMCHkgTknwXoKoVkXBh+/O5HjypzlQTH8UmGAWL6ucktSdeTMCiAseklYOQdoteZ
otLsvCEb8E0oiGJvV+g6tEVDKN5NWuQEErgABfjJcoVXjZdaBRwfPnZev9kbgM+fftT4iEQhzEJf
IiBE4z5JYsZKzRGpH6DwyAEFNPopj6ksxPF9P8WkiTy6iWgW0Mu9Y5H+xqHm/xlc9xTDZmfahFx5
fIR7RjjUqq0tnJU8V3jpSJpokpdtgvfyjmlhTutfx9IginykW5tDnk8kODYG7VZjbJnw1oKCRUj4
x2o/Evs9ec+O/Tt4BN3Gf0dfOQg6369gQd+mcy/gIWVN1WJFuBiiTqpbmlDv+zMBIBXlJtf3MGOf
X4bmVMEzVbDxIuG4wXmzrC8tUoH5g5xCANpg1Ye4Hl+SxSGv2iEENBXLHaz6HrvnAI0tNtOLLmWh
SScYZ7vaGiuUCwp23SW11YruGa8ceFQlztsnf6e6U3+F5XgGsQLRLvun8Y6JN0BMayfOqQlVAs5R
zE65RLr3j1QwKu4Ig1kKChZlyeUcxlI/7Y0wgCdb89fAdZorJrVRGToL6h6bridDzdxelFMQU3wr
ivMXCLnDGcWm5SSKRO4t/WSN1TqPLkQD/w6tMAuwfG2zKaXIvEHcmnG9DJeBprvxGY3SQWaMJV46
88LdDDBiblrCUM463wkBUJo4Rieoa6fv9+MKSeO3jOLVcUWtXMk35qwQDgUmb6X0yx7/kjT/wtf5
7jmMokAFQN18Wa/UX32ApgTTr2KKKJ+6T8bR1mKqka20v9dQad+QJ83xPso49ovaTryHzM9UDKgU
T8Ay6M5j9eEFF8loHx1BysBm8spMILP9OPF3BFk64CAnVm/pS3/HL6hbe82ADj7zlfsRD2ZE8Q41
/+d7veLfAsq4Q9yLy9ZrF9pwAiPMs8M0l7txbvES17d/HdN9cXDT0oafBzMyCjYI4FOf6rkrcmE1
VTe1+qB4kdg4McEj2xCp8ZJIHFOj7kyNzZ2p9ODTGGDd7cQXJ8ZRYrnORJLWEIIP/MOQ1MydcJwA
oI91lY7CmVtIuGiOipw/pnurr0R4nAJHSyv3RIu3jRNbo0Bt/SbdVNcS85kXavd195n0/UxH2Dyr
OQjPcXJgjF4kxwa8r/JSlYxkr2MCNzNwtP1uI1UBfoH6OyV7MU+UljF//QEH61qL13wbHkSwTrnq
ZDp9rXB/n974S5gOiFhghqL62ZV19Uooz3po/diYjtUCIUK9tMT70sWRlOol0UIQtRUwT9QJV1dL
6o+/C2rgR1wl8UL9ZOG7lJtCSsf17jWRMdWDpo7iCE34AY5O8uuSkHSP4rtiFIS4lOkbbCvO4CQq
jTvEvL8O4Ww77i0yrfVlu2RTP6u/5Zcc7w6zpaFj6g164siGVA5aav6I5mTBT5xfcgBNFGOCr3Yu
pIG3MbEbMz8Ucq8x/bfgH1PUeQN3LHZdIpSQ7jSAt516oWZiTuPQ2+7v1lmskYAWWzgxg1CJGN7m
dkxAGSRS7K0lMxPkSChqJ+Hb3SnFy9dk5A7Eiad1SwYXUjxAZ9QeR82l+gRjRr+hxGusg9wL56Bj
zjx+mWcv5GZr7LgL8jsJrQ/HcmbbB+bjVnRNACp5RMitKf8yekx4oqpz9bpma9VbWqwL4wi0xlNU
ZAPiWzlJl+igM9V6iuitcZgAxPtPrmdpe9I0jimSkruvJq4xyT7A0BjmXeR8hnqhIjBWpyCXGdIu
1xREtsBwAWedQbqBoEZIIGkobb/lZyilSRUAhQ4AS2SR6PuVhhzcbI9oP65eaCtz67XgevUiOZ7i
SokO7J4/tOOhQ0euXAVpu+ES8KOgZXFrO4g29uehAmXSvUR9fyYE9y9ZHx+uukxYModecHNqsPvn
adGLZ98eDM8eqL078s3mCI4k3dRsWW05WmamQfI2/jSsTqLLzSptwRgaiG9jhsM4/mo5M+StL2Rb
kl6+s5poth/J1SS7Uh0V5r3Qz27htxcZhC6UL11HrAjx3dS4dsTzbP3yMDZkW3UJY4ibCSltQLRs
pPSXQZcivoJxUPNICOBUz7NrdYyyJVL5CZzA3xC0Hky7jyn9hu0yGZuUoNhp0ou0cFwjg+SYXWA7
GucvMlA8g2FttAuB/2Nu6c6MGznCS8obWU5YZeFdQUdOQTPmm8t91bBnILWyjLvWa5X1vHoqlexH
XtjhXlycE0rQA+ZQKEy0Wxs5OMLygyxDAPn9Sqcay/N2zrespceHXBMXxnNtaV0tObt+iKTrHuWW
+yNfKNHMk3ICrt+nhBqMfzKUfX5AHt4AOIp3coR7mkibZ2pV38x5oWZwbBVEsMO3L11Dnhm4l/cg
NUK7K8AIQ5PY/NgtKM1l8SHJ+q8RD8MHqAxVdojbJAC8NzJwzx3sXTiyKFcnIzDWFBhf2zHxBFmI
PV5oT09TCTXlNyHlvi8JoC1QfeWaIQL6GcAFu29arE3JihH6+LzxzWG6LPNu80GwiWozHwSXi5Nb
JK2tE/5/dGezM/K5SsVs49uFxVY02uHPSsRk3devgNLA4jYioQntkwiAvycZ22w3YXbDgpeEQGY2
NVMRmtmztjE0caWY8K58OqajMFrEBinEu3RLRWPbFn7nhGjr6GUsmF1ummDh/H46+tyYKeZ2ktkD
aByA6tiMX6girHcSsTPJ+c4tw3SGVdtPxD52bPTp9HxAM+iB8tYwl3lnX4uzFJHwOr/ah3OAvCZG
PSLZnnhLTtnJ332OpD9CevHCcicrmBV1SdbfQJzsvzW0pOetQp/uGyVQF0l6u/N0tl/g1hyDMdK/
JY9ngn965oQ+GQ5o8vDPrEAevjdZyYHn9VeIzqNwC+1v0YX4nkGclZUDOOGBddzHDhp3C+Nyc7x9
PVUlAYyjeW4o1Iquli33XdGJTcrP415HAw+32LwR+6lC50oly1kTa8KVWATMHwsBBwUjkzoXckyf
32y7GFjGVfxLMhmSOFxihmB04pCMnae1wBszlL8jQnNSFC+0e83yJBgQTYlenkXQHwLHPLEweFUQ
7FR2tQQFFr+OU2un7pHfhqC/YU459+0pHPWGRamNxhh7yEClb0n0X3QMlAn+W5HgMF9MP16AHDc7
s7R/rsv9gtWsm2GqUGEPcdV8WY8uSADlOc1X6G0uD7MNDVBfx37nOYGrM9sobz3vHtWY3Nmrctlz
L9DDwcCmmfxBYSa+wQH5zQxiNsDrGtXTKSHQ1T2uqWGIoOtdZrZfzU/n3YR1xDf0z2jmspj1wJDY
xi5xGcL4vaEpMo+DOICcvzY6uTRc3plA94nqTTHorlBoNrKFfq5kMNQpDU0IE5nfLaSu74KQquf2
9sRwL2CHVtru2MTA8gvkqltMTPzfKpvfUguUj10xl9qvOHc3Via5DwJtTmoJoDn78H3jGotCLlgo
UYb12OUCmMpC/1cMjJ6YesWxskHO6rOP/WLOTdjxJGyPOLHYDB17rGU1Jimsktu9QlC5ekfQvoO6
nS37bhqc/bZzqpWAQtKj1bQyyPd7DPBtCk9yvf4ZMMf5wcO0WUQSqC9cAUdh26zphKZ21VyiEJmc
3yUAQCEdCAOG3TU2mWBHDwj1a3wcSUeTNF7rI7dZsHyowCmwQm0bmyW+oanZEfse9FyE+Zv/YcjL
aoYfVzgYf0S2r9bjhDH5tkMdxl3uxaN56vXkIk7Q7g3T/peXrfP+WFUd17H5qi6DUaKLbG730NUZ
pwzXQeRhCVVIRIQn7pFMoY+Zpkdi27q9K/it9AjPH8mg2Tvxtu56g1OaNvdpQMn5wf6DWHBMVzXB
ffoa2Rj1s3zBUeD/cvzG+QsV0YxBrR6P2YEaUODNuuxzZxQg5nDmVmzfL6rPc0/NZroIODyUu5/o
Sg6eN2svktmtjwoKcedq8IVAB+wZ433kI7vBtMN7rlNSR3B0bRW1C0bLdZzTBMATH8jWjiJwZGfS
+WSputZOvLZLfrpnnqcpOGLbdXvrinl4/3U+5jFvyCb1R1T1mPC2l1KY7FUTVSzPA3nukVbV+OuS
riHqXpwV0xzC98q5RxwOwQ2dEUykYi874KA/YHFjnmMtjqmKr3nX4N7Zu8aMATRHmaZ2P1Nw8aKC
TePrPpM43RMV5bF6FN5dxoKQGAbHagl2Hx5ZIFG+AO5rzvZ/HMRo+m7bpPQUYaExRSDpouG99MI3
2JAlDCksON9nD2MpLbN3iex0hhdc1VEb9DHUbiYQWh6vnNc8j8awB5Gh7wPaqFeIb/LDie1oXT5k
M8oUjH/eGG03zV+qOTgXExHD7aDFxAur/9y9a0zn1+e/FCI1F9NcGzRnq/Ci+hUMZGZJnYxvFvLH
wJNLHqbYZHXDYv1qTUxi8zVzUE920PZqGaERw/XSBjMG5qKbvyg7lvRJ0Yh1gafuhQnixPEimhRz
9cSaIxP1TdF6ykOCYlT4Vc4ea+4KHYp2ddSYZjduJqED7q70e7iD9S8htxofTt2gdKlKVdS77kzq
Vi5+bWfuYyZ5qsl4hLMpwQFT24vIMKMtQqsbilBzrGMOYSn1S1OOsJCPNy+NdOvfBlIiCMqsoX4C
aSi0hXG3ndu73/F+S6uw2J604vxAHJzAEnsefTD2sK+pIXrM8IVnonjjV7kstInJd0ngPKjB1A4S
tZGUJytekMzg/z+8c0lfBPgongmejZx3T98Fp5z8CDa8DKIiel/Z6qn6N6wNMS6YQmNOhpTX7Qve
NtY7Dqj4d7PHKKgvM5EfsIDmgAZs2Y2vYMxhOut48kRvJPDfhYdMuTgDEw640djFVkCys2ppWO97
8/G/yDK6hJPIFh0/LdvlJb+Twopi37UPVgS94TZs2sJv3aHHE0AQN8TXhLqL+o1sM4ySkZJzRt9k
HES+fair+vNUQhnfQ7OAyhk59F0w9rKNnm+PqrAl5Am2c0c4NH8zVknPA8mVc6GX7bxYBG5nMvY6
NjtTiDJrBmETJMcVyc9O6i1plHm3BZ/J+1jGcaGlFAHLyjX7cyazgFvigHT/DYpSpF9s2dm/6cy2
fvWrJgIjH3AnKicp/4N46Oe1279Z+QUNgOKDNG9I+paxa0Fxrh9hqRZBV3xyGs8Z087VdZC+m++5
4aISKtQFgMLFdCOPA75XTXx8jCHKTCrNCL72K7jHwTv9WXde0mCFpzMPJaoXf7r+WqAz72nfvfCE
knfmMLFm87/oElhBrRxoNeI+lgNx9TF9v33bIWrLZGmGpu6yiS//Nvk2cR+UdELC9E3MNkUVdwld
v5CL24A8WsPyDO+akrltl8K8GHRqr2Dn8CL5+jkOTcpOFbJtqswXA7CPdSm8VYTPAe/A7h2XHieV
Q4+xGek2mX6sws2AFfgJhRFAZP1lqefbHtKK7pjzxeKj1V3qOD5NUMfpaF5Hh2QyAJ2XyL3KRc35
mMDOsiXDkfDJxe8OHqo4gSuedEoJAIQJQp86ftcF+ELIdnpYhLIo1n2I3ewShzOJL/cw8dR9uo9u
Bs/2qsmrBcrf83m9fCSbMWNAIjWzfBralq4FRqg//xwbkaal8b9zUswtLXVfqHd5vLZaSEnu6Ssi
swiwvTVpqhMklD726fJF0oU0g7aku/oeaeoXSKy3bdfuUSqJa9+WudySZDY7DA5rK78gGbp7RsCR
Q0GXmJdywETVW6mxi/J1lQtvPOo7g29PT35Qs53YZPyakNbUgWkcjAzjzQX8c5NOtB3DOUDnaThl
crx+a08JsViSmDcQppO62aKYK8xWu9k/6OLs1gv3t83tY2OuFTqqRchdlQchk3kjwZN7htDWoCbg
fU+8Q3wEpxNJzQzXH6wXBaXkm3c2aQrxQo89XyZPj06ZXHFK+m5Tc0uZd7hF+ekPBy8TEFFDwwSc
Wfj1PGuL3PG6R41gqtHwDMxKpdXX1w4m81PT2b7EtlsioCb2daxbM4Yycbt3RbsvogmenJWt1+8K
NH8KuM7Qve4joWaMHyqIsxyfuc+6DHB/D0NjldY16xKcGHhrFaFiKsPRvhhTetCfsYIsxPK2O4ZK
yTQxdXC4ZEg86mgxPxcIVSZq3Xa8C9G1C7DvtQBg0a5kFkntQCYuZGAEWGtIQIdJYX0aJJUNzHX7
PPd3XsURsX560+HKOkNBXLKx7jjaBWCDWLR8ioBTK2ZXEhVK2E1V/zSBynMJnIf4HLdMaVCwePrp
7uWy/amlTx91rMLaA61vUjnoIgIl2lfYllNpmJ4fb/3o6Zl1+r0PuwvT4IFkQ5CUUD2W8nGQOGXM
O7eF8xmFmoH2jC/uJyc4GrEKpFYx7auZgTe84l1i+VMDjCF8Ls2mX12M2UeNO5Dnpzp8ZDrTJLZa
W4SuozjZDY12W5DUzuuHF+Orc1lwT5QNVUgjQl0lcCP+UP0FHz+Qv19otRlhu4daGwaOimbqlGYT
vRxYqcimuOBK0JE1El7kzeNxdQIkW/ha9fa6dWi3FHU+0+oWy+QyYoYfMN3SKXGrLARpSuPXSpAg
sf2lejGvGTq2pQCsvmmn3ujm+LHBm0uCCIf9xq+Q6nYJZ44umxsA4ZMqflbSRd8N1UAM+P4tC+vD
szpY2mtTrISrYf6yEcoDKiUcaVbe1omL376AjBHS+TBT7UaEdY+9OyRBmaMEckMuildx7hW9WTiJ
Yxi8Ams1zABA6Um7j1MxcggqJVlI1/k30YrdhnY6Gjsw2h+Kc59EjmnY+Ys/ZaDTPlqw5qN1IFLZ
TMI0KPoygNHoXqeDV2xVJjyRaqPi3BKrbcCan0cpAotJGO+iA5SLftdkN5kphB89PYM6rZ3jLmXv
jpFHS3YNBRKrtyFfzJ+Nu972Dl0GrXVxEKzLLKqyGU1cStoQAflPuTg04MzYMpx5DzXDBpI13SSh
LZuM+aOW97WYAeRUYia1ksc4nMTLjUoQtYbnxM+T7XOczW0BOzKG/TdqcuvoodDfPejEHL1QgYGt
pxat/++bTUv+jbzE1AFCk6wue0k+kSrqGf2IleZG/GdxC9Hx+KcLVL3Lg30HKlFoBlqU71t7Tlpy
r28rjZpBadK15S9Y2C8+X0Ye0XUX5t5AFXiD03EPWUT6VaxKsGGEgchYP9iFU2pQbl0dE0924Wcy
kf2SeessL42PRMWfCgt4RgHQLtM5QyIQK18WHFWSttNLWWv0/aIBBjWTDbdrBuxrLPFV2JcccsYr
OOOig45HU38gNtkKZlBCNogFSYKyEsXUFx8xSohvohpwQwSoxaB6qTWjiXrZDQN6v+tvhmv/rRwQ
2my62yrz3ir9nNDnBSQWhoGdBsxZxH+GO63Qqb3m8y+4uGNDfjKV9GWTlmhTsP2mjU8wR7maMyOy
GJM4TeV4a+X6uY2KINMLD7bkaFd1P+zpUcHr8BqeJg/DyWk5/MyNsomyCrjU02+yQOmv5dLwVWxc
tzwnjL3hJHULdMx5DRODn2B1IK5s5zkwkWl4HWxx8h4VzAJ1/tHxO9/fVUqB1kDYnoAw8VQqIrX/
/iaMc+tYUuQlEgSuVW76wCZGS08gkB5P8/xhKqslzLFgQIxVdS/B96OOheAkE6xtV655li5faIKb
aeghgQRgrc+Oxn5kOnRB66NYw/OOsA1NlDFTvaXNsMYMQuEDqdpHQNfcVA6GzL9cSdJZrRWWx1Xn
cZpXuPHu0Ff8pL45w8jHGtduOq760hrAfvonkwjdlOVxR3aPBIulovKfk8ELjb0b7TDjEUViMu06
zRJ0ss3bp6Xc4swQZWg0zvHDpDW/R7+D3MxUBTRcBOVNI7+2WxxL3FPDPrfCMhVKUG+b1Nw0qxTs
gD8TCMJjK3/YcQhXjJIOxewypv26V2Eb28LbIpC+r8IAi9p7T5mFBw44/ig68JvhSY/ZhO8zBC8K
XxGHvaSU1IcOEJftwNp6a6n2JvLtxpMJU5+lcjIOzYdmw+bxkKxyIXcHGN7suaNTGwZJmYCIBWXr
JPoBFDpP8QSatMeGXbJaARn3qSDXS+E9bSUAhqR9gE7ttHf3aJ753IMC1ngDeDH37ntTLd8jqCA1
gYEfl5NtyMD3IG+6Nx0tUygmN+hFe07RhUjKZjvM2Y61Ky80lu2Q3dOccxMWlWIyzHxPrOJUJRUI
oUxHctiEpPerkp8V01NUKGGd4AW0nqtah8hdGPUTlTstws/rB3OfIEpgSf22QjpUXsebjS2lBCTv
O8yxZ47R5XU+PIfurgpz575IisWM7GNdOSKkH6b6Hx8+ZCjDehBg9c5peHjKr67Je/jo+3eIefgT
Y71R1Dal0oIEDciF3dMqbO+hmHtQKBfdDtLZ13yqH7QUxrt1DnEVtcV4Bg2drXgMtbfhXOjaB8P2
Zfk+CE4Z0lzFF4gMo2Ee2c+4NLb+pVDcNiKaiXNsYxms3vJnRuL+q6LaAZo3Ymynot3Z8BfCSvDM
bTZlLjYHYc6OQlIR4hlT3dJIkVAOI+xP/lix3A63Q/PD7aCrMQzaBLbKVGVwZ1cmHOo6Jon+N1Ob
6bsDUJ8xrsslSoRC4YjQ5luMLNpu3CJUaJ2kkAj0NGR2kPtdd0jiyhFLeEHQawKkCg8/HA9wmQsP
H2wbnQpb0H4zALH9gwwPR/dr07i+n0gf2+h20myXGwirPyDJmywYCZuM4tuEJVjyp2glsX8xIMU1
pD3Rjk5IWzi3to2/Lo6o+Jo57bF5sl6xF+pB5roPJV+n9ENDumGWz+5mvNOkZomSyYD4g7Yy1OhS
QuYiMMvaIDSt1BwVWS/tC/jHKAu3VwkBvI+pSCGAAwSMm/37Dq9DwvLZxylOF4oy7BjjKo7U9qYm
X9eYO/B+G0rhbQIIx5TZ5x5QTY2dFaOh2UpeGFqG0DMNOF2A8k/qGwo4EzGvotEGY0HW+UhZNHbk
JNT04qAbQWV80Qapf8Ktn77HIkojmX2IKtxOAPPF/jrq8qztSrE7KEbFXVdBxDyUBcBP6bA/nPjD
tjDaH0mXknmLgBMfKcR9g5hUdJ+g1yLMtTf3uzsFsJtYxpNwFijCWmuci66W8L1pI/AFU0IJtdk2
zxcJqGtJl0J0F06Q9Ai+B7+QB0cuiif5qJV6Sa6GJBqIdmJMaCSx8/wvoae0+ZYWUXgF9VnG8rxE
PFZWuyIAILNkogQY5zwfpHttNbRbFkZBZqyP81NVg/CU513Ef+5LpnXTzBau/myJhslwiC3X3hfL
PZs40EsTe/CKDxMRvwnlUC0SEzOzdTvQT6D2rK6lYuX8rLe0r3NUcV/QpPdWTtFklHtA2EmF2WWQ
HZOszZa6d7w6btYfcSJtD3tPUC+Ju+mR80rY1sQr+1BbioZKWomHe8DaRQXMwa7H5lkgAqukEDpR
KYlxhj+7YzcsZfngfte91tJUF7DTc6KzARKyBRBEri/QYi/HDG3CI/+o3X/yp3lIKXsVCR3twI0Y
dGfYOiZNL3Rf9dKWRBW7P/NH+OgiLj/pwRjTKCqdGvU/53Qh3+/kz5xvMHBU2dSg7OF9cvoWqtaD
7HxIGPzatnLbDJMd6Oiar0kvhOr1tBGFo+DwEkZGOVVP1KLPxHiMruI7nkH8LJwnd+4VNACS3edS
DxqGNboSF7u5SgBMUvHMHU4t0+QFAh+AtMCl6eTQwH9IUIT3dkhrVQ2PVJ1gJwOnICkyoge9EiwM
gPmJwaLMXN7vMLZoxd60XSS0jN8PFwi/BO0A7xQXCMX0HwEB2rkL8P7IMoq/aO68S1A3m2yus8p5
BLsDN7lwDbU9oP1ceaZuPAA+Rwutdz70GwTqQckHY2NrOlPDPg+THUEfl1G0zrBliifnYnAJSUr4
yNqPFURTkdBHTAAo17oZTzCOM1sNucUX/2Xfo6NBACJfJ2fB5GgNHxnZ3jMuxgCSx8RmYbfrMWbt
4GG0g4Cy6ATyzTfAvw/8EivFNBDnHkotPAF3B/Op/z1wnfYhCu3yVojJ2274C8UKpqEMnvGhIyof
d0PQ+FtiPGGO3fTPDdQDRuAPVrBRG9IXCXQcFtTZiDb5k3wcH/th4rUEWt1L8ONMyzArfQMEvwgj
6zhozlsmW34+L3HarpiWdj4Pw80IGrEg0hGVUbqaB/302cMDApHigkQv1ZdvJxF9P5LdN8HHNNvo
IYeINiSDh+LmLDTobJL7XY0C5fXFgdTc3vOypvOvZgZy13nJv/qIi3Zd16tQNbQefmrKE5yLQdng
fOTAxnANQDgpOLJIB6gNgjEQuntrKU8ptNENwi0jaUG89YeFKtpHaOnHe2UJv4r/O4gqZSP6W1kK
U86ebcK3WXiM6+Kvlr3rf1ROckPQKqibsqWvBo5j+AQOX7aUkucaWqvWlQt6YD/7AvSXEBk7az7a
tcy+BurF2KaYpXg+9I1CT099mFjQQ0mshinonkYUKVE97gF+RpDHXxmgG+R2N8XrhY09dVahvAo8
DUi9VwWaUf7uTH95i831zzB3Y48QOZP4hBh132HPCRCTNBIGwInih1a7wxj0WXqtRnwuGrsoSGha
ydCy+rsjYjzokI8DyxxiMBxrblU/Kad5kOJ6JfuRaQ/g35hJ/KFQ7Td2fl3u5RjLxBiPFavknKh1
YIRRC+8R+8xQ+3BJtUMWUXV7x6EvK3h8jmguZ2UmZF9lVjq1KQJtuD783+azZ1XW6jd26Q3goZYH
JtTx/IFgospqJCvcWCpZpXr0v/8urambkkXA9XoGjggOMkBcvhJzQXGwb8EkkwbLsha0RsvIJOA1
z4atc6hjHHDl0hv3xe1zgg2xuaUyXa4ODBQWG0Vt3MXxounJrfwqdLnK/gItf+G8h+/+W1XgkR27
OhjiXohidPNFOw6r3ZR0UJkC/zEaA7cIcnC5qGCxlE3XyK5F+chKBLWCqzG1xkX9TyfpmI8sytyJ
Vre1JoRrx73GST8d8/KR3jR/9ER75MbQr/qPQhGnuGntGK3gwpLo5zwufG+guy1xF6nIti75LGyH
86nSQ6X6GuVlLb6qg3EWF/qXlQTBjG+y5xSByzwlVsN/jTQYeRF11TIQzqvf+xM3CywTiNIseBn1
1AmV+pm41fjwSq9fpm1DJpoJEzhSZaEzq3meF8VSZz17yUIQ2ka0wxkbPi7KT5pv2NufQYDu9VN9
u5b0bh3JUfhvKeo+X2dEB5472uksekxDjpSvLiIKtIYwCHpLRBsrsCN9psGMvh0XOB6/MLq7bCwC
g7Jhkqg9odpSWDRc4PhxAiHzncPEhKeCSDO9IhTBEFooe20g9/icoeGmpa+8pBxeBUCmc3JYtJEM
7zLttGgoajv3Jy48pkp7RXthB0cvVhswo2purAlOr2yzVan/Wh5PJr8HD8Ld1ScC+GmcRktlvmr1
4hlsd2aZUl8G4QyFk1AtviCqugE6Yon4a/p+6BDunJnTSUQFSEpmH9KuvdUvunY/AMzvnsWcjtfY
svzON3kauffXqeDUHFaAWAok0dHsaqBNhgCGDQtQFlPdbCrOmCbkAD+XK+adzxSAdkrJAcqJ5vod
J6dKviKxJKDJc+dYetkINBIYaqmxJq0t4W1e29yVHJnhXavo5ABU59NszZ74ik9RYa5drVlDD4Ij
ivzbLhDqYU8BBRajRoveCuUJiIuzPJwWab4m+M8dJnUubr+96JFJNTGJFmirmRECBia4y1GL6RJ3
2A62Q0yQPFD/qT2uBoKgFQiof3uckFfNl+sXfvMuMdL70yFN4Iq2krwOjPPnbJpYog5pFWtqKmfA
4xlGo0fgYvwxS37+gZOqgOBNB+XG58e37rY0UnEWmE7gmAN+Xfm/AV5mMCVIZVKbe6IlWWd+FbdZ
glO/iK5ph1j3ihaizoYBTtGfCp6a5zgdsjP4K/9647ttTcPtFjqHAD0ftVXzNUj2IaTfafN4M4A8
hnTZJA3AzLq60lizdbUhNcYYZLcZmZa06Ba5MwQLnBQwGxODfch38+snyquI1N1mxsu0ekU0aDHN
0yYs70dW/QQt2Tp1z4KMVfPDFkbBrRVALvT0V3Pe60+fdff6uX0Azh3AP2GBSK92l0JgI6jsirE6
PpVGFyrJCbpIOTGKvWgOP4XoDvAsDxkvheOn9yYi72eXROlMWSdtVW6T/dIy1Ztds9DGbygUx3LA
sHoZY8cURyufh9IUao//rdeKLX+ThqUH2qDSDQFidLWsvPCuaTCRDJeLvr0jANadyceJy5U/Lnim
ssgTkvMXwAyFYpOV0iAtUtOSI+xwXY1vgA8W5U40O/iTj+I7WQlwaR0bhNR5G/Gh+aAvR4irh+ns
RZPtXDwKCCLPTbUxDyuXISX3/vxL9dB1+q6WctaRiOZh/3Gzz11NBR7AlphFq5VSruArVorF5uDA
KzVUzL4MYodgucvawUhnKUILlD+4Tz+/2l6I45CS+9rKPuflKwhTs3Ctr2vc4Gu756BgCmwcqQx3
puFMWyENw1vigwHN0D6fv6r2f+q6ANYSoU2iZeGnK6RpDD6GmaXJICUB5FXxJ6P47199VRU2ZgJJ
HFVl/DWf68/YJkjqVYOHKscWyG5KjwN5x3nBsXp+rmdxa6bQh7ND4HHpHJcGqKXtQdAuo+ook/+z
r8uLmVecZLMtivRa0woUmP19rxXpUnaeJswba9n0NjVYLxVOwHZ1rHrywEW4UtZKe/A/ahNhujZ9
FfWeK7CI70uPnPfJ2Hgvp4ylS73AE4cYXKJZ/GiUGf92NucgwsA2Tf2eZR805i4HSIkfPnVas8v2
+6SRf8SrVGxSIxSMBpyaiyR6QpZ4dBmJzBrKZsKc1axsID10ok5ZG78ybsiJVq99yQwlk3zpsJTV
Wo+uBIWggGFLI1aNcfwH2LhA+RcMdgBHw7OYpm7ba8kRUBbj54Ov3MbGP16lXj16IoxAFZsDIuDp
2/dpAlnbc13xMHHhTZK7Bi4nYcbgHNi/c//nsGgddJ2p7BAuOY48gBireisOlUO9cJIpFQNLS8wf
a57QFoPuFOBM6qwtUmLHm/3dVzxNeUwBFXrbEbRR4oqBYvj+ljsKFIkQ8CVy60lLg2z0EIyVNKLl
eCdjLtnOHogbUle+FYUaHpEbGTCMeH0xpedeTt4xCdNtJOhuX43yxRVBNLe1hAW9x61/gkC/oT5u
2MHB1dw8vvfsbi07PC9z/e8BDwGPDjuzd5j0DE1J4pxKJEnQi/rPe3jiCHgwNrHQM9vLltQjRxEb
IGIQFryekFuohPjji5moccqVMlHyFJujVTk3nQSoruQgfl5g89I3V3bV2OkOC963oIQc+6RjxT+F
w3MjDt2CLGFH6Z568DQwQvkQLEZOgllkm/CjnjAIYUqrP4a1to4wZSpbYpLLVg0bjHvhuhCJyV+p
tFfkI/1mhVwgpHZOagtefchY2p2XjyU2Sk5Po+LgG1EsxDR0oXPTMkhW89w+Op/XzvxSsSEildI4
Om8QeArg1kxAw3MYYSGt2nKK7KW3vUF5B3rBkqIP9pNEE9HqYbPCbaA+zM4xPH6HT2iBQ/OC4RNd
QEq+aWw4AXGEn9w77zlvCPDBGfywe3tcvZlykClGaujYbZycCFpaQhWRCyYVRXKRTp/KYyd704L3
tgzJYZMRasbbL0+/yTmSYsG6978/x+cqca7cLu1nZ5diNE6Hc26eLmscZplmLMSV/Qc2xFIDP5tz
Nz+ZQylCK6o9vM0jO6/3+/bwfdhU8gm1nkqobmdOH+YOaj1DyPjfL08zE/E29v4PdNIpz7iGZ4go
7s48B3BHwvVYjohfi3QrLvfGAJvH3oz1i5sq1nLCZ0+iBbFYl9zNedss/SrzdSy7a3mp0XdhTJDM
Jr/6V2VKTlobqDdLs/dt5Vx7VqgKYpI32UMS8VACvPprnuXhfo3gZ88PzgwrePTK3/leoDr2uP5C
Ph/hVDmFmhVzmeDv4Li3iqnLo8mirQylZ3GLzFeE0RGavEYa5axtF+GclUguB2ASTMpj78KgzmLT
1l5PkUaEoTqePCB0Q/qdiIN14Gbxt8CS4RyUcY5u6uuOQVdJ2ZXnnwoR57YfRHE5rwwXcpgctsPm
tKjM+V/pcud85p2y414/XGaDcvGUZ1cLGKIWGDUDSeTJJrDHRKacN/dbLy++8FSjsVmoNm6b+bfL
spY48JUK0JX2JZ7yW5rH4f8TJ6RrvAcCaSBFFaSnkJ8wG/7Phhz5scKmZ5KXa/6idXcqzOEZicgW
OcOON+XwfiF4btGFFy5Xj4hNuGuzs2C/gi1g3Dya2oq0yH+PRGecjr8WnlxMbacfecLhu5C3fGKu
1Nquf0DUqBLiWUk3r5pKI74T2F0uz/z0bcnaO8j9WT049CQgmtvGjvnfj00VFdyq7EDbFTWZIe67
7/qYNgWVBDzZkYRoX9b6e4dFsJwHLt8vAm0ndOjuHWELZHy/i6TdHz7lR4udlVKPYxz5TXvkVjIC
UY66pDg95TXHPbAIhyjcguOSIU1cAuEJka2oZHeOcathkoeCvsuW54AC10cVT57tXJee3N5lM1I/
Zfa7IZQnSpyIiQ3lI8QePM3kbPAhtM2eeozeaHha0ZSHEYstqjpW9s1uPMCkpRqHofKvUH+M6Ugs
aUKV3I8kzkHgjUIG2/CXQrVRJhW09YzCpqNsNMU3Dqo38SXLmaMfJT8mJ3O1ad7sLswIl7M9JAQJ
mn9FqJp2DYU/3eibQeZvBFV7kuxdFaK3YeWvqqZ4Fgeh+mtGL//qJtCQc53+eTuUDBIaP9H8Lev6
CzR9fu/RflIX+vPucQggDsDFHesAg/seVHqeNdrb+Kb/CGo6GhcTehcXpBKNJUMLfO16nrgt66Cu
V3Z2VWjPuJLTUJgtqhOxiS2/xhSumL8Wm+M9aM7mJ72ZNVxgfx+f94DW30MdHXLybEnnx0gfJw+n
7284X89VQUP7CY0ZUm7ST77ae8xjNPhMVRRihc2SnQZV61Eu14S6INXuxRAbcNuvt3B4WPncGyZM
snD48LKAxYO4pI7AED9sD6eby5UekO3qRax3Kzdk/8xk4rrPzo4KREIov+G1XbMgyK2R5JnDx2vw
41p7XdkvnNW85AcOAvrMFvp45gQJSyjMxBy3EQQ3SWFRq82+jymI3DBiX789uRlmUVd8oSxV0h87
mu5rBKzy7i2Um2LufJwQ9zCxgJAiqJTa4dM0ReZqjiWegB5tMSf2IlxiNtA5OXt1Py3M04QpMFLr
ynD++V8MwIYAf12eKwkqeoPT6kbQZvLLr1IqG8urHWJvOIC9o7kvIEnCvbHMxXcoYaj1xdV1PeT+
NR+eShyWnnfZxfsDkdj6JNOFK+q96Ak65DZqR+1CNjMKXebbnJHd7V2xdvQykhy6qES1EwcC+vhn
cjHmCUXFBPUROuXf2q94wlht0fQQoWRywn/c2b84C+NGm6PCTUKg+MjbS/8PaN/hjLK34XWvq5Rn
RNfAYFFKZ3FlguqZ+8r16mHHmElHZLDjjy+4khfZnIKxZitMR1SjxLwXvgDhvEr2YNuERJHK6fUi
wN8vcFzaX7F9YcMq3w+9CDn1zBejtHRHX5FwW1KmLoSXP5pbbaQ2pNtOSwbcatWRDO8Z5HZR+bO0
MhhMCHaFPJIVO3RogYJ9M/lylCf5CGLzCEeO2G0GwD3C+u8HAp+0t+GpvAo4MvICFc88dNXDBXNX
jck2gaNSar/r/6kevuaa/6txi5r4bRHWi1qoyeByG34H9Kq8J3JBtAMw2yXCAnkLUVxzvjn71ULK
kKBOTfU5p7Hach3VOfiiJRb7kaDkgQj/As7oe6IlsKcjuhMthdjWVptG1KdNbkBdJ7UcoqHuQUYy
e8dP+Q5iZujSp0d6q8wPkTMKU2bdAYJ58pO0s5J2SyfqZNe/WhH2mSZniboNMkgajyz22dZBoBiN
HHAru2lCRzML4I+dQknS/LxKau9o7v8g0mTEsppF+cp94DAOafyPi7WokBBsITCARHTZZ9uEcz23
5oYLoZq+kNvHr0gBZXV2JP9QnosSlYXNRxPOy7Mfj0K449OcSBiDh1lFbKgotxIShS1mEIgotfeX
RWSqgiAqth8q9nMIzKtMYPtAwx81Oy/nSo9no4XNHkL/v7ka5BL//RFlj0W0l6XBeu7yxNteUiYv
Dvri02ewpJhSZ0uy3AU09r+69VrU0lPbYHLhhc5xGnQDNWpcrzWPw58FvBkTbmn/TelqMSFOqlCb
UuL4h5M3bp3ZHlXHb9Li0YldHO21qmb4BccuPEEU8ft2ymQ2MToHOKuSr0BZ86MEi5HlfcX0/MCy
hZRM0HuYHM0R1arIoUz8ru/2zLLAJvEhKlrxlRHGLkKjPnzCOQhTOK5zZns9JV9lu3o83o47YJEj
XP3tzugpw53FggIlZzvBZQksI/YlTvJ2FUNZsA/KXd73WcuF6qa+DgVdBFuhqPSO8E8Mr+H52L83
vciq/k6m+4ZIFs/wNLNfBxrdrTAu1wRq7I3yqws4nJ0wJOaJCs4drFu3OHwDrkikQzcPUApbx5HT
UgtYOe2U+tszBibCQUqm4LkeIoCkvR8+0MOIxpueP8Q3Gt1DjfrMAJbA942NQ2tI0puX3twT4DIT
DXMSOrC2eLPDrp46O0Z408TnJnzjctkYHF4aVK83quxyts6jRugcUUUj1ocK0UfxB7j1Y1gW4q7D
jWeXNff5C4AWh4lJAGj8V+T7Bl6llzNMxp2euYGq0PdiCtDeThQtv9MDsm0HwWbLJOBynEQ0NF9U
narMklch+RKJMHUhLuqvx/iRJfOPXw3oOBeGeNFFmx+PdOWpFzuWi6csJb0a9HtdbkBlMk5IgcqX
IDEEMjrlnM9gE4rwJ+a/2neI+vKrNcGe6zT72pVrKeMQpPr7JifVmZTjpRSaBgtZvb8KB18rWHNK
YTIJllxBd2C6qjC9lG9k1fjjSMnKOyvlvc2TdEkL7FKni/F3JP2p9xXP/AM1YFuW/3a4AzVHUfK8
v2dmngsFhHhK1eosDsf/NJqlzBcDDEFS5tVGDfydQjCMTgfyMBXqEMVb2npUCoq4yNGOxzXFVxJU
U1eIcjBVNhmxOGlmXHiC8RLuRQNFIyDVauMxNZoVPOEBrTHKTuQrc/d3ES7nnhX148CHkUFupZLb
7g3lJNITAPSmBrkSjCxOS1HyoqoD+i3NgUl4tnV61CM8NlJRScqJFsz39aozVnN1jkjqAAUP7zCD
cp6ybEf7n/eekNEjjQXM1EMxdD7EtwV5zOW2Y3kQM+f1RhIZHIYmS4dbHK/UAi0G3LmvYFtN6eiM
nPA4fcM+GnFh1OiHLwPg4ymvcHZqBx+yOQlR2QjHbzISRX6C5G829HbrwpCMfS+IRsvJHuw6x65T
JG/ontqiXn3rBqASOBe0MaTvL+MS1CqEwByL3bBqNNgh5ZWPDHGi/eH/lvFtGLeCWnyZVzJHTLre
7TQF7Y3IzOQsffq4RbD60GkZSm21OTFrsV94LUHig+DhK/q5o+NBtYZITeHQ4F9DvLn9VRXVdCR+
zETxGaZLuQXua8lEt7KGhV7PNoKRUaklcZNQehw/Lhb2FcE7zt1CvfUFwxnaSfAMgK5poWhZ5liI
QeTA+MNWgyU5apFnaCdfFVJC/PzkZZBcnyMUNbnJwvGnCsOqHO32kyn2lGv+AmrDh+7OFWJiP5w0
C39Jah3N+uldbw+K52V9q5BA1al4DtRbjvvSx8gWnqMKhmhSbA+3GIvEEH/PK4hcjQu1jZVy+Tj/
ldVJb4eO0qvn9EEtE9KX7WiGOw87RZIR9jwosbtDpV0GAIB7nxhKd9VAlrdcX1yearBM7umCtdav
ZCPsGbIJ5tMVvO3Rzpbz943KNZoTn5IBh2wG2YLIkGWY1W2lpJu8Lay6K1rXEg2BgbmGnJfcbcCz
ys+H7EQzH/tzScK+8ZErkm4wRLu2GoQUhhcC3RTBu1a+z0M+PE+ZldTmnYPGFqE6rZFchs6bJiPb
4WIszfpIfzWhJbd0WlwVvYDKligA5T7sMO10uDkoCd0lxdkLbpqcD6tZq/dlPINAt1TXEClDhxNO
e4Z2Fmaze4fdT5PSyhaF2EbJSc/J1tEO6rtRKUnLGy2pLFuBWZ+V19IaALkFDDwkV+YLmWKv/3I8
ErpHdBpH+Uj36dFGLFQ+RLkdUlVIVadAlwmV2bUTXlJn7YzYW3MrDhf/qNfE1ER1h5MQWEK4HiqL
CNVLQgNvHp34m4/axekgJhzt5ous98rViqmvjYuhduLUjoJBGoXO8BCz5mRzIDDguORO3n8ZsSif
Q9dv3o5Yg4vKKtQEaQI3bj2ckHrT5kwlyWjpvALDH1L07eFubQniUVC27wPXPNhEIEA8ybRz+VA8
qCbxKRDt/f9s4WTe2QkqMilduRgv6xCnyTHhXFpGFS/Jl0Ows4wySqpbBWcQbCFAuGcFXvON13e5
Id9jHND081bzFK54kTC2ak9HOPryN6zfCR64+Q+A0IqVWsj9u1ODfe9zeR5QWTX4jwfCJP2ctaQR
VWylBOPs57WL8pgvOHdIuiXaB4iIA588K+YbNOYTIzeEVL/rjPyc//6lDykqn1oba0521vNek5bE
AcL3McfNpGWkEgrMt3bEeI6dV5WDwJXUaHlJAuj0Qk4YEk/S26LdMx9hHMblv/QLjQoWw332Iq8/
NlUGrdW5AAtNrZVce7A3P6QjSbaVBcBMq1Mhz6oG1L5FIM/qKrLQZ2FJAVFNssr1afoJojgH8FyT
h7Fks6VLEJq/1Px3rGnGOWq5rSbk0wI36N0YLKV1AlRXBifTF1q6lRVy205Jj9xmNzrBI6QLUJNa
lIM0LjVXr2996pSzBAo6hvTrJJcPVcNKKZ+6s3/7OtqY7p654OneDGfx2VLsCN029h1rU3ahmEQz
oHxgcXXtRD/htAtGZTiGpO/cZzGKzfeoauQV40ubtOk4joiqDAK/fENClsbYF3p3C9ZIS6kntGLP
Sge/mDnH3o0kFPW+8O4V5W8F6XGNUA4zbspa+kaLa+bWZ1jVR6kaTpniv1wP0q/vr5aMAFocYSME
hJRLqZPZMgFh0Q6vnBgdlAyu9qhd0ZOg0sAJ4xAQ6hgTDq6VxTRd5cv8dL2bnJTh5Zjou1cE2hy1
KXE6UzlA61uYcrLAOxx/zUep/Eu0cB8gxG09ju7jvk3XSn5NkuVx89ZV6EcWG/RMGTWTplDI7Kii
0xHaQr8YSQPEKV93aLdDpUNJtCikwGTjzkO3JZyGZPItvZRJ9+NMQXfhpkgcjuVS7Q/yv4JAHdUp
TzkdpSF3aklHfXw/ScnMNRD9iHY1rbFPYFbAVeQg+PBGEeJaB8GH4v6lM1CBMwM4k/RRkQ82THyB
1QyZzevFKimHlJCEk/a1R81qli0xdw2+VL36E86QdMuX+9AXEA6TQPqKVVgktk0oOfYMLHlJbV5V
tN4OgqQs+yHMk6sQ0nQt/Q9oRXd6rjeI22s3uB8s3WSahYxeAi/WVqBnj6KBzGlVSG4n+t9GneyT
/rSI8lCV8LGRGkPDFSYEsGPY//896h3DE3SiQ3j1bKc3N2jyewYrKJzlFo+7inE6w35Riv3GjowI
uzBHH/EP65NLDKT3Vrgtr5MZJgmCmv0fLBOv6EYMSg4fXhNwJklCJspKN9Addva6sHO8AKTzxbop
emFldVW0oxcOAaspB77r0DtAvDuNT24fPkN1zk5MSSDzuvMwy/OYpMEl3ojLCvcMtfYVWs/nqeQn
K75m7XDr1JKD489u8bD1wowLd9Qd53cqSvwSp0vaTETaXk0MjPxPOA8XSFI0zkL6A7e4S77To5ni
KZjSZijBDH59LkCehFsVkIqI9MYg4NdTgiTvlitNX967w5gWOSaEghkQ4pauVC2exhEaVLyAzDKf
Z+08FCZsucv+48ppM2TBHCfSHpiv22dn3KTZrE7ex3bKTbUjRR+LppFtz2BqNql1OOfKkt9Q1qHj
wQwverAgkRyvS7eugN4j1GNJnKfn7dfuq9myJIZmFm9TCJeK32wGnzw4B/RR9hwSwoFItjA+dZwf
2SKykZHQwS/Xg/p8cbFbs26Dm+uBKruhSMwFNQxZWgcVlv9X5z2rJE//393WxtZMhMCgomkbFOQE
3vfyGQImVSQ8TCz9yVbnB0rzZkn1RL42JCN0gyKX0eZ0KqxT5aKXeMQXEyDiMkQ8/8PZcD1KMinV
Rjc8sBDVVTCVjJXaAMDs9e8X3IHxBbMZg5X90/NJ1dxzJkMVeoyLjVFasPNGfC4fTt8iKAgjkxi+
nr+mlJbUWReFT2W7Nb7rpfSYpTJvv2xlvyyjk4WqHkhC+HhNVT/q8rzGu3AmbfUHukOC3kKvf5bz
t5A8/fQgyuzyAILGR3W3Y6fO0BLOQB+QmAPm4k73o46Y+dXXZEhVbLBRUG7v7wp9doPz7McRIX1I
UMSJen1q8lb2/18lkxQWN66KPeiqqpgd6XviafZpO1kkLs6bTSCHcLNpESvUEIm2fFZ/1ACe3DGL
MDLG78KYdHtvXDzPfKVYnmK2wdyU0V4D529mxqymHcujUjnCobyiwjd9WNnEkjUJBlJw6oSGlB/C
M6ApBifidDHNaY2pw5vYqG1E/g43kHfSHsmvXkEfclUIWnLL9nUYo1Sk5OCmOidUKZ1S4c2Jves9
ZL18rsQMcQqrFGQQEnAEdaOUv2JtDsZ0fIUHia4mrkYh3pPEYfrBai7LfzEnGkLnt/uORD2+7SX9
ecQO+FoO92rqo3nQ3MDzPQHUSO3twojvDL9Mn/rIIXWhZBaimyxdQkBmn6WjmQgDa0HPlEftyPkE
uJYInCsEi0fZczJ45eOj4LJkf96dWoQbDSRyEkx86H8rl30dvug9lnCyZShKAeA2aJSqwKKkvqq6
49ec6Bh76iRZXwKwoX+xqxRDP0KU2vo5Yr+GJgR13I4pcIHseCAhm8Nrw71Q/mRgdt0x3filsjIW
Ei/xEL6SfGKgQPuppE+rbijYlbD1+s+19Ifo8d1VRLMt8HhJzzmi5WW/gGhEhZV8JUhE+bJE7u75
FXAeMB33eEOct74cL3MuAVvuqW72joYdxUf5HKEaP2CkTo0vzzjRYbnmIAS74koc5EP7pL2UXWze
ZD/VEVnphaqbVNdHZy7XtOiG/HwR9nLkLa0XPRXlci09X7+3vypFwzUSKXIO0oa2Otld63Lt79/k
P5SL1jyWj/aJwuuHIz+OnKDqcCx4RMynWpzWaqyMrhgKXpX94qbHkRl8Etu+DiTUAd6QIV9QUUMg
liLtvfZi9u/GqDaglheZgn3C5TIEWtCG0CRPR9ZCx+9hUozmkGS0b03nSaL79w4JSMxudam9mRI+
AFfYfyuIBSvpbB/6S0pElv2URaT14WNblupduO1vwwAd+cOF5doCuMwRH4zS/UGiihNrMpMwkQNZ
ni8FagC1aOaBOCVEIonsyw5z6torW7O/YoPSkOyfrbV6lPYKUXENRJ99Nz3GNYfrI+/TOPNrmxAu
ftSwPUlC0S8oufULzkC+CAsqlg8pxGXP5TKMLmdkAhnnzWR/2/O6iM4IlCvhmA66J18y/Xmvmcxh
fw3ohe9YDNmbVEiFRHjjy1Rb0gBfuDaObZj+ZVmoJFSPv2lwAMEzGj5GnlVPYRO+V7kDb0EUcG/5
gY/ALjVEmBF5pRrWSl9GnXOMocLtwM6niZ1oWZa1rNlozQPlFyBS5JcPBKuTbhucfdRDWa8U81E9
CKv4qw3xzf6bS4dzoPDMk2HtU4R7fJhe8C/c3w7cu3pBxR/CbYPaC9ZV5MHqjW2OYcLTES4CgHT1
2T1vh+JXG52BZJqrc7QFzKyCnaudg9d50S08G+uTmYt/mUg+mcAd/xM3DXgbmCJsESz6ZSeob69K
shFvQlB2ho/1yyouMKc4yZlKf5ctwHX1tVSjeJ7Lcb0F5EallKHD/Db1oipAVwS8l6X3O4S69kQO
Dgg5iFwZKItFccVJaFj+Lb3yvgZBHUVryDbmMCIVF4VcChUALYPJfLgA4vXs6AiE+EAlnPZypDia
zsEgS+w94kKAZmqylQNq0zXLsINiSL405QzSzmHbPVuyOSK4VOCcY9Cjlt70vOCctfCOwSxzs5LU
YdUuQfWKTLsiAMSISdzCOwYHCLIwR18LuhT4ZKr1tJ03l3gQ/c0k52jhxJAzkrntztpszmG9oxtr
Tn4/pN3/muxvBADP5R8xg8O4bHMRqFpI5g9i9dq5OTesZ8sAZUFoOgTGKdwfAnsoEbVTORbLbEPY
gEmKnvVPKTwllTjZry1nSRpZ1m9SIxQ3KsL/HZdUD84J1BEPFQFKWxAxgXPVLEuIZ03LAE+JsFtn
GzcBUGIuHsoBN8/XdPXwHpUZ8G1P+s3BzW+XgWOCKGYYEuNTafQCNyz3/02C4wRR3aBTuGkEgz1Q
n9kSZagqA8a1gcvNo15FrAKyB9ZcRCRXulCq5q3sRgrwyGgfo5R8AN8KaemBNVOY8mTV+FML71eB
Iw+vT681Kc31Bd6HWhw6jcEbm9CQLF9Anjq33c4HVy9RDQDTWGtDGCa+ViJZY7ALxpvp5vxfNhIW
+E0LezauOS1vKOS0MQcKcZaoDUHQtncb2InohUWfa1H5HV26+tN4Bj7InXoBy7NMin4tMwpN9OEA
0/KFXz872FLO5RaVpkNGbbwiuAHC02DTERXuRBERVf2hO8CjQ+vIwehc8QhH/wqXipubzsVMbVdU
h3jTdGkMCjVRC7GXUjaZKtJ6YqBIy30tj0cG7xewo8XmSxOZdlBQnMssuAhXwrw6vd+Ab+LqNYby
AItBnD9tvroHdAErMJI3f+sctKjPbOXRC0v6mq3wHYoqCbs9OCvPYvXCKllok5T3uy+euTdOAmFi
0Q5hbx1lzmJ4/sKkqdiTSMXce7It27ma5eG4H6CElpU7yzhYIHBOAMejRSQeSHSM6g565ZAWm72g
bOrfNl9rb+1cB6okNUNmkSr3Yz777MbV+1mcqdmVJbAAUtNJcADmxZypd31VikdywWdTGZdwfG5e
Pf9GZJGW+Pn5vbXWgXv5NWaalpPdfNLTLkPH3SNjHglWGSU07XM2pWdn1dZC0u+uTk1PCkWgr5yY
g1hSScA04dKq/XYAwBFIGy9p5GXiofuh3qeTeKf1atmU60VUOr/Nb+wiSsAor6YQltLxNYGNkG5j
y3QZJ6giaMwEtXjhDRm75vT6t51lEQunquqkW9bGV+QmLTPa+AzRHS2dL5qJMlkqG9g3Gk0xePMA
zrlgmaMv0CbU1Zf0pX2jIoHmUpOapUMYn1IrswNauTZ2h/vG8CW8yrNaxURZwr33O39oEbkC6wWg
OM+RI6t/f04JfRY4ewACn/wYbXK/Cc9EDinwiWQhhfUSb+j6xaMVSvKAv2GLOkJ0ENZVu8Hq8otf
uPTuf8bsbcbW/Ot4uZKhBAbmoGS+ZLJZVG8VLUMeZ/DUnwrM8nl7kdHzUKvEywnJMtaYeg0/Zosb
hLPv+eAqFGZ4TUkGfIvBQaTa0OlUb7j00Jfiy9Jy9VSyjOdiv3hmXmkfe6BT3vIOUcJKOnktrJ5I
lR9TlF3cKwC6fG3DfoaginbwSu9ixmSPjkKxqGzLpfQTMPEvGA34bXiZUCmaPBkz7LQPiKoWGxbd
us+wyP1QMqb8yKDxqfonywzzC1sMqFIPDqCZjX+/5WxPMZgMsTtF07g7aLPv5r5gv3Rb5FB4pZSP
yqQkrrCSSrF+nWzgTmwJlVFY4MFZsVD6C/YcPHBXxbUP9ZxBKmlyRLSyyapLTwmFF5EjO0n9vp2R
6GM2BGhM2ieBVQTtb98wGPVKZ42lLHEJ9NsSVpA1K1l1XiVhTDMpcjIyEK4Nez+/FoXCtUnAx0dC
MXSpJ5wx2sktzos0+q34eOthTmVM+0F5/S54N/vquQ4WlJSe9RJpRVVU+m2WdxxLAc/3I1Xn/H+A
Kvj/gplWmhmdGFfPSNXXLseErIoN2Iyg37i8LDsGFNRtuTJpYvLpRt2Id6eHj74p5LIumU99h1QX
ywhWks8dkKZHhTWUf6n+AE5xGhgK6gzrSm2KUUjAVWrI4mrKBkYkPqhacreN2js5IBlHT9ls2+tv
fLUw9WlRMOt4yiRtgU/qq2jKBW7UerEEED+w9pQtegxFnDAIwX4//A5JkfaaB3Wrtb+eBTCKphXl
NqQ0bQg54j1Qh+C4gp41iW+kBynNEcg2HAqO63SM4kY6cF0JxwnBBglibT7Ya4g8A1YEbxxSoMOZ
udTDy2HeDZ7tB2DUIODYqU+HFoohR2yvFVyoNpZ0zzb0eqflDwb4WZPxo/FjQBzMAZ+oUWAlfZar
e+zWVyCz3hT0dieAqz1o8RpsiyUet90iH2OiSZp8sU8tBzkTMEUfWpmeyZiUBbXLM6fPiWVAhT0H
rDUu8oTKr4pnIawvOhd8PZ3Mg5VeaSmhUri9SoGwdLvC1jq+oj99eU6NRfT3CKK+HwWoAdPPvNfB
I5/8FB1Y7PZW0gYjaSG0orb5AfKFPLBsNQl2J3vfWeWwGeldXAZGCfSWPO84bzMKpTnSI65BJXAN
+sZ8cqZsF09u36jy21f3p74tbFVHcnu9RwqMbGa2PxX9GvuKbEml40P6K9KgNSKCi2MVDa0myFj+
shQRmrRHbTC1tAawpu+MLd6UTglHkVjf4Y5hNuc3fCSkQrh9uiiP/0tBa++DsHKjntwiawZp4CCB
i9K1+9nyUoIYcxjFuh8WGXMSKesG5JQVKXaFhOMHalmhl74kTAWKFfHdZzCBgq/O75ltJr67CYnI
OmMkXUp6wvx+Cp9Afl7kNMzxDTBMilmesqtCECc3fETHgqyrflVtvYsSZi03h6kKl8A6AD2kXqiu
5wWp9zhaumkjgN8oEJd7LiSpZVnrHvpuql4QEKwPuHpt/UJ+N71lOM7Q3Ot+DZ/oA7sP2T07LtZO
+tS4xONXo+E/42Mx6M6j1LxaoUKOfBvn8B2uS4X063r/QzthWgX8ukv6gl6oJavQX1NiPheVetAQ
uosTxshGof0lw97UX5UkSvtOTbVDOCNpzz/fmbYEvaX6SBfQDNVisrnQM5YvXXXJsbfMEY5LRd0t
4HOude2Iw9mCphdzEG0mfNWSc7gvceDMH0SYmTkLDRBprfKRqqkhQ/4O5NQjAwSAzCCBZmZYZOQl
pxAnc41K6J4HIEa/7HQZIM84L5qpkkhGqYY+zXYCQrvmsVqRaNWLA+AHav+KowiUdANLELD0nC1n
UxNOMFdS10AK7wNdtMxUYREURJ37WgpZJtCWtyxf4xvA+HHTT/CyII9/o8BlC9XiOpYvQWYazIht
eR70qnCLkGZpa0v0NqoDPkkyypSENDTd5Ed2lyg+q7AA1zE8PB7HWIhNw5In50jr5UYuEICVkC9g
tk9x4PURlbM9McTRfSZ1z2fO7knDlEZ4fkVbSwMimnNQ8BB8SkKu6Vn1n+cormq4EZdRddd6hnIz
qBPsFi1b8lJvLIXEvi5/4VbcGRhUSNMZPNH3/WaiSvNnd2kaNUscJ6eCQXF0WRagcJtqvH5Zq/x1
WCC2G/DdNvkhqWvAEwoDBgW01U8NW9rlCe/xWHvcLd27qPxGo8RnPMIAKZDWU9F8zV/oOVXad9vp
gOmN03EP4afTN1i3cCKWXad/QyiZvnwrcePdMYL0mvVej0+pGwr9s2MlOHbk0RrPiLr3KA4V9puP
ZWln9HtQYCYQ95p3vU+2Jy7/YpFLpd9zPYq3s6bO8zPTOPsLpAS22BAALH7Yi2RO2r3ytl3PA4nQ
zcv0yDuDh3238l430RxzNw24+R9w3vQGQZMKk051AIGVDpv0SuJmCgjU4j9Mq4JvkdSunUmGwEk0
uc/z608xNyI9HtQByE1ctUrVeVM/Z2XD1rRgYKjtRqPcmTkS4djy+h3IJOcklBYqPnZ4qSz9y2sj
USj7FQ7McBFSehYoRdavnHoVoSP3I19GcaZOqrTwKOpYWptwM27bhWVEb5rv85Y5Wg+NSYVrOs5b
ODxFt2s0rIXpHpr3o+UuRx18J34wdQlUEOjuXE/RBe+6wnxbTibhDa67nCFvX8wuJjUYIA6Zeh6w
MQLqAGfr0gpbvyZKnqTMIzaXEqXwrucepSdscJ1ajZoThhNz56pKb0TaIN+gWHiV9NOuDg3mTMBy
87pin9w9BWtJ4ZmiCl1Pbs7XC+UTwKzS+PO6Ykh92W6cn+BA5dU51bBsYuU0+476sXjujR20i2EU
f94NE5xsWjKMu2INn0r8dsGKa0F1zIV+fcLLdtRdo+u3MzPPDVB150pKRoK5IP2in+REYiVZMqid
y6I3X9YJCVkqGFvKnVOLFqqzgtKXcCwgg5uWCFB9s//9W5EZwLCDxXSowqrliO508+SJCeJdDYko
KqKVt1NhGDsc6AyuEYbHZJOavrF+EEwtB9x0Fa4WyXSQlTc0Pljuoj+8dOvdyvmJK0hLJwo2Ai0V
E4jaD1NdTvRsjo95zuv4Pqs6rHrTFlr7v0GkBmNeyPLc99MobKGWyAajquULM6nwGw0aNOZiyScl
NVHgtzDk2tVDufuPaQHTO73tKjRgJUocFWY1cmkc4SSAAZg9kfinmP39LXIrjsFIuQIE3EfNV76J
YRK/z1nmrTJsV+4sx1C8M8ZZm70G8qzzZGJDGgB+8k09gUrHydmh15ZtsJc56Qi8wW+npJDKBR7S
gYl7qMebP06vPbZ05LrZU4jItVOhfhvD1arsv2pzmb6PhvgoT5UOjpvg/fw2buKXK7IHQCiOzS0u
p3Ei45W86wX9oZjwxHhV9VufNsWJVYig5ffqhxwvz+BLwtqfENL200xnKD18XVDRZNhAH275Qjeb
eHt7+OEb6ZkghVNyzZI/dzG7cROkTDcKA24efELq+W0Xrxcbx/bOx15IXA+fWXGM86qItMewaL1Y
FKUzAbOWN/ncQDubklJGqu0RyY+HFfmV7i7ed4bMEApg15U75hkxSkgBAvp7UbpvTcLVtnaA0Vu1
1AdcwBeUCL7SqsyGrdMwG6kZCY/4Sj/WV2UBVuFrPYJKMpBDyGbKjApyiQCLCwgk+PYlpqV94R4Q
4jO2maOIIPPPNZBiayQJPDbIDHhFvoE4yOrMQtC3ncQ/Fy3SiW6c+huh8CPtGf1nZOjAya/Ye3XH
zqOFod5+drCLd18v6Jk3/79GtgR2IPDSqLl3lgelqPFn+LQAegXjQvncCYUAhyhrz23/pakMWybA
0Y8JdWpvwD6xoFvWamQkp837ahNd0hNbjYHiEpxE0gUQL+AAABmxD+dHrnqDjz3D3NDiaJ9bDI3q
AoGZNtIqDdCblXr63dtNuwfecw/TqrU6HoSlUXrTgfbKLYEP/yr/SLkLeue9B14IWqsT5lsL/b2L
zk3yRzlK4B07JCsVEZTW7c+bmxlzlZNtsiEW/Isqz+Q7GxykDFyu3jeYSG+gVZh+dX+QQbk7jsy5
5IUpbo+fju9BZBzbL6SbB2lrYI6hlmL0dZip9hMQe3fIzx8P8upHSCPZkOgFHvrDYcuKjbcps8Bv
u0Ca2q9JQxu71WNm2wbG3T6KHmNZjir8sDkvecYG9bMgBO34U8vuRh1vlddo6ijEvu5eET4dvWe+
xtaHuMnIZOlk6jEsiD0aW3/7Dp5OCMTMGzqayy7h0OUuvkDOfGymtCiNXwTJf2MZFrnjSkZLyO/d
Y4Mq1eNfDNoVqsYyBzn3nR3vpX9LfIWy5Lxq1qTM4offwN9xpA3ViasdTHC+8wlVFtjO/HYDLCxH
PUllEzBjB4HOdAqcLlC96lTzZ9l67Z6CB2NDWUgMxtUMNs7r3M1/XQU7w6PEJ/LIhO/V5gatCk13
qZduarsvqamwlf0sp5rLQYTI62K1eBFWB/vueb/qOxql5o1TVajauZ+hASkJ+iXMr+ztHvTNL9IY
YXAK+stjBtvvHGvNqnO3biz9L5sjIzcJ1LW86oJUddXCnKrH7gYxep8vU6UJccG0VMFCtSlctpgd
4R6l6yy+3G7bHfeou9iULqhoegWRrjJYbI+Wh1hjtPHzP9qaSD40VZPGU8QcL9g78S2RoaE/ikDd
5/dhnOVd5zVjVOl96mprZmBfD7n+/mGekSRxcFwDJJsblV4ibVboYuloJPdJiqD5AhjAYkaOUQmk
iRWZeVQLUVhqsVKjbr74gQqsYZ0vuVAaWiNDM7wMlgSBaPFJ3CopweFt9DIVyLJSAxLznhaE0Ps4
DIIZxdq5hCQAWCg0fC1IgMR0QTM7C/hCLk4wqkf9zxuI4uHBnwJHnDYZGbio7hjP50BpnmZZX0Nw
MIASzLNVIBQ7LQotmsFlaRexVgvVX9hlL55V4DxiSzj2EsxpPA2wydEVRhHkmGMoTN5F6+YQMxMM
1eS+GbqUkNJx0jSAheSYJbcFqpr/rkPGB4U2+ZC3h/saAo3ioNua7Cda8Lzs72GJhwKDYpSwB+XX
qf74MYVDSboM6qZUdSYwNqOk/aCzGQnu8ioXL0PE3G4lxznwZarGoRjcOgDK7jfvNw9IP/Lfredr
YOkrwQYzSv/YWdkYAnncFSDmt1LLpB0L9twL85fzM/luhuMh7m+C61ROVISy2yBfPD0EyrkoGfx2
Qah8gB5XJbEevdDycEZbgpxlFsC8qx+0nxpYIYFUAKxsmFdFRK7Z2/L9gWR0f4DL/G/K6K7Xmlo9
PmfLdMBJ/Z9/Njh6QcxAY7Scz3YQzcODhtZonPwuJY5qkoiLbC6ONgp6qGMlnTV9sj0HxHjGLXS1
IfYlwiB/Er+o1ew6VpIsRnGHttu3pjmCmxDdkAfFh7AuHicS5sFdXlUHc5qZYCvAXzFLMMxCVr/n
TsAFGruvXXisNhBHxjuAGqW9NyGWlYTwSmcjGkfhwKHFegoeArrz6vTEd69gkpN2nXC9YWopQfRn
05ENmNPTvOEjkzBWTdYv4kth1iSE5k7XsJQZCgh1qvJvgSkXZ6RsmIl8uTecPlYJvq+4bQeMPidv
xOX7DNcHNsApGu1H0vEmTDZHTMmWBC9RD+E0iyP5eKAAmzVMwuR2QHMyjg2PVm7nV6IavRctgVFO
OWt5qzBaleASDHZu1CXNlBa9ZDic0NdZchQbCRXDH0p7SodzltRyVuYxC0ccc4cc7CyLPjtwsQhn
q/mdF4M0HF5H/oNRWMlkRoUcAa8Fplcs4WjgTAOslKNdZFoXn2lE2EiZXv65Ib41q0fkjvF96VlD
h70TWQp054bDBxpV4Mso3zBFf7ISqc4mXyqqxl0ZGfWvsWHN4j77znJ87WhLs2zH3MuoRM0i6Oae
W1lvbSggoo/Qq9wz9xruFZzHbUyKvbQkm/Tim9w5/RTOvk9Je8+QWoUNEyQiFSHt55AH0DbLguXK
kx4rLDLqJ5tsx60xAUr83jXeM4LJQkaH3gyNUKTrIPlp8Xzxlbve6OXrImCQkD2W1dAxyG2IwOAS
O+/bUCiXWCT19DVNkLqYiNYkAewnsAAIU9/yLj/1YJVIlcnM0J2RCkA8mDKPVp++IsTvuIlhB4zd
tZNDwBC10ExZffqt2wjuAfShAES5Y2/Y329Qf2J+d9RX3oS+ZTxJL3n+cgOzoajNXul/HPh3g7Qa
HvP019PhtZBWWITclk0Ab49nBq09VByUihDnu5FuPsTZmE7OqnQLNSdLhQjwBvtFGG0Hg441wVJG
AK7NX1f5PZCFTaieLeCsDCcvIPAKAiNP96CltkhPlxxlgftOnGLtcVCgJZGH6xjIkzdmGJMPVmYG
Z8WJ6HK3WizmQG50EO1KYKuKNxZxi0dHI4onH1YWFewwCUf16OOVXN/I+twdtw2MxeXZ9ryXwwcj
tez9vf0xh1V6bE/6Hb4236F1GOheDKr6LHFENKwB/F8uh/BI2iKnHad8jSsuuLkR2/LanpmXTwJF
EK6eNjuSJWA/8phaINLSlNDWbNqvQrGxnfxrH2CCp7iIeZKkoZPHvLi7RCJfPqzmXpkhh4i1rxEW
IH5EYmvGr+JdkkgHXo45NcyZVWqBmqavKoGBOgti+7JeGfxEDG846dxbdFfU+hEBF12JnDWWSpZr
SkFlwwBVQnDfMHwpR1oTjXPW7L3/1ZKwhamQctqK4QAI16lN8svR3Y64tJV1mXunuML3ZjqsYpV1
tVSzpttqkP5UsjcWXImNd0pFwoGc20TTXxLZucva8r2E6BXBzy57Ogek20DuvOssT61lrk5id485
SOTkUUxGgFdXSt8OLKBl3Rg6ACEwyDr+lLJBYYNgs6L9UUH+dzPA7tlwgRU+h+dPQNw4z7/ZTHzA
lU9zxXN7xjU3b4M+/c5Lj/ygvOMBK84DJXOmgfNVUeN39g9cMmhHjQQD4vrrWWIO844OYrPmjKjS
hMAJ5ORVBdBdSCIuXcm4HTx7vmGzwX2YO0Vtma7pV+gLRMLiUiaQQizAtKJpCKbukOm/YJ05wvWs
zRBVWs3fX/lIs1NoFiAOjHVEzUMXDpNjSY7adL/RpvytnejZgdmGgVjs+q49C0uEHVQsQYuNHD2w
LyUV8Fmjda30eqXvnrXjcQUlCS00UnktBhUA6JAdYQe6BwDWlmIYYQFlcFdseTx8GvvLXKtGv5CB
DsSbPU+iroOpBn8YAvLaJnk+ub+B2499gEFg2Pz0C59ajJ+vSTywArMVoUPJtl/P9DeCSsLSF34S
R/aAdbh8tNSRqveYR3OCi9TPIjCatWqgyVaJRNKo9fHa/2ymCppRrw2yWLNYAWSlNpFC7qmWA32B
kKmrQ/7QxJAGB4ANkkLvLiwhVWD8bqDNBIs4UquGMk1juXytlA8si2XGyTgIljQoThmNlGkJLfPn
PTPuppPTZgHqfMnx/gu/GXc7hVvZE9W7TWnYFy0L9xfYiIvGiVkYsdl6eO4xPKezsYKsTLe9c/Ha
eheowF+XUKWqtqTNWITi7wzdluewgskoCiqSqMZvTZOpOXGfZ4MIfZyZIyhHMWhyJMBKd5CuU7lY
wI3A5qsAvD/XQlNSbgR6eTIslFA4pnELxM4WbfKpJpHLNWX9w/Y9AyqpU3sEDOLO9nvRAXKF8W/c
bMkLu2SVARFG2MVcaQ0LEwQ5EAFvgv7T/eF3P1mFtkekeaFV1wIjJcRsBKVg2XmNI6GH4xmnQRyy
MzPV9hODYqZ6J6ycE8/PC3NoL1k26J7S0zeDswP1NcYwqeavU6QpBS9XpXvDl7qsytAAXJwSiD1z
tTJUHWfU5eNEW8pgV7n6JMb8f9WFcfTJy8B+UEhqbsysP/xB6csxAWNBT0C7SWcRP62HeaGnr226
D/cnUoOiiomsAC9sxFO01wPln+iF3jX0GkNstBdSsTW+8HgZKLaqovkMMxPQhkHP84ymZLmbz6HG
qsiDzcH6bTj/utLAyngYAF4JJCobycMJbugs9rJ3mXL1DbWwXVjB+XotVd4S2aYYwHRbBJ27wmqH
SmzdVO2JGC9es9DAYgbghtS6HSZck/A34lSdwydj3nuuFLW0jbHdO7Pz8vXj+JAtXpFzV0txroMj
hYhleKWjY6Jae31gg55Bi2qIVkffk1zOgMx31iOP9GPK+mA+v3Bdb/ajWh9FD/YW7USDihXoin7G
Y5fLyDBD/Qtys11MHe5GLEbthw1Bz1pZxwF3mHAO3gcle9g3hDjAGYZwjx300ae3PcMznxBPZPHu
YR8wKHfOPkz8ODUrRXUoqmAxqnbpu2hqeZrEhZCbGrFzHcNx3qPVF9IDNvQ0MQ0onNXDNtOCSFkM
NBRyJV8z7K6LeTjCW3pQSXQn0+RbjGdTkigvohgg0Xgr+q0LPvEztJS1bp8kROOjsNhqRQwpfUaJ
VTe2v8lGOMUeCMQmCFXIaYZjqVASiYhMOdeGv1V7e+cUagiPt1jasfd0XAsxv2dMsuGaM2ouneN/
Xj0YWWuW+Li7CqVdLPhdzCmL+3YPFs8DnpsLOrT1AGjxToyyvEdO1PLFZLjsofWIMUm4WN+Y/1J8
w7ApsKQZiqV/Hk/bmnYRxmzpMIX1cdxdWizO3xOxiywnKfTtvOxMAju7+/wtUpHCQu0c5K3awUuK
9dOC57sXLPn81wzQN59eRqbGAadKkj06MzoQiSnSjS8nzgKmwuM7IY4NZbJKm6o0rII2qn2Hy1Us
R9iFhc2LbOVvX8pkEvysUq25SeNqngcgsyCrifupOe8jAppWXW6bE8/v1QVkTDTnPOXvSp6YwY7j
rtrkRxwRbNQxWmaKqeVxaDc+9cKm2Khl/hYXLD0miZS+seVhxoMoV2blDkY5CV6nPgC5fTneXXPm
nnRgX5lfpAu5SJEVzi4SqyHH/EQLRgcAKJUJF6ChNk+dqhNd0YdgVBLX29yik+JcOzfj4JY0IuCf
vTytzROjaZvE79VUK5smIr356ShGpXUfdShr76+KRhjSAzPut61Bmcfns2HnwW6HPPxawZNA2gH2
A17dbTgAXtML9+5doIGhwRrRPA7cEfDmSYwHBn5D7vmpO3OHb7YKSnjrkKL7FN+k5FQp4u8xtVze
+QFYgURrkm+azDV58aqHA2GZtLcaY96nctFt1T2QSjy4nC9ym3YShM/1N7oXYGKuWUmzdebg/Jhx
5eEOHaQeMnELkh0Bm3BJvbHpUErG5bS8qCIIBaQrPSoVHLiqPi9I4eobgrNhELq9/cCZmH5OApWv
M59CjTjOyC6hsOjkGs7d8ZKlzjOPd1CQjtmVmrFbRV+xVlm6enEGDlLCphIUiLmVgYE2gxtJnmb/
qsEBT8v08NNgXe19ewfmU03weSpqW7WxmJTemuvQAsew/f9uyzZdLfcBNjCRYZ15LLoZRXbJtNZz
+hcNHHcWk1NrLcRcnPWcPoJJ5MmfB7Y+N9LY/sLiV6IkEzFpvvvs9dDXnmWdUAAd6UXhDrv82p+O
hdQHcpRz3pCEh3DCzvfACUqWoRltCmJEALcny+2RHymFUlV3wuj/B8yWX0KyS6l9J+joY6oDyTW5
ZMXd8+2lyv56fpfm+TSHjfFoRVDCnQIjCloE01ku6htX392GrKEM/lAjf3/N60qgCOgniiewObwc
vf6+I8UEepM5moNYyExcjd0ENggeDx31J4rHLh83VEKt64DVoy2nDUMc7rzSC1ZrAtu2UrCGr/WU
NH+p+MjDuD451hjbRvvfK4EZmnCUU5p3CDD15apsLDSbAwKHqJA4Uno8rwanfKDgk6MgfFtfHjCc
kJRoidv9Tl2TqLik0aHMQZ+5h+dwwhjupduHGjNQdqMQQDs15+Le68qsRl7PGimOV/OLPirPg2SY
MDiA4PF1BL0hKWkNmceNsCe6buMx2rJCGviBpawHMDQfoNnPCPuL+hY9n73jjX2t3INXd3hbWQxw
1HeHunGSlLMKUaQsGwfyN42IMB4HYKOYo2x+vHC5dG+g1cK92Qdrnir8xukidBaHrebS5CStfDWo
RasdTiqSYUKxtwtLBpiPweOAEaIu/zd31uomedezuRgocFwtclx3lKgfQPXAVkdmnayBEVnoUgEY
FkFnp2Iqp94KRDbhg9ccN4Ayo/Q7YQSA5fqH7QhVlEY/WMEFW/8mCPpZpDMvctfgWdiAOblW6Q4L
+9qbX3dv3Q6Ov4NfrZWWgylee1fr5X91iKOSenMG0fFslOX72rbucSEOYeKfjCBbI5muhw5bpW/i
3idHv/l/fyQsTq9jPS8IfAFc/qa5tWJvqsXid3YkvdoFOtH4sArlmTt6pfmn7+t1FJdq1SqQbkPt
etpufvkl5dIzthq4AVeBJ2cZnkCaLoJ8UdCjY6U3Rwm2an6C98yJAE/RHEkU6dWjH8oi7iN2an+j
BrtxLd3ZOjX3e1yRqFvHr2/hThQaG/3jvJ4gnpT6dVqR9IW377GzMZn5mGYv2O27DDDXLaVmqu84
5h+iFjQoDwnPJbDGgqyGGhIFQ0OMRLD4Aztutin8U883tXK+kwCfve+/1OUXOfXll8ElJFssNg55
KzOfW5m9bT6jnBQwxRP5dYd2IplQ5P/HT62nr25iJ2e14fIzw/yYgqIDZ2tunDYm0fLP2TsJCn1M
ZNsSdO8vXTL/WukGOQIX2bpLGpBhz8ED5+NECbSoYmhJkTTx/834poZjdOCiQUZdLeE0FsXgkxFD
n2iyJwOa70l+VTTdy2cuneZkJoM8MeAX27dt+AEeZtP0ihPI7hcoUDcO7z2amCR0k+B4XO6a/vSl
DtZH8lCYxqNbCgQ6A+J8sZAolMMCAnekP/MQn+OmYMx+09sCe9sA9GaCVbn7p2LHTiQi38Ori+8U
QEJcCsxxKoRKTIYgDDiPakmxy4KOKr3544xHk2WZjqqu2VnoLFU1P5tiUP1MqDC6raYrFAl6mAEo
R4pEdmczbbd3pCmUbmQuOraFU9x+BSxpHdyzUe1+dutHD0r7rBIJeadW3g7Ymig4jDkjCxjpqdd6
DK72T0XlxUyiEY540hAVTdDRPJ1sZD8S4HIV7Oqi58vkIV/auk2RBXJrzpr9kf0C3Qi+7aaszJvz
eMLM9cUCYDa8a3k6/Zu77GLmsi43voHbjyTrz4m2FEg3FkI507Pwx8Ox7yEkaMGZI7KZPA4Fh079
LMWuqlxrylop7WEY8sT5oiCpe8MSai2HHWahP+kwiJhMUDuyfKyEZMJsc/3/dZySjw/Q+zQx+pl0
2+wepNFlhpq3+kw2seLxRf/nFDLtQ+8aqW0Y+3lF/Xm1icwPTyO1I75wCvxRWtaNseyDhEPghvMM
BlrE00+8L9PQ/58FyYezZ14krVWrY2TokdV/1sSc7HwNzjRszx4j49ibZVX70pNcXS7El6s/EfeE
847MA6qog5KFxRbfy9H3EA0kxOMWRqGA5koAsYVfAOkLjEVp4U47+TxrcIHWDsqcWFqnmKz4UYKe
P3glG6YC0wKPq7A4lN7+F1YGHvW6Ry+1gBy1z037lFIXV9N33bLPN1siOEQJkZUyIaR5U2GXKkdg
Gg4iCFFOwagVI4M019HxYghu0zSCjyh4uK/1QG0MnsbE/BklVdBPqGpanJzmaS3W4/8NNdOKPY7B
20HB3czSfJELfAPCDgj0GlAHJjapN4dfCMlIzcYwNC1ogACC7Zs/iLqz5fAvZLFri9tG5I2TAnZf
RhVatnkIxrgedjq3ch/xoXfEV0dOh7mfYMslY0NDzz44Lgnp7fji3nDutsW3BhetTDdO22W0g0eX
oSW65GzWm+B6NoXzTRI4jSmAXvxDEh3tWsC2xU320wmufLyB6d0PxvQp5LJcYA+VXSiEZWWQmaxm
OnoB7I7RY1TcHRGIu2r0N+OvgGddi920p5jRGxMt28piwowkP1sbfGnID8tD7yzGvfC65AVOMJZj
iigbD+g4D7vMdvklWj4EvyrBOSIvP6zsrmobupUZu7kdWbY7ewWdL3CVuane3sPbtbyy7KiE1E5p
3ZXqkKq/5fPMjI4Zn7x5QPbw3Cs0wUZPwpkZM8qg1Tyu/v2yQ+8ouMQt3GZd8UM7wXMdjow5LdZX
Yzbw9zCeZoHp/kdsIWkF68XpjmuwmmpFywrJN0zR0qVr7ymik4U1hMoeRkPfTh/H3RwESEdScy7E
xxH815eJ4vBXIgnNu8PFQ0QLiVGoUrSAfyozDHVCGsm1YyUFpj3hT/wnbJdNAxLmvjRKHtwKYOVu
gJMm7Om4QowTdnwe3jfHPFHsL7tXlMj5gfSCyuewcLW2LzMKi0VY8dQy83/EYJ2m563/CimpQXza
wmtaKhUVfXe3Go6HQ5t/dbkjcJ4J5lucx7MP/VRkOHoDpksHxr756sa5OzgXxC17skA2RMZSfb+5
Mvfrr0I7xmnST2n563KuTDCd4YTZ0rCpahh5I/Uyc0Dj8Wxg2ktCchpLpFUGht9i+fKh5JgPB3ec
inHzq4Gun09bDJAPg7zINbjN3jqeYuYtDtnD+W81FfGj8Qliz+uTUQjqlIThldGV1+OJOco6WeUr
nPTSzZ2j/lZp9h23fw5uRxqG1xfnRuRChcw+lUjMpKBQvBYlvR2pELUfi7Jd3LpoJXIKx5RyBOpc
MxxHYz2kJHhvA1vE6seydpDPMR6cHP3SJOM/Ep/OZrtHIyLtS56uVX8tYp/E1yDwbmkOD3z5+70a
AK7hYWZRzOT6k/u6zHhTWqJ8+FCd7XePYZU1dh1NuIPA/IEqPapBkDKfYWlLY/eEJhFCgpS3WnIf
o/I8vNzsi5s84bDrJPI80WzEzFhZ/TGvgY7mIG0YVkyCChLqkfMyHei3ITwR738aj9zo72QurkAW
i7coz4Irm63zGinzlNiA4L0H0Ma10Db84CW4w8XPCvhRodvol97hVYZ6Es16y50M3B9eE2P7r0dY
2u6ESTQAXw8oj+NYavHljqwWdU3MRrn9K/eVC0Yy5pUQ8nW0Dmgyy7z4HMwPfTyluu0HJ2QosdbC
UgYYR0dpbZXSKHAUgqUCIVezaEkkoxpRuhKD2M80uWq9cXCGmolw60Fba+JrKGXJw17ZV2nhfLwZ
idiHjf4Sq2HgbColJWm/sNlv55I3Tdha7ZBlaLtGUpBAtvpfsDjEW+w6NNHaibKjgeSN5tTasVSr
KAUESQgwJsMSW1HRGZPuJU2BhcGDGSPpWkrpP7busV6qJ4zH6sS0DfbaTvAHcfIELAHhfp1mfxFT
eKse1vKOrEyoYs6u84ydWIyFWbm4y1ltF6O/x2ytNYOn5rcWMPhj5/ffS2nFOFnc4IP9x4ymUwa3
Q9Lea44DiTWlBuHk1PC5kJPLvY1ZzLhh2LBUy6LNkehaz0ltaGSp3wCbIpDr05U4P9jzDG4r5711
4qYbmVMYfVaU8k3eqjH51Xh/JPvsqFuLgAcG4EhR0N9FrUHqMt5rrduir0jmwp1NjcOqkSuKkDl2
cNgGH/hWkxB6F9xGMFn3SdBTavaozfw5/6+Nv5n+0j99fk0wdoII9CCpMMAIoOAtRpSbdyin1v1n
z4y1co5E/wHYkRpaQ4u4O1YegSF/hA5ZgNsd+kX/hfCdVKl26qaa0K/Ng1SrESyZOZcKnjxCEzcq
ThEGWuvv+l1vGjBx7biX9+Er2cgHZBQ8yMmp3D9LSW1HuI0PD19O5BIQzYR4shhngvODohG+jiDr
YM7oQxUZNsfkJJolR+9r8sGJnKHDmmKaM0Vi1rp+gdbU6o4HduUoiQDVloz7SQAhqihoXli8GQ+m
bn7i5UczgFXZ/K3rR2Psn6dAwL2Es8znwaPePZAH5nwQRnqAuRjhIACYcuA+7Dc1W0YNExgVOYaE
9bUNsL6OZ3Xf2S+CLCz4rF71HFOAztJaASTqtKv2NpidafPfcRAra8LXS8Ob+PVFeUVLB4gp/Lyf
irKidsK73RepjVWbZeoasAtoaZHktETv6jRgAEII1WoNxAjf9SF5VLY86n6yZCWivsaQhtvx06wD
pmd6fLPdExF4bMQ3uoxqr0X01YS1aTw5+BkQymd3QUv8MoTIqAEwhit5OBn4CuYIXD5nNAGIT9d9
Zy3aDOBfBOFiY6lJM2G+Ie45eGwLMSkZD5FAeny2Uon6yk2/UgdoEZHdDGbMaiynQZTRx/DX4Fpu
qsMtwTM04eSbT7gXyqLlCG/szkRLDIPirNthh+IMUiGZ5ZqKu9Oue3EXfkP7vU+zpfEZNwI495eX
gXLpAeVRHm9yr4XfEkdCmZ9DrbARw8MtpAGd4q3qj2qx2Ud8t8Gsny2p1jWJ2zQvlgyfVdjVaOWi
qUYDR0b13MAlvAqxGJ45NDEMUDwPXT0WY0KsR5aXm3N3JZkGtdPdHVDLf3CKcVnZ3/MwmUf8/hHw
2/Wi0ufCdJsQF4j1txRH5rcnbOzg6OcvuWCiXlUSdlsASDx770/yIM7ccl88VIoZv3a78MPErXLw
3qGuSKVEMWNWuEtx1ApsLFyWVmxG7I8i/HulICwLdJLVf3AzzsQ8XLutgvbSQaCBvaXm33lr25fI
IsqMAcIodFN1nt30tCmH/27d0irFaSpC69dDJumtBg4GFIoHwCRNd7VVMSY3dYpPGHi+AS6vqaag
5m/21yyrJY4/n9dcR9aqNQCaw5g53+8+oLGvxyX9G6fXlxvfakGxtrxN1pYP8KXFiqqNq0qezznR
GLFMxc5Zdstsi37HX4O0L4BXBvOd0PrsKy19N/1cshcjR2wnLccbwrnwWQmM8bJmcm3kTMs8tFgK
Oke6oFz8cwX1QXY7+KJ+yYghYrsd4+9KxTFHGOSzIE/qKQin++/crZgxxHFBCwbYo2XHfGCe26Ie
uXgLI9D78X9s6RT1U+GUS5gQ7YSxmEtkrlr8jixbbl5xrdNb0MPrUuyeTmO4TRfGfQ87kjUgxIcL
BVzmj9OQxJmxdbZlqdnXj3WfLt6uLvg5vnIu9N5PIjux+HLQIS840aWHxfRw73gs/6jKg7u+ygkh
bFZUz9o2qxl1sRbuDh4TkGfnan0P42exj+GU1nhN7R9XriyeDXP3quvmMC8gL90survX56aHLx1Q
latMmdtYGrVaQvt4RdCge1amoNEXb0B++RdcS/ddVHTEeUWhLRQTzMVwDclyEbNU8/kba3e2aRRI
SvUrnYOp5NZ7Ijx3nyw7oXuHfBxYqZgo0kmTfzQU48NWMWIT50JNxpk/yzbKy0jurWdI/mDxsbAn
/7hoyoXOv6Ac56dOEnTrGomBRE8DZ+SmiBWAWYtZVye7c1yrHUyISyKUXgnoGSmYMkKGVAa82N4J
VnYFgGBsu2OIqY4kDl2LnUs8QmG8rpZomXy4SNy1ZAaTYpf9ois+jdZvklbku5+Sx5sHtQdfMdPX
/rIrsC3JSvpw+8v8l41MjUHEIFa4P6zwRjLITTFulBPhzBY1j/rD96u2UDAO3FdGfdHob+TQu+cJ
l948GH/buGgyaOQZ0glxH1qh3ayNko+m9kg3F4go2sEusPweL2tjWE1rWZdlhu+ebaM+QOHuvK5x
xjKYb7jQKMzEtxD0VaTRzfMEFV7yvnANpN67R334+Wbq09o68KpxoYh9enIPvEJHEpYPl7ujpfPr
Y9jLfdrgcWNAqt/Vfbobvb/NYq+XeIoKUuyzWVqRAXrjYjKt/LGc0j5TUvv2CbH0bufaATjd3y1D
pof0wx1B47coQjXdsW24ACBOl6CCIafiUaMpvzJpClL9l+jCWlGauQZ6JnDFUPXsXSgMyTJWUWzI
2uE7Mm2XLHEHNkNBDTkIkEvKMQN/pxSlWczLiXbzO9L/GBQ2Scmy6MKoxM87qktgUQjCLL4vUxOh
KdnZ+PEQgVzQPq6eF3yBU826SeddBSEIQSzMgd0wGsGAtlEhC5+spGFqfLQsNUpdIPRjvAk9j7C+
mEW6TaHwdnJ4szbxYVvHedxg0kIiaPzbbVtmqeISpZGSrdKyDl00XGXvTHegPt40Q1RG/7v52OVQ
NssOPALNJH60KLGEl0M6RHZQ9oV0Q8kaOUIpfoTus3nJIfLvXVvNFC+7BXI3t0MEGbVhJgJFTfWf
ccR62UouG0JzHipH7FDYLN2KXOlRjgYPQf5UjW30Ri/zrEVu4qqXKa85dDTa7FaLYwgYBUIoaqJ7
W36CIoEQTeMorz+v1dgisct9hPww2ZHJfnlkIEjag849btnMGf009Vp1FnbohtG1FcdRqJpds8wq
+Qp2lTGAkVmu2r/Qq3HDg0fj+wI5vp2C7TTet618tqM+Pu1ExAESZPUTgoA7D/JA2fXg7Eu6B8U/
9RDfeQzwSQatHtbR1Hg9fPsu2D1zP0qWAqLZtPrWxUvRrupHVsFUVf6+5K2Hxf0Q5GAq6YOMYYHs
NpSaig7mfG9AWinn9hgWhHLH6S0zYyorjJvSzh1NN7LoN84YeWGLEJqmKKKH3cogX6kV1FS5dyT7
l5mMLRWvkKejJ1uo57gufB8J6wRvSfTqnTfRjxM/B3m9aIbw/pIBtRBcgv7jKqElqA1naXlGTSPi
oxw5wsi8EujZaC61FJ6UqNmm6JquTI/7LvPYgbSnYiJ48LykzV/qYAWnM20EwbKadvLDg88SdEc2
d8Z09W1DC5TSX2tcjO2+EAvyLjgS2dVvLgVgzuy2NMFks/24ioj045g6v0+az6r7tAbzNqFHIJUj
VlrsToG04l0ZLzU0+oSagRVP7hZleYWEE4THSi3XuKfKBxL9gH+bZVmBybBG6wsRSvQlNQH0HGEu
kS5Y+FbbjzphZrnw7QecE+jcHWUIlyyrii954Ri2YUI+fquaHfgdtaN8VCDYLf8t2T49JOpCKpjL
KIgAP5Wu6zIYQK45vhcb/8Jb0ZKiYmaGiB8xPdCCrC6zR+27fB3U/jGOzt04UxAVdynOf9+VrOtd
QeejIRkBeip6iBwh/I5t+aLDzjtszIgzFxtsS/r7L6WQfS7Y6WpAuWYgCEvAhaL3uH1tJhgseTCo
gdTj2SyQB1PA4CL8IJn2wU/Gt3hG1SM1hMA7pXU+h0i2McOnBppVRBxiMu4dyjeRzpauCCZk9Wbl
Px3vWJ2ASUPXIWdouzh1rlWfgmqo+g5j7InXDSZZToYP3QJbehd6FFEcZVvMJtI7NxJ7UxceGnQ6
OIUfI3uehk2CiKHcsOHHjbjDUhu942N3/cmv180vNULDBc2UO/k5w/PHeXsWQblV3HHev58XB07Z
yO3xvIGbUPQ8ZOgEPD32vWlVIfJHt1gqZj8rRsXNsJpiG2v1rNMXvg16lJx3HZUCg6dXTyn/RkTf
GG2+AkiLfOoEQfXFpHJCszpJdkNp7YesMOJclqlj3/EgBrEB98Vx+8cSgKf2kI/K31+W7kQBGEaN
87JpuUWRRpT1VyI95VfCjeOD7BP8/VI5ElCf2ImDRk1TL5D17YEJjc/ZtL92BEWWhDTHfOHQuXI+
OZB7CGDk82wyZFgeD9D8pK+8N9nFmouy1SPL9PEupf/5dt99SPbOKQUyKIOXmgvqig7tSbmSgNmI
wyN97Xt5IpbBOxHyYvn66K/LFJVvs/OIsjbd7+5xrQ0TAfFdHP/AFpgFK7HOMzLl8E6FTmUU40Ma
FycMX7lVZjSm0VH+vLn6Mhzn+KTFpmVJDEAVApGn2CDO+npAtwtyDSap2rnAZ0CPCrsNhB55seR1
atlBLTxBOz3PSbzfjG0WDuq9JI5R1BcNR65uy3Bb/II9RjWChelGn7wdR9Iz3ZVQcYvjAntOaTYJ
MQiKSTQuFEY/44Wa8yYIz7UC52e9xFda30VcJdBhEEupoEf5lc1fHJe7VRxg1Hsui7PVWH/Pz5DO
u6xKqydx2QAtjNZIZ+y7MTC6naKsGgt/m0ohZ2Ol2jWRXZz+U8g1RhEv49Ce65ZU7imlhRQgr9Ra
D+oH66oimHj+k9yRNd3/Agz1aAvlczcWBqAX50MyI/vFsUilT1daVModNr9zKoTvfJ7pZwK2z3Db
NYTHxOw8GEeE3Vx3NmWnQXAq6vbRkGt6+Gs6bGkxAN5SvdpBA5AKU06sDZm/inySjt8tLJnqz530
kHkXpAMI/1KbI2eewyqLmjrvQMCRf6Oe/JzLNHprXE/rBfi+COpH3HunEkJDfiQKzVN7nqbomM7Y
W1CayvdsOwMstIeEHivmdT/eK2DKzpKUh/o/8MZ7WXj9l8iPGjV+OAMmDUtLU5h9WrUhoTfLT+4/
6sFMs4jNOGmpP9GcfAu+H71ArbvPqs2k0S78EBUtNSwUNJsLlu2OHc4M5xgpaQjS1bL5tY8LsiRt
XM2J8lknrc2njhnSHravKDU1PlIp3kDFr6VUbg8SUrwxwlRF8mBq5dk3XWy5+cyI/uS2hR7DrgL1
RPMIuvBCr3QDfEngPa6JMgnq5sNeLq7Cv5ZbQBK5Im2KCYIf8FbYVoM6583TzYdNidRipf0wjYFt
9kxL5vX4F3BY0TYoDKlXKFEj+IfESFEHhgHQB+1DwdE5Jx6T6G8uhgBlf8Cy7lgg1SGadN3XVfmc
h1wwRxjPP3u3eKaC4TTg+JA8Eynjcd2+Z1y9SJTYCnXgiOOGIqkVQE0vt/W4wl3GSXej6/AIMmNi
fOQVG97L9nbT6RzGg0sczWEW1EjHEQuOGrLTCm548WonR3M+/ztNSJjYwVIhAVfEhOrGQdpkjkB2
/5iTUnbpcYB7HKWpGwO6TKPX6qwtr2xUsnRVropl9HV+mASWERyM7jJw6yY3gmkKbYzwTq9hIdhl
05jT/F+oudUkgTkhCYSxYRRY6s0GewimbuIGIV/bPuCcPKjY+ZHpufZG9PSiXaGQ4h5em6m2zBnM
HRWGEcmFCz/DETTuCAsSjkVs3WaFTk0gExCDoKHXKQV4/8f+ImYFykvcI7pEenCKcLojOUb9jmYr
7F9Iyc589KaI0/A1pu1s6jyrbrlvln5xUCilQWCHC6nBu3SvddREmgDU2I1MFiK8Z69lXq5igT8j
OlPuhcBlx08OnvmgblOlbjhdCu4LlfRlaUkfVQsZKDCFb3BQL2uWfiY6aA+AjFHjGkfMMAiH1YLB
hW4YsHmFYc7qL0bFXdqyv0f5RdabR65szPEYYJDOp8hBl1H2EwRzUOdo2cBSB0cwzYxrKnvNUWmI
6efYZ3zbXg8d55pCCIzJ6yAEn+WRz0556Y5xwnY7teVLPEIHWraMThe/SL60sn5tuhb3WunKrSBp
qkzAo938meI57e68f05uECeHvsFRpv1+suyGzCSaUJYrtjLI7+0XT5t5mApPJiESsdycUTtztXps
glJRaMLeYD2z+FJ10ccBYZjqLvOkmP7N+pA/qzTdvbRef0z7UOEwx2itwv5ViW7Dq2WYDV2cAeMb
bcKNZiKj/QucTC4u1P4nCQaLOhfUdf7ulTNGaTCL8qAI9BqKfN9KNZjfvkWgSJGF/v+sy+U8Yr5t
1Rvh6/jClp+47NCeVE+E0vqHYpYEoE2VGEEeu1EjgqMvay7jGMK4N0TCw6NFBPPemBC/AlLBqfaV
3QWG1tVWU2BgVwL0zZK3OwAjHuCME22A4U0q0J9mlFhvNpiDrb6ZTCHak7VMqOByjcBgtdBa1wnU
DH9RSCR7hl8Gqypd2vneD9oj4dwqBsgmXWcaMXBiEbvflJGSrcYWoO4HNnJGcSSk4FQ/ZQzRyTsw
/LmvRjVqWb+Rsh6VLkM8vbYYH41nnw8/5oX2l4jNfzttexlSKQN0h3+ZSXfxWpEglHHt/SAtZrEr
c+tQt5NVrvaiBe33aZ64g745NVb20h2cD4O4N8TPPeeUZee14ezxtxQvPcY1G+iBzHuCWYzS5qXo
7HnGqeSDhFkhyqbrOjqvQgQoItVE2FRwnad1vPvSChpg8fMcMIHT4dqN5q1EXAIej2LrkaE0FqsW
E1JFKzhGYe9/4hRxZuVMmgWxryrDnsfdU881ce7GfBAgEQsV5HGM9EyfrmTAH/e2qQ4Ru1XJ4jag
pr0PmPFEgr8PF645lImB2enjHDWlkQ2g+9jgRQ6c7ucLgr9QY6L1PYql8k9BeXttKfVHZ7l78Dtp
/VQPp0v2Dgd4zEmRM5vuBBRChxXeEMs/uI2TUVLpbm9K3aqbQ6Cp/fd88eoOYdwnsPjJYhbmg4MU
nqlx4O23faxgyDfkgFr9D2YRbUbasprh3nsDIgQhc9KsyU5C7lZIzsEgeh5NNOwGDM+0bZhAcrOT
Sr1yZB2wER6/IiKVdRiHyckH79oPFjrQtjAnMPm8dsFu3Rk19MCiTgalw5NY8xRl5P2VQkjPpNYz
De1drTrrd6CqJNtvAVXEujxUnsV/u0hZhHW0tN6iKN0kl8VmS60iTZXBZFGpfIGdr9JZs4MfwNOz
yoq7Gmy/x9VF3xTw7WjdbMLVC/gfW4NdbsOLgmzFHF/QCZkGY7WOtsE10wHMEPhLEnK8BkxcuChG
SfVWkmlpgvEudhLzYDlFjjs/fU2zgye+Ea0GSWWMF+d1I/MypT4Eqi6yKYCuQhztOfTFScqM460h
DVRUTYYSSwCFo3zsu8jCiANa6cosmyFdJREvJNa9IGwL8obcziIJgRLjeeBH316Jpt/QYYHfJhWV
YXPT/pW+Te2hvyHtfadnUnHybtloYb/3yg9mO9eJHf8gqxaoztfnjolsyrrXKPn/0hOuOJqQWeWu
6OhVOKoENC1m3mkdqEFT1qSNhh/zg9sobpt9yueTchk2t7RQ4vzOux8Csbv5k8o/8nPMiMtIPX7o
yJhBHsMF7rmbdLIPpg6tS9JPbaT2Lgf1MxvUtqws0+bAVDmwRJSLMejgRdafr53PYr9tcG4thqA7
0n0RGGpdNjOaAglr0UAL2rNDQFTeb+DwBbegJAvlv/xQVKgSJU3kj2P/rt53O19D4Ia4FojxxZjK
hixM6mWWcSPR67Q6jBb5s55uXPWkZxA884kKM8LmUGpbdWAQwduIPEIbctU11w2n1MK7Xkejqey0
+agjx+qon+T3kWLj1awpmf8VVTAXyiZOe8fG+sj17EhSQbfM1A6H4Emb/qVvfnJ5jUD5fwMS+Han
uaM061PwfFsDSaZE2ox/CjpMD5d1kudG3B8A6BMXfqsvnKMg7aPZeZjwOK2JsTAvOeHTP9l8axjP
/hDYBfQ4yQlOjunpaskSR44X+ozPEGd6yYBN/secrz6nrfS/ZLctpqZhQHau/8OUlYCoC4K67RrW
XE5ZIO1hBi3EX4jCS98URlPNXSKFyZB0X3luXeCJYfye9W/fHUm/Sw+5tXYoI8+Q+aqQr3ii+kw0
OzlXkMF8aiq+zYwX/G6J4xtpohJt+MUr72xaAEUaSxHDZFdi9B97pGSSALTsSt+DKCanuHcUoscQ
tU+jGesfkHAtvD5unTIhWYy5abg58T6bYeYwBW5ih7nO2rc725Dmrv3I5/rplzKwTnc3dGwk7pVI
zB5VrPb4Jqeq1HKxIQT7JoSA3aTFO50FmzXxfaShrdR9yZSZ9uV66Hy/FEH5qjECWgz8NemhwnO+
jbKy/cgMCfn9opYSXAgGauBdgbGROE6sNrlMvdEkgKC05Mx/fyTzPHpTO286X+PEvNSX/JgVOkt+
uhSpQCbOm4oB3KBkvm4QoyaoOvNPz+34Q44x/Qy4Mha5Ip+XWZJqbAadWedSrAxVDZajXXuhxftC
HylchUyAFR4mpWQOPzwgRH1hOidVQz45irMBfBZ3B3u1I0/AqMa/KoZ+gENODX++UrVPBWHTYBRS
xJhfAmgk/VSA8WLgUJDuEo8vRYX2VQqqk8u6xI7pO3Y6xptfIMtVseCuauHlhvTND6tyNr1I+a0n
zJL5nF1yYDu2CirM7iFh/okbz4mw3nDirr8imrSJWDRmiaHMTXSP2bnr66Yix//t2mEYYeOIx57H
/8SeKji/hhjtAlJeEPZEhLtFFNfgZONcfFVM3qIpWotc8AovPjGshMpOcaA5a0iQl0t7UsALXF+q
WvrS8oyZsNYXlDbNhptFUSGKixkvAGwd/SKDKMY1iGY9+gCdkab23rPGb+o0x82JlF6fiKGiR5H9
nxLmM0db+g8rjl1WQ8LDWjvTILE3B4L2iexSCzRANV+CnPJE5GF/YVfneo5UIKI5VNp1FbPGEP4Z
dyPqjkHy9Zm27xFfS3w10S7tVPRI9S0y6+Hjz4zHVAiGPwcm+zCiV2q9l1O14fYvM7Yfl9LocnZy
pPElqvvHQa1ML1D+hNbILxeodR4JdGGiGiDb0EfjcuXZzKiVBrdOt/QLbw0xaVTnXgBMOLuAGUhU
Sf/D7wA+OhIAAkhTMCjgXMLbu+kR8Ea4AuCe6moKQQ2a94eoT3MCQp0kmXiRzZJJPrn58sTw8RuL
jvFT4KxEHuegkjEfxRhfSV4TPRoLS+S5QB1OVcfnl1/nrWyyXIibSwS+0uSeFIS6KwWIh8kyj8TM
kO9oSGHzyR4Cb4/nXVcoEQnRElURxLxY8ZGgbjhJLMo6dh6GzhzDsoXdkVUg5DMRDloZ8Tp7l0rU
OtJ1v8VHFcQVoVIPZ16AY/4qXe8eIYuaJivCF2P6VaTVuMirLWuQ67VRWsTdCVuHtNDEUiTGTzmv
SKd4Lxs46BYA3VyKF0TQEPrH76gyhEphuggXQcnpMq2jO2Gm+vI1AktPvUz2fG8lA2a7KZhhLHkx
Lb1ygoFt/sBxgac6292Tham3T6R5jrgAMAsZ0KvF7R9DrXr1Ndjbg0cMqxzOGefWeEKcdF+oGFy+
wOrXLbzX665hx4valJAwlmAiKIZAnAm8LjaRVC7SWCp9OqW+b1kJ19929/sqB9byOMjMh1mz5Mlv
K7JcF0VPsf0Kn33GwUE56Ofrq3SBRECrZyuZZtvakmPHlbNbtm9YNJYLB3IwDTBkAMVuifzR8wVb
rE+rZE0sXGfjG8adD1wS77/8oY9PRvzxtt+0L7xTOgSdM2uMJKmto9yLSsrOeGSZ7kby4PrCpFic
kn1iSQieYPgVLhsCAmvANXaN4q3iIaUBMrcCr2OTEmnnP+CL5BfS1Elwh4Qn8em733Q4fPkzIc/l
o07CrNIIDlm4LvObRUAh0ctzrhMD5fmwSoZqK4abF7xW3SPRBvxnPewNB+kQD2YPl9XPp2BDRPsC
6Fn9xZW7vJbVTsoWpJNYRh2y5+ADyLno/n+ZMmH+U/zC7/AcDGGYxSQy6Rwm215+/mJxgnAfPoVh
UkoAaZ7JoOwQKK2sdhKhtznSfuQDZhhskAm/XcCxF3hbT7LbJadUv6Iw0BGX5qxn2obvPu1MR60P
50wJxBw6YnLRMKAQHb9gcS2xEeCo8mKhWDIxXFTm5eYJjy21GeVBwDVr/xiVKtdN0p2DGoUATrQx
us33z2J89LBQTvJTI4oAcx9+w90M9Qz7rmNyOZQKu+Z/TAq7jOC7tdBA4p/9cCOFDMVCcnzkMKC4
Kkyi1Ul7SAYxQFaszCr0SvxQSIJhWJjVZYoZy873IHep8vddOi4jSehLRLcRVMuWhQnq0nFf7UE6
/Vfh551XzxLZNrF/Y4dn9sc7NesiXulRUeMzmausI1aSjNVVXZgdUmfWpR03U2jM7BZytsIfucvW
7I6b59A4a0vbeUgEQIjLfhWgv6GC0Hf9+rQg6OpC9NsBWi1nz1Jy84e6igQQnkdqUuAZ1+NiU/m4
2VLMa3iZcyKWB2gs0fbF9m8MpNii4KmcBkgC0BdE8TE3mx9tP7oqBpaIlXN35ALNMNz32knv9WuB
qFiWQJzhbzYYqiLGFXLWqcsTJ1ZZ326hRkZKqphtn0S1g+eJSpa4w9ind5tqyu/qoWTqTlkGFUxB
dNPjXrKbAaJmVeUQqC68rtfBRsNNrY5t2MpAzsbucTcFdqZuSjAoruVWDAAw5fV34MShkmzjFFSp
5fV8rsaKmt2enXkw75E97v2aTKvXkzNJRj8d49n6Z+E4LO6I7IAPLEgW4F9J3jZc2JIpQj3PM2QN
tyS1Q7uTa0CKVWAaz6GfdclrM6X4EQfknDl7sfuQ8343tXPei6TGpW2kTbv74GLCmoSDz5zuX/7s
VznqGtZyu/Z2LsU6E/nIkXqIsJ+9+dkf+w3AAQCi6FjG426Vee8P5Wxs1D9E7yUYa7Ifvrgp5JQ7
fMQIFXOL00J/9oxnF9jcIkaLuuuanEabRoj/8NEK2oYcIvywl1N43m6f4YxUNQWh5stJregdidcY
4XQdcIJ4rDm8QL19VlrgFSkX0BtaRO5Ecn7RNwil/H363bSTHxCVWcEorzdh7ebVjfgjEdzdbIOT
bKjXwPrRwmYUdj6IIImGuP9kdMIrm3dJc/h3YlgEVuYi64sraZWpDUj6Ulp5+R+KrABXS4rW/IL0
ik0gW4JbYzGSTkDZWQER3ha0olVVsJ0eW4MNVUe3NsR8TNkjyzRrPjP614RZH+UxnyCg6/vkMGrb
Ll0Y4yIxmdi2TPD3Z3BngQhy1ShZ9udMcsUfiN//wYj0j6SUUKwln+GBu/RhrmwHb87y0cAJetyq
B09dgpgg9P/2ds1lrp4SsQa/4+/Dz/ZyILvxZwnE8dWLCIa0dyNPmz3dAJSP/dJej6CEeGtGNJHb
B6YTgO/hcHvrHzJh4QxhFNJNdTUsYikbSt4DUqyIcs3DiduCP/gKUrAl5dXpxE/3ZMTOoNrAYe1/
NCCNDR0vApM8UcHgwtHokqSxNrxUb/gehpOQom5kjCwqs20QsdTlfDGeA5pFgJSECnLc1I4SsbAb
vNMkb2U4h9j+S4xTX/4ooxTvsuTXMi6iPqncDsnexctIl8Njj7LYkNx+5979Ev7Okh4Ka7DcR1JH
Ru88wbFSaVZmz1cV7M/+ObQbDmRuMoNsiBUGNKYAhllRfBjHwJLExSXPALjojgo3ik3E9k663VWY
wYezvM4V9aBQrVEMLUZ7HF3nQAAS967esC84RXul/+DxQ7g/p0KT63z6t8qNGXz2TWCoga4bgEWh
063bu4vkHQyAeh9Ap7HXAE+hPHlhflvvnQOU5bReNHAOWiuoUOo71pwpi/O6v/NeDNYXTvIYsb5b
0X9EreQJv+fvO2iU38uSpW5ZMqHylFd2eJAfdvQ6IGpc1rjaWEMGfGByPi52ZC8N7TzshhtLFY4s
EqJ5zW5V466t3SwZ/lhaXPBhXrGCNTluE8sFVWLOZ32s2dOdJKxIqdZUv3qgftRijHW4kZlkTXf2
zIOZaTYUt51DhRx1NXTOjF6j+Mku9qTEPQVb482HrJ7FMBYmWhI3B7IkHtSm5tXFwCa7M8aLgjHK
GcjDqzl7OvhbmtkPfsa1W+0664uala40kiLwpuoQd5wIRLgIcL9nb9BXGI/62PbRmpnVzCRwn2Qe
B0dTU4gBzSr+b3ZSMtTpCZoXJeg3kjMgdCJckD3PN9LbUaH1I0X9hASYgybN4CsrClzhi9lJIp38
VBsFHdstWj5uFsS8LRSzg49VweFMZPQSvRxBuVgQQS0znCOv395D1s7t2C6zkVlx5ATaLTNNyTbV
QPq5Sgv0T1Kg2YxNwi5MGCRV8XfglkjVDBvkwOB24b+rNU0LNSNc9LI/5x4pRZtdoIfwzEM9D7bd
FT3p9Mzo3DKgBitVJfDGV34YXDu0xbgM0gyUiPeTA6WdQAn6IBkgP6jlEOw/u/FH8bOW9geg0WO+
lRmkNDXc5HoucyBGMJKDY+H9/Vu6Bogqf8I+TWFtak5KE6P0tSH0h9JAgC/TK61hHpF490wQ03jm
FAgddjKKFE3F5WBTGbKw4te7QCBZaiaR0JI1hfwmTH2ErSAOBtjb0UnPSH3tde7Q2yKsNCVh2jlZ
URy8MkQgiE9dFR1zwoy5vCnNR3xcvoWH9j0ZxpQ0fAPXq8s86DM0eNvlsGbELOQAR2QfRjKwtw+x
0xylSfg16qf+wALAoaJr3LvAcFr9FOSerXzFPWqdnj1hhTK0TsAuBxZ75iebxlWvt847TLYFRI7s
HUdwaoWp7PYdTxcb9iLlRcRHWgW6uXXkP7mtiet8TaLKNRjC17k3ThiyHt412qLMQHAmGtHsTwBN
WEthy7BO6cfVt4WbkITYMy/sciHeEXwHUZLgKtpsc0sVp3Y+M6appuVW9q33mwbutMC2yNDsL7Fi
yX/xlM+cgiTyKeTvaFH7+ApEwLUPE89N3eZTj8n6R5V+IsEaB33+CbTMtQJ9JFKREMPZazBq51LT
460FxRtgtIELSLrMZwIMInpMGUJS67hxEK5UPl7VMrAfJAZUCjo45a/huvXsfrg/YgTX7MmXemdB
+geOeZ4BqGouZzjXUZoX5rufmlKrl1dcWFQRXZP0jT0srssh/ayU6fHxueXFgG7uOWVjK/DrC88B
x8ry35IZs3+kZRa0LP4Hq2B74vTf9Sl7N9UMHWg8H6L4vG6dtquyhD4bdTNtWoESbVUDhi04s6vm
MBzVkcoeCqcpYnaZ6ISNR0m84+RtSvCRS0adGRX9/CJuPx2rPpq9Cc1SOIC5DnWqWhBetIzeI2DO
X9ALGx4dot75F7GvfCoKvh3OfpXbW1ocXET9EPkSuIwupwmnvxP6lFM/HTjgsIIkdz/nUQ1S+juo
8agU9CfIMXjWJZodse0/dte1WR/VHuW1oCO3sBfEBW4FDSqloCCN3gQmFx8WYVOdE7gqBXpwF6ij
sG928eYwNQ8I8eH+gcHqHYNQASZsCZmUPL2HES/dJOo9Wjs9jxhCA/XpiRuhrEE7vzy6sMzRsRq5
C5V2FBFWW5XhkHNryX2IGuDv5mvjzLLe1m9WO4QtaT15SywS0Ti1c77Q+JtwvNidJnHBPxgmSd6+
BZrzRK04+KoS1+PPK1LdKeKKbW4qMW8YAo5PGUkYctGMpyTCLQLRxDK0kKko0g2WQMso8+onaheK
4WXTm0ENRtSIhaPXnOqjNEYtvj24dg+eydQHCjObbdZkJqJkTsliVQxU/TTFwh+JUOgjJz6KzI/M
kgTn58MpSozatMqXNj0KH+DHz4/0jnpbLPcxIixG133EcT/8431OMwavnV/qy747OVqSC1WT/pRa
hXaIYoFF1MG3toP6WVRqJQHFFU3h7qR+1hSbe+tm9MoHYeWA+B9hLkQhNnbH2xQeyFVxxeeWcXmo
4AePrWUPPPbz27rZMgZ4/W2QjsPJ77iHI/uUAjgVPPN9vGR/dWEVDv7upbIA2ax54AQ9V8gaN3XS
yLQEFhKmkjrMwGcKnCBJl8CgVXC++dpezm+mW9yRA7a283BwkfcxRjSYYjrDvlTX5xmz1FCYiZCF
tEfu1o1V/6zbwxvC9IUy+TvgswcUTuCpRyCy/AaGa1sKeE5taqsce9tRBsn5CbYyZvx7j1k4mdKW
u18YvhelQDEKCTfDFQQSo42NY6PGSL0EHEXfTDaSas3Jj0KBuc0MP/uuK0QE6AJ0ZZIXKOa6Z/wP
/vE6zsjAKKCJzss5UnpDsc9xTvtK8mY4zvomC+WlISDZDLZBdndzSU5evUrh/Za8cJCDcblQzMH+
geJI6MP+RwGbFkFqAxHDf3l/VmnjNJJazlqldwotHvoEAypXZqW0BjvD6DPlArwt79ipci3npXFJ
5XRhy7SbdQ/oEwrK2enlEmCgPoyIVxbj0hX7eGqRVtxCMwsUCuaD0eRJJzT37JwXy0DB9WIn3kmq
p8W/6XnceJ9Nja8z9W4uLYMXJMVC+2ald/qI+EQf+Ya6SdkQ8H1ZQP8gTr64JdLaxAgv3CQ2Z8nZ
ILzq4NHKDNEKwNE8i9nW8ZXQjO+SnyVhowLuVphaoQGNIU7JcgIeD45PcsEhY70NehLjmqKf11oa
0gNUL43Rxxw760Z6U/bzTOPGGEMz421j+PU3T9n9YEWphzRN3dPsazHnqH3VjArxoT3bjRHS+Z+M
TNVR/gm3XTFRK1oc7iKjg6w6ioCL/YGsNsdSkV0DcTrjwQ7n2/RK0Jmqgvh30vkbAIqU1BN7vy08
L2OXYFe/2CqcGNmMk/ujd5mkWai65WYAZE0Og9CDRcLifVlPMZB+4d2I851pgaS/XGN84HH/aPYq
pKqz23P/UTb4V8RwzVmaFDok2tQfQZLPc/yzeiI/wcu9ebhq8nfSdjhYbVG6tQ7cgqnjWnMEX8bh
ee3M7BLsZiHK1m3V1gm2gMUkwXZWDQsbHxXTvkBm1mEYkIv2ViHP4YAxYF1PfwOZw34eRCJ4zaJE
E72vI+Z2ZzVf3IyzAn9L+s+647i1WJMPM2nHGxn/u14AdL8q/1bDL9/4hr0sfdMHyUzhIK6JpBFu
9jLx/O9z4Ft+cqZXAncab3L8Y6PxBI7kE4Ucvp/i6xV127bHoDoFX0INOOXYoeEzE8E+EDdJiCJZ
s4yMz/4LbH882SewDQdacINoWAUDHtrPKj/u82/5h8NpX7eB6JW3Jk0+sqaNiQ/IJTYVXVg95JAh
blTgUgWXxH3lUuYmw6U+R1PtNP7TcJCRHdtMv8Apfpm7fVnv3BUGjKeMtx++msbz4w6+fzUhz4PM
JC2Os1PXSTO7GwK1gMskqJwSoqmvBexPydGjp9jHYXZeAf4lYdDzpO1jKpC9++GPw5c6u1yevh6A
v7kJKmbWogG7V7jBG3ZsLtpSJiME/u26SDeuzkBRkxNV6uxxLmXVlI2Sq/cHjMyIp8YRy37iEgpu
+Ci65Bdg9BKltz8K0yWYRonVVQSSe62BPqib0cc+dgIkf/u3AqUkRXoPWtK6/hAUyt2/kRht+VVq
ufSNEY8I/xhI4aQCOD+zmxzfeoe8JBdqlP6JzyPNjqL9UX+/zMaRfyt73Ai9d2crL33LiElmy6tF
neO+hS0ACN6NavC2uKaBDxuOnNnPGj5Do5O8itkuUFclGJ55DvaafxTODZe8RXnE0aUq6jwRRMy1
BGBCGiohbn7llO1tqYKBK9xQfK8MMWe3IzwWEdiO75bgQhMI//WkAVHGS2kMYm7Kbds02B2iB64o
LaebDinihjlPvf9GppWhzjL7L9Agffs5hxJjAQRNTzU9UN/1LU8CeVNZ5rO6vHwKqYAx4bs41ud3
NDLXT9EOZw27MAOlSOZUL/xG9zcp6uohZeghpg4an406pAj0Vzwu+1n/zTOQ1bBt+yCcap5eGb/3
+zG56sGyRCcKenro4YPEE7YwC5WNHgczC6X64jDm4AyfVxXzeOgVFb6yGjIlq3KAXkzY286tK5Uf
yRIyi5omP6ie6rZFX3tOPejxGYfuZUjVe+WiMy6auoEvIhn7Px4gITxvb22KBslVdT9JjyceYC2E
s7Y5lnY6LPgYggvKlFhh38fUJVDnw6NpUplK5D836ROEwwY1VpRx0x6LAiEYdp1s12ycS6mdcjM7
kMZYvL486kU7E37nKipoMMx2K6sguI104Ll9wcUDIgaLPi5EbznaQ/Ct0qreWQz7DvHRKkbkK+h+
qIEAVEtJydP6fylWmNi6MKcymh+0QK3H6TFSk6FrDIunr8ZMFHUnTdm8KOAo41rnClzwxOZNNPSP
iY1A9QyO6xt3MB8Has/a4hlyeIpWl6/xEWMGtEkk5ArpohxjbgpCPS0IvSo5vxTXMa/PtEVFCb1a
P9nxR15QOGe2FrhZ86UYgQqeCQZE+pBCHj+OeKtPco837ZRPy3igtS4JQamlNtNJ5f8ztTyUd7Zy
2jfWBOkhcf3sn4aqsJN0O4yxbLXGPQetA+jBD2T9xCgpU0QqkRUBTYUrIg4uOteXhZJYIWjTmBBO
R87ZfoRKuvi7Rliy0PSas1+1B/XjTPa5womTY8NlAacFMOs6y79jxTsBGFRVUrWQsS0XOjZT6GE9
mP7fevndOZq7msq5LjJlKq4z3tneqvwosmkNhbrQN5mBRD4P/OPuFYBAhwLeO5GhoxCDV8LdF9dy
zIbcDkqqJMv9KlynoObbB0wzAu+RVj/sz9eyVgZFhzGLjFNxNg3pcAptl3FlGhOPvIVWAjfIO8Q1
C9RW8xRHhM5hqfnUy5m1dEqn9211zRPYwMHOphsKFuwr4TmKZfpdd6FNOPmcjy8WsXQ+YdiWO9Ft
AIXLC7WKs6qAojm1dnKomoEPJ2lz4hEmLFqkeJYqZoIDYtcixRYXFFzdztUrKRCMjC9wkzwx/JYW
W2tVqIsm8cA6jz786ruE6oJ/rMpe8+V3PQ6i8TJsyLttyygd/UAPNwsCF4y8rVNuGSgB3WZ5AMS8
MRxJ/LrXjmu7E4yaO1LBvFB1l6miwf2aOWfTefPSTUN85AOQU1cfwlSlvxeew843aq7MGLKpoabP
bdaJmDO0Wx0lSWe/TGusjpStrJ+bX9iJWGj9Y92wXQ2OtzY5/vlYZnF/0BFBq+5AcCxTMBYGoTH/
acIzjY+bpzOi+I1zpVS3LwyUlB4bGbBlU5JcmiFI1yhtZSgOyqTUDr9gh4HQeC0Ifvi6CFPYMlyb
Lc61Vcs2CbVWBZdFUzCanQ9wGeTMbp8Z/hMnvHNtWyKQSwIpLNv9LQJPqsvbV6PqosvRyOzIlyRr
ai+f1KMWrfzvHKXtb2eKcpBn4vNTpX6w9Zidn4Z15x1iTS0ENCB4PVwaoFkHnfH5sENP0FE+8fsM
95AcnGdUBqmmzcr73GjaydZSqNJX3iQJAbn4SyBTdzFlqG9SDWQKelwcnttMKOplkxYiJmnde7KJ
Ho9W4FeDw30uCctme+xsT4a0jAhfQONAvO9t23n/HmRkQhdaOdLA1O2jkrmZNRLnDXX2H3+oOysp
sDS2TamgXqLwJvIvhNyYksvlbwXlgPsELqAa1hDBV1XwdhCtzz1H6f3FI702zodMKhM10ThtUDT8
mfmjgWjdCVlSWHS1migA7JLR4kg4Cp64td8WzcYjOXWVtZq7voAgoeraxqiqcr0vnRAH9Fqc+jf6
W5PgCIYMyYwjMd13PDI6D3Bs7lamwczSJ8FX0Cb7V96zykpsRJuK9I1/99Rra1w/t8+V05VWNr12
hLy3hdHoYKSqoL3/vMonr9dl3K5CjvOml9L+67XwXGXMDJJLb96oAAVQ8On/nSnAYYI0x2Iinb4A
7z4PiL7Juz2+sW78zk6HjAirq49G339Sng+XLskWWskLHAShptbXOniLNdFrv6+h9j4ihiBBkI3g
FOvrMOe02Gj9mutx1NducozE52aNQ0APJcHeReceFlOrUTnF9cfkluYyJxejaffgbQ4HTr7jYFCe
YBcBX10CTyGQ0nwyUgo7AEWELm9gFc6Udt3i0T//aR+loo4ijcNzGK93hTJAHtAk0XlXkKkQsCah
dLCEDHd8zGWB+BfeNzEaZbXS293CR6ofF8BcviLejH7y0rtFQBs4bbPbR7ntqWKGdpkYEuuaKFeQ
yA2+F/sk+U8TaKppExf8x/BN3knk0bQuDHZ7fRuJE3j3x2V8LhgClCDyeJe2hb4SOmeyyUR5Eua/
DUa72K8KWKlhL81KgHh70/1fwHXwZ55vhcVLKo+Muf+IE1jY5DMK79vDXKzY5oCDkAr9NP9Zgw5E
XKAlmQfMSyl0v9VMz0QkvcaGxxelPSiJfPb5wws1u+NCThQYwRyn9+c5moFrTZRUbdf3rOHSuPRI
Ywh94KqXBkWCNp/ZQi6yfz1y9Kf18uFLDnptYAEM2iheMQyzSAUQX10vTrPzDAFNOqEZV/1pZ/iL
WJqHYjVlYiHX/8tUZtKhKOm4QjZQOPAC1vs/CKZD3L3/791UPEGLUiY5TJKRe9p7zz7CycXB+N/M
05+Tx3aIlnIREoP29/1eo7Dna97XWbfTgd6PFX5jVmR5QCIY7b/nhoJuUcXc7fSD8yml1OWgXw3M
xUaXPlZUw0xqKXW5zlNcP7t1BJdOMpwDI5+bvunSGsilqucgnCFn15F8CZiqpYOarkkuU3w2jF5O
qQsQur0QaJxCvP1Srq6JOiDFNJiAwkEgwnmrhnTizfNaf/6cDnie8ccED8xVyh/75+zDzluuBrO8
N4+8MC2VJelr2MEBJjNPBVp05bKlYM3ITFu0aB3jBgUnMeLs8PQM8MhQFHcuOunE/Pvald/50Vq8
lpog3yI0H/D4g7Pp0gFbOwS9DH1nc1/hjEif2/uX/7AiCzdk9xgjUr3ARdh3iI1YB8TNcwBzA5eE
+q7y4tXgm/2iZdZab/74KU6ItUm044Bpb3Czv6s9KrOlKMbBwgI641aGacdhS4SCEqtCxbIyhNKG
6BdBIadYFpbVA59/MaWeUFXQbDPc+TyhvD7p/pYGIEEi0UTlu/nndh66z1xctPlA4VV106eXIL5D
CUP6jrKaD0XwpFP5IKfsB+UptCW2/r9wVUoaCgTBW5o1u59nv0DWpVIRHZm7eIhvvVDr5d6Mr4n5
f4OROuS6JAQX534/1FuIlzgW5ftKAR8l11uKM+LZc9LiXZ0wV6j6fDm0Y2r83oy6pKz9MPClLxVM
fY+hFQ6LU0G/b7gvo2ZYiRox/fDn/Au2JksbHBWoK25LS70Jj4hEReA9KgzlCt0cMUWoCyXqQwsS
8bDHL6QH2yGCRRGhGENMEEyRqayM1DLWWkOOe9tIIH13Z7l+TLUdzVC0LdBpokQMmaQwc2Dsn72E
BIgdh46CEg4VR1T7Elo75OMivk45vzTzOjde0DW5480vJo0FfPcYcrqwiTbJwx68jxQjPsXZZtdQ
7fieSNg0Ctj83IeKBKT0f0td9tjinmnRgASGFCjueENETp8lzMUTG8NK4ldAh6ZyYxmrpPf5qrdZ
X2NlUk0ToK5JmJGMNQQgIGPfOnsbTgdSTzzlRXodNBSvijls37knblMABinDY+NMGAKwfeJWSgRK
YptGE1uF+JVX0o3Odel/JB5/kMZAeJoyQXAwUnhPtumzcobjkoiLa62PA+y1UjsPv8ArxUAERQN0
xcCUzs2w7kjSo2dH1nhv27oYQf4oOkUogC95gr+gc4MmM4mkelNF8Eq5DYFXIkLq9KWUFUMJlfeH
x+JE8SoH72m0ZkyY1hPYrC5VsNax9ZnZSF4qX4EF594cYKpD1kuCEXomMW6gRuWJmfypn8a56yk+
8hiGBPJ/hnM/wZyVhdDNB5IXSHlOPsjnAmsMt4wMUegVV0jNtlI2itNWPA7XGH4GUHXsRrP8xWd7
49mW4fw2Cz778q00WACqQRUxmeD3j7/mkm4UhITJwELDbmKL7y0WfbAHfmz8Z4tAFa7TPpYUIAOt
6XiFJyQuLLvckJ92Ps14MrFYxo/8bkvLYEtB2LwUGs6yCkeR/MPR0rLQseMSdvWo1sPdOHF6R6zs
sgXI6OKZ5GHp/FAXGaumys80zA0Goag1XGmSNYL5Gg8l1za12+mjhtcvgPefNPWpztBB4ccDQN1A
MwA14E8AgeAoRgbEOP0xkZu9ELfgNXN8X+useJCtMxYo17glgsLs+kJTHkstZ10QteLTLlx1FWei
zv50bG1Td9pdFF8q7mRP+nRpx4ZW87qtLEzIGAb1oQbhvwvON1iIxpNwoFiXyDGKOF+PkQrj7v9S
cB9kzgLA+sQzu+ybi6zIbvMLShBwwGyEWrn5n8+K5rVBRnhd2Fi/Z24KNHLATp7cde627EcXuhbK
nkiPsq6q3qXGjglEz8IQNQkhQA1sQ0H/8V5bj+qXtjyknuBaDMQioPBXuNiVLYDrrWziOS/ZMtAl
XV+q2zkj6TqvOmVNbgQgAMEunAvRiSaeogC7EUQUBfIcQg8t2C8KMbAJdfcLKk+GI0YLzJ/neGMB
BsH35Zhd4zcKyAnZ5WGIWM9HoWyw/MwSuYiENZXhAsvTyWuFHcy0QJpUCJQQeyKeCpjup/lfKNTr
+TxqTg0oV+S7E1fgv4ByyyxcJS1tr7kS5q2p4Opr0ym/RnE3H9rHAnZDLTHYuiqVYYeq63G2RoeK
lxiK70qEztQsSMxTdZeTGhIf1jSi9BPqd0GTuKklxDs9Ya2jgtEcQHEBtO9cJ6qqrQC3NkYMZErV
2iQoGJEpdIpz2ncxSGs1ixddmo65snPTfREAVu6Qc3+AlNXbpUBdygO8a1EHK4O0V+UZUEBevZOQ
YNJa6xWl06V/4rS5sADqgz8fiP8HeenAVzmvmyOi1we9M5ckwLWmAYesVm/5dQZs2hygwv67cTvX
cq9PN9ULgodVf+HInHZ5E6hAA5tUT8iwluqhBCL8Nm0uEMREft+CI/zb2fbdMycgXiSj0Jzeq2rf
dwoxRHAQnWpoTUVb7EKOYlnuE16/YTlhv2LL36TdWrczCp7SvMmODrthiToLOaDFiLPh8hQS8CYg
Su70jR+2kKHECjKKkKsucZUD9ySoKjDfCUqalKZi5k9JnPfdZmTu+UIUK3YwCiSNBcIVF2Z94EN6
im+JqNwp7z/GIpUDniuHcnesBY3/WmmcuTp1HNsA3iNtcN+wdWpEOGDoMLtLs3BSezROalP4BMdA
uu4Mrn/FD0bBlJO7XXtcQ0uYwUY25xmUxYHDX374w96jivHo+Pum1Kr57h0Xf7zl4/9Bh/kbX7AP
uOM/njpG3WCu6mUmjCgqg56fClRxnPz5iyWaOjw88yTcYDNjRCOs3sFlgUhgf8Ijg2MqK8y1NJsf
ODUhpLMhi3/ELx33KRE0qFtPXH4HP4vPIuWOuFD4hlwSQwy+yt9dpg1U10/ocDyL/DcC6jBeOJsT
W1uX58hn0Ev7w+EGh9FXS3H9K2TJC60qeX48eXmYaY2CUEA6Ll/UHZMrXMK92f5YRN6ujin7pDgu
52pWF1WVetYtmH4S2UvLKdC96CDW9frasdeU25S6Nf78i0I2udobpmesc2Hqfo4OuAWPzy7cPqj/
1yHvCIFE/D5gLPufEzsgIcQ5K5oI0bkiEQKiDHWIvRYeK3KvpMTEovogVs9V5cn6esALIUihRBrB
UqcWM6/zcSXCPlD6YB3duJBARonqAdonLgK+CzyZ5rjOwvIa3N7yMVj+45lAXmxyWGjhLB+bRTtA
oeTpOBdW+iiKYnBTSyn65ljUB0mJx/HUR4OzLHtZZmq2Nek+cVkLjbiTmZN0yY5LWwkwdLaSGY05
om5xtP5gOOJ1xTrMcmhEJdP9qhJm/3SOrovwW15aUuwt5bh0a6U0lcO1tQW7oOwWRzg78sKeDxSY
RuPODg7Yn+/X6Js88XG3hNQ4EpZ7iAL3YXsMINWKilbZB/QtH9Xe3ZEOmBc4f6ppyvsTaWsX7aEF
poFTij89p04Rv4et6TMbAr3Qb8ZkOKbxTdKE1ahZS5b7JJlqxDNVKSWbYVQDtFHpnVVRnnu1fybY
pG9r2S5cEmI1QTGmS2++hJXC37B9m9Zl/rtOjKMGu54x8J3lYlt2N2Xb1LOsLuS8AqSKIMM2U3df
9J0Lxc7lOfpJJeK0HQBVbuA22OrXg0pVL2RswURr3KrlgH9TcarqZ6kiVrQGivxYTG+FTSiC63KD
jeHcORa/ywv0Fx118eZYDYJvfOQ/6ZG10bk7X1JeffiMcvAacoIl+pooJn49uaUYhzBeyxJNPBGs
bCl/xcGzFhrfiNAC3aut386JdALhPor2Qh6EfJItcPHfOoTxK7spTM/aEVyPmS0BKQgqfWkXD4lb
M2w/Zuketzv8/P3N2tP8vL/WS1RY4kgGYQ1Fq45rSJ2ShptTYfW2P2edHmdwHOUO70kp1p1E8DVE
+zy4Ih3izinqVkaBv9oIqsf9/F2qWEPp0EetFb0+OqaHB+056XmfPns6NqncC8zYT0YUQlea7bjW
10yDxzDGfLbQJ4kZSAUFApMeZWuGV1Um5bIZfYpXA3xE63fGft/rKJkC1oIyFpMuGfLHMHdIuEH0
kpOfU0HTyIglOfUw+4sMpFyh0K00k8USp2tXl/DFE8B1sQ5nZDAX7UXBhyoOKRwJgF+KxUtDfKxN
U/GTB8vXUCvC7or7muF/JOrK8tcAeKB9nrnrY3RMcwrEdnWuNpDGUBBgDAb29et0bqy0QjgUWBMV
Txx7pK2Y+K6hjrbN2djItO0T+ZXp4WQdPzRCTr24xBA396s24/IGUDHBxcSROGjRQmHeJ6cPGyV4
Jv4h71OmcG477YX9tFXyfL14ozSmP3zHvlGCR51GjdGRt6aVOdzoATS5mCFvxZhdJo7gDVDjB5S8
AzDQhx3CASF8r/PsrpKKbFYWmYKIssFkhzNmfgG0ZgorV4qNmWfiPUxTREI6k+f7V51ReJSdczHs
dRS6P0H5dwQXvE5/LUQg4U7z0gVJsQsa/rvtK/MqXo8+QulD5GxWpxNJ/HjNZt/ePTm9XBydPlTi
awFbIcUmIx8iGOu7rpkh/SqjNEK12/DmzogG7YZGPIddnqDNxc6zZ8bHdKCSzyrSm5EDvnq77mHP
u5yc0zaGoI0L7g0kwS3hP75GIh/07frhlKotLqmgvX1vtWGNhWJJylDy2aKVsr4f4Iw1gGmSypWM
7S9xOmJCjUEeClawWMF7/4W7vWLdD8RqzXt+CammFpu64ZCPohzQUBDx2crhwdCn1zg5lS/O32vV
+/p4k/iDYAvFLJSIKcPlvUlsJpIcZBV8TeFcxJh9cjDUwuISpnbJ6DIvQWw7gb5x0W9kW7HFuG7q
pbpZaKCgPfKWS9jmU5+AGEebnnlSuSG2UiqipgF/BsExLzR7yNM1jULe+9edEM103kZui+dgMVh2
KNLI+xDLAhYEHzNIzGMezXElBpTMK5HsGFuLb9jyCzMdSwdBmjxaFUtLb2e5RREnAhdOoisti2fB
Q9UXjOhyEDfSmhVLbLIOiksNsHmzZADNOFSgXzl/88UDYGmYvuachFEmCAAgHCaVGaH0jBqCWSub
9JSUPF/68521IZeJdl3Tx1Nz6xobqvnum88emkCWFmY/i8YZFjzxLoCPf0mqy2LLtyGns7/uHaWM
vAJNJYmzPLAw0z0peoiv8+hOREmGIPfFXvqy6uo1RPClIGmnfvY7sJD+QYlve/CbQLtjExDbTLm8
5kFiYHDnBwsPfTnssc1FY7swNDkvFMrcGThLAil+QcVcKUKJ+5cBC1s9KwR8u1hwlGs3aTqr8CMt
8EOXcvYoegRfGJzLYz/evfuuGmx9FSOfLoC//5ZpaRvXsDAtsLFuqmAHCruOGwO9U19enphcfDIT
qTFkduhsTPhtw9Po/VK7Q1KPFQXuVbufUMo8+D8WjxD6R7rIWECxfVRHX0Fcx6iWnqPabslq47+7
zsHg/GsMTBs8Ylcz14q6YLcxhBQiVpgAqylV6opjn4SbI43a8KQ1Z7ZfhsSrF51q7B4wt8VlXWPn
3IiCTm6eCwzsg1aTSu96CkHMKQGPmi8aNnAvGRWFByCKd31OsQRDiQukSFzFYWJNcpIhAvWdqttp
8ioGFBTxIIfEXuPE9p8K5XEdt/3x5ObW7PHddZub5R09DZx2fh2M5dp9JzZ/ulVI88a5iUk95sO/
mMUw61zDG4RjThBmKYsN73IObAhOFwfRCcSJvs6NkdKhcbdZmRMZOuwHN37+7iUOq4I0mhST/yuc
oXd76NhhTsFwi3ae8mtagCTXKO+OqVaVWFmMr5jL6agT+F9wmljbrTakeeYzXvyO/PxmBflzp0Oi
zn+IJmiRDAYbmxSyq+EV7NjVwgV9DhSracnFxTWy72fZaAThRPAIeTYFARstNpyqXqF0EHv/rB+I
CIuOVVMESE0PMPTnG8zu6/0YgHqivb5Bki8T0le96OdixtFGm4EcR+kJtfysHTjdEhhvNUYB40Lm
ZvohH17Qky6Lg3ppzHMgHkmT+maDAwMlpoI6nHGr9bVhadg+vZTw2ULHfVjt2Xpt8sNsXgo7Gczt
irld/toX0f0admML1CDMBxxjouOqpNH8z/h+KMv2yhVAs0cPSMGlnfZBSTpEcRLTyWldTRcRqVwq
NPVhMmc8MnfpGG0MIopbibR5b+JxZ4Rjssrk0HdoUHnjr1996z39owVQSYAPzXOAPhV3Y9N30fJH
U9MuoKMG4abWX8NYF4W75VS25s9iIgqy905y763sy+Cdo23DCC51f46V+jJHbyQ3LI8KaljJLKM+
xgOqThNxbYwfGJUNLJBauOc6RVVvTrvCENIDZZGLSWc7s+sStPE3X+qkfZn6bUG/Qlssy8/4/I8G
tiuWzExV0PL66FBULZw9D+Xg/pBaEJ6vymbOoxddQgZ7zWNhSE3Lc3PCG67GU/L7WXI7Ld9+X5z4
YL5UxYR92wniKb6aDwA8lb7gY8F+7ZjjGZ5gL1ACmK6wwQ6O+0UCCWfoI6Le1DbPfFHFTqa3WqWw
FEhxGYTB7WHpk1Jv8I5ivPdcEBmZIjduBQsfpaaq2f9kKdwiQYCpEbgxjRgyEuBhGQoiNYqcPKnt
IRY7OpTpSaR375p0OrH/zHb6fGfAQKZad2BQB13D6G5TF50oH1SCMmgO9ZXY9d4eT3GsxVmzs9J4
P1XFPd/coTNTyHMO1sOJQe8uNDVuBUE4b8Fs4eRPKkr9sXp18Sz4QKKxO3PlAUFLiXIE24EtnqSf
1m5SFO7OZhmlnlGFOq7CrXyoodcXzXPuxqdh2ovpPptvYu5ynt5LV9aT3T1rOyJ5zcLyYtc4XV8m
uNEcSg6mg69yKUUJA0YBXjDPlkC9qHrXUR8Q8bFAbhxsJsGvDafGQ0fteDX466qFw9nKIWUahkGm
bQ4IpE/Kq7Bndn3dYvAU8SWU5p2X+7pmehdbwWqFXKxLXymaixZ7vIQ4yvTTsCLVLb7gWC0Moy/y
4+oMD1O1W4dHYtudiqCuBszgelgaRsCAXMsHiHswE60vHR3Clk7LlCHTPOo/pW9FuO06NtLHZxdE
tr04jWREpZoLPPLNOPSXKeNOIZcdXzWh5VgTkz2o2Pu6HX+wob9AGSYcoWaCqXgmd3HFULL+7GWR
EqWbRBYXwNPc5Lo1f6+64QPyrUP89AREdy2XR+aH3B+kCYNEdk9w+7oSnJni6isAeVko1vY2sSX+
Zdn0kW6pjBb8d8ZRzn6WpxfG4pkCTsu+4J6KN/HlFe3k+TsvdZbWgE1zlY4JrVpTERUm4mfuepQR
z4wZXySohaSG+F07pRor/2NzCqaanh2VAsjZ1s7kKE9Z3HfIKCCVE5WB6lS3jW92/78dc8V4vKVH
DNrNH5BGCmmW7oNno1/+PP3hihnFRdmxvDokBfjTNawGWmCDXfyhWlVT7vmnNIvrpWPwNfk9ozr9
DYsl81N5wgK0m3F8Rch9TXk3UAW5fEYefCsyn8NcMKQsY59usQiWOtmKRecd2XyUmz9fwNLEzcOt
RNO8xmI3hZfCb/KKgsSx0JZL+BYK4Zd/EQgquWOe1SrN/0I9AaY8nM4ZF3qDtWB3K8TnKZai0jBV
94uMfsWl3CIvsrvN9YzTdMTmwaFDw9CXwVefOc97mSNxzlFe1eaqEwUyILc6t35HcuFfPiRN+Zlu
/QZDmL5JPG9nMjMdFJHRm+aV7hPuQXTK1/zvearQ9MWLloMz8eCbjJI63jqzLEjIrO5hcPJCDhtM
OU7Aq4qbFEIpjEPSjmDoBnhk8SU9KsAhqeNfeNlqJJ937zbLOHJEahZgc8t6VI+3+K7h2ngcZzZK
bm/zQF6mpaLjpQwJzq/pSKPInUmby10ji5K9pa1gUl//U5aw1xtiBsMoCVR/rK4Z7m07oAk1OohI
jeicjgw44WwDfzkZz+heNNmC3R8+XDdmYKWtxNLMa32YZdEssLWhb8WIb55Orkb35Vzvc5DSsDI+
kq4dFWquuetdW04bjYYcP9EfvaaSKpT+4rmPZOjSNcC074evd800qkzbf6XoPzwIfA31cjfA50ZU
zR4xKCY18eIO7i63SIGh/2/Fazoz/Dm3C0xGom30qePbjt4RgtjLFDhq7aVLjbSBcoBWVpT6GGT1
xOg8lYb7U1TWTzIQ+6aSWOYB3/5WfWGTOrDPuWkPSCE6qSMmIctkXmaVTSQLwyFBOi/KDOXrUHF5
SczuBSCsucpr209fMEpxCoPSOJyQEy2PtAJEO/81cMgIjDnhv6sOMgtFhYS2Zr3B+gVEdcfvbwRs
/BHr767l0k3duNPqOZOjn6cFeBwG3r+e/18MjVLr2Vn6SK8pe3fb8Zjo2qnMyKnnihi1ma8cDHoK
A9CudLBDlOwT3MHvsD7IDFmGI+4SUJ1vwp7IedcRfNRpymPhXOwA1rsnSd6M/EEfc37PQhENi/+k
H5JhdFHTuTfc3qVz/ye7wC7czITfRV0+TxxXtLaC/ebChm0Lzb+rWarpJzlBrGaTRH90kGedqsVh
X4vp8gpQ2Z74zO7wp5QiAyXNSzyC8R+v/VfbJ1kFqDwvpMUeByxNa8NmjWO9ibQ0x27knRxeEqyP
g8unJ/RwzEbTfEjICw0dAUoXsIPgKw/UzuRIbKUvEmX9SnjvKesUFh6IlQtIHDf0UtpVWLszmPCn
y93f9RWmVeqvVRz2SlAxXHbL61AbyTZ7iL0DEOTHuKG/9pQLstBmjBsshu0Show1ayyZWW1Fig9/
NzKEHbKQmEEAKIQNaI2Nmg2iP+3wBRvTJr9rQGBRDZIv5bXi02lReG8A35oTJEOD8PNC/wFjzS1b
7c/bDtJwAfmWaqUu6l9n0wPZZZ2/2+QTnQZuCBjCe73n9I2j2q4NpJhd2l3jB5t7CB8vnpC+u6PP
tBBYBWnSbTTDxsO1joNw03Hwfv7Cbg9KbI6yxZXtgdKTPfQl4XYkEpKZLbnoptyaI0S8CBkg1Gw1
gaLxTIwj8xBfM5rRtyivfQamMNoNa8+BU3WYYonT6UE0tK06KE2IivHpNn8x8e3U8cIZ9RoPYLt5
Psovxnt4z8wnPEvaDOv08uUevdE1Eu6yvKX8GcQVnOS+QqU5MyUZG+AD5hu4QYcjFD3evS5xaeKu
DdGRIX1eqtJWikSO1LwgwTLe/VLZrA6jVhSG4g+fJ3+B9KUDHIni3ySk6PbIX9nLXYSvGe4r/xje
MqgWol5PHSx9R11mohe/0fv+EAaboumCDVLfCmI40kY3YlFQpmFyRBItglAeEZfMzzSJjMu0qWUB
vJx6ZNioZvU1VdPUyN1+lkLs8s5S9HTXeqJaKn35tspEjkgPGH8BQcZuzYJFxSgQeZp/KrX1HEtY
ZKfBPbS9hN9wtG93OA6RBSgcCKJlxfV+A/+x5mhjKBS5g2Ke2vnCc0xbUZQd/GmNZM+ZC0ZQP/H/
yvEmFOZXgHW48mOAGNQzTr7uYxC5QPGRZ80F6wtec4+CeF6qNfTV5MMnSNNywhA3cSAAJtXcng4O
067a7a+BiaRRK5N/ONvN/XddK2rL4YJTFWvDO6ueeUaXsoLsaAAy92TSzps8OWa1yY7WCg1jMOOY
pD7m7OqivL/Lm2wDtkvTfYxFJa7UTYR4hJinTK5+DP4xcyn7pPReue0EsI+ZOi1KoxdYv5/Gdepd
NfrRY1Iw1AN2xF0EB0HDos6KpFjImrMDafvIVF9KvupRYsovQG6B0RomL8Qzchm4WeG1ka00j3pI
I3VYZGCmd4qN1Z4fqZ3TolB0me7fNTu56lXXgEKNZEZi2u71U76NliDWobjOQ15cYBCfOqCOcSkZ
enaMA8TKaFjuyMW2Lpx/OEuvHNDB7h+Wzk5xcFRwNtdfPa3WtF1yynVwqUrZFmc1Dfh1B/qSAUhl
y36uCWD+/RTDsHpmyft/QYbwerEC7EhbEVXsXtR1AKigHEBtlZZGFivSykqhU2pZM3tHRLLQRgCb
nt2/mlqMk5ue0qkcs6d/sJ7Q74z1hxyB7go2RZ5+TITm+6kkrwB5aoABYKC8Q321ywgt6W/lXF6A
Uq7rUtAUEsPgeexQ5mt5R+473TWmFjUinQeHj0MXknrtCo8zB7OpoMlJlBLkrahp49NYAcTEoMAr
7eB17lsTjB0CPeXJU/0qHV/LJMPphz2RitK83oqzBJ/TqMxyehJfd/O2OYp25kfI5bsamh+p1aCM
Q+4jPdNazBXDNIlRDj7tVOCf//uVFWvmiIifxU3ZBbu+pffI/LgTnFwQ/8EdQBLUZTNPrAtBbfqn
V+vMORXqQPj+Jo/OXFe3FhGjU22+kIfog+BmFps/D+YyKOgLHhQ/PJjrWzuYs3nGQo/DA7e0itUk
LsA6o8BUtunl1KwpTrCSdhxLDR2izip47lAykkS4I7yH/YFp5Ssc341P9wYH4YJ3G+Fp2y/54Ag7
llVAKAg1xhXzm84XybC2Z0B0r/9H/+dZJ9aQIYWSWA14i2Ps61BNJE0CTEROp19G0bK4Mnl0l3Qo
eLzUo9Ga0CJnlEUqi03i6jyvVtxh1R4VZ7t/yzsbUQPR8gZpgw3ue4AjX/t2u9aKdK8RQ7EZB5q3
O2NEMzwXLHsRelKrQf3n+1lWeLFO+dyK8clP8D7qlwb06GHkReKe9S4G1unvF5knM3L39XM0oLOA
xgQQPKbRSiXGJtGnyWJ9JFnYnIfMN5R0rtvcIkElUZzkQ4bwfwszShlzUQaiKh2cv9B+DUt5+Uqb
nRtXEINyjg7UKX1nA/BEdrFmrcocuDltAMG6T9VBVxbe54/oRLg6vF6ZPJTClZURPscRU/PeOOsL
tccXVFTv4nFWFxP+kQCuvrkbT3yoEjgtSOIQtCEgEBgxVig3pKgjaZki6F9ctu9vvXmpAbCEjnmH
SM8bUVXb0JhjGPsumTDzAd7oQ202X4u9LRva9ZurrWLmwt+f0k/SxgF86tHlANOG1mH0HC8lPEL0
zUJ0CrnqZFp+JLZI+1HRhUmEZOfNfKK888vP3HbbN9ZUbhP8NyOlhEEOLG6GRmeOqBgfh/9aK2zG
e5DFKRCJp6qNgltWEDNODJhrCHt1HsOnep8roiyOWefRca+NEWBlhJEb6h2n8zifEH0hm377RWOp
cygy2Lh8eK0JGwApgRM+LzoiyMwXd4Ekj3qmcTEAPo8A+6Q1wdIh468GrNF+34c5HvgWHN+xzNJe
jTB5TyIvQ0tuHL5WNDfjbQjUxxxnNxhCAzB01QnTZRt76LwwXoc7fDGzvlJmw4BwrvsiGVqEIDoH
zNtzO9UzBvzDHN49shZwrPGXKDfZWc6RvgSSK6UT5UI9o/+spVlw9ew6g29EQJnYysDK3ve78YRU
FGF+M34Xl9Z6oKPIkZF8L+LSKuP3vEdDeaw5XdlSOtQ+X9PDYENWO1gL5u5EczmaBkzZTs5kqyO6
8KLBZ9Ho3weRcrBaVwR42hYOgmr37WYbx/8sp/lqXLog9g4d5g1RzB0sa7dGw65y6PRfklO2rdsD
Ky2gOFXbguzJ6ELkitfJKSLHfo81Wu9ESP1lEdlAsCDu0u5ZolcAz6QoiOXGPC063bnft43E9O7Y
fIwNufyZuFDpB3NoKW4ziYRSkcYE59wWexc6XwCpw8Po8UheqYp2XYzz3s7bfz8c6oM33sKcN8S9
u2+96EE465U8+Ad6ydJmJ3kN6LcQ/ZuB2X9Ugq94Qseby4NOm+vezFqOT11rl1ZOX4Y5BSDHjaYf
ChA354pq69KWq8ru2yKTF5a9oeCiX9E+PjOFFGf6vsjvzxqBArh/n4ifObQ+KpPHLxueMUVk0lNr
1C9yTPMv6+7ed+zicwqqUYKWXAYeYnZAupi5NkBNpPzlEgGgBZTN4+cWs1IlFeb6NOVZcBU/v8z2
piagM6DmctepBv2nAy2INaZlAYMuHew62TY94MXxmE8yf3cSD4K6Lp8MiaDqiMKeAn3xZTOW0e7H
34Y7qFAvHlwCENbXR59T3CsqHqgFFhBcu+J84MhwQEiv9jgMARj1gXRm+ap3kOaaTW1A6lK74jIy
AnSF+bUaOnvRwITWPfVKskWhVTwe5Le1xf1ti1fK4UKCRZJrSFiO0P/TCQ6VO6pdmoD1OkbdLgYd
LECVtSpq0F7d/agEqpbHrAPuPFUB5kYKgal2EQJOrNzAM+A250TNUFhobqPAx+NInOcZBo6I085a
Bvafl75ATpZjPvjl9ghdrW/nvTty+5zMtF6n9cmuVm6VIAWTiLbbVijfnqOQ+aYUTyfKbPds2zSg
G1E64TJkONqlSjJ72I2l453YUcDqdzwrplAwGdr50LQ3hzW2bPHMbV9XW7jcoD7x23ApN/cTjTm4
cSJwIvI33FmjpWLEAlO7gekWhpidKudQcTyMGoTvxO26kjn5W2mj3okEWDPUZdsviD4yoKPcIBS2
ziMQiflreDXc5oGOXPVrYgBzR5eoaksf1pyU0X2HqSL7oJHiME20ap9+7DSaNUIGKYcNClrbhs8E
37NFC2btTkROhvuJhYcSBrG4WRcvY1hya29xKebsO9jYBnqE0p78uZm2HjF/NrpXHBXDim/VkrhY
6FwF4ulVaaD3O6wc0pkpEM6zB0MdSt+sF0LbfbPjoKgHdRhH4/lVOVmBj4/gZqq9uBp0P7TzIlKs
GoliOC4a4Rwya6kQ2moRqLX7bkA7gYk/hz05NOlolU0vh3EMEv9olcI88Kv0YFH0pMX6HDDdSzXd
zdDN7x1m+wzzOpb5ciTfCR+Wc+14ycE2FZflZ0kdcwz9ZPGfxsK44PSvIHKdFyXAvuhNYiH+wY+6
og+Te3W8Y6Z/BYZHiDzc+CDk95YFDBc8CfPDj5YfRj9DXEezTCZhB5aEVTx2f95KR5GrLL+asj3x
xF8bOXBRhEWfh/lrslefnZ003GnmB07xwHyAz8KXCMTetF2XoL8DGJVoe4/phX/aqzrsIacO82rI
TI6KmEDj4Km9CcoY7gBfEvbvsUj08BvtzLf9Iw8Dyg13WEjAA51x6y7f3YZQNoxTrhcunA0qnfy2
tfM7bqya26oemf+Ub1qMRXAY1FRJxPYdnbhcFzPKz+Xxb8x1hDFogVmL8Ry/jf/Fgv9ToTKagOIC
4r5+fCK5v8frcbkGleBKlg+YEdlxWD5xLlUvR00ECNYKbLB8Vo7UKf7KKSCPBT11Jt5cHugJivbn
N3dYUqJW2M1b2zMe+aASjwCK5ZzHfhZjBEXaJqVn326RUzyUCIZFezFaKGqaRO9hxbXU1PRdamDt
rYz5oBpNKWAXAmINk7eQ7bINkBZSJmVAagEbUQH2yS6WKObQUTeSGAPbVTT9VupCxZpYZFnc8naM
9z/01yza8LGLYfpiPzxPQ3Ep9bWXCuK6uamBeEttz49MzJE7QRzKdcanVbsEHcavJzkkM+wC2YXI
06X9/UhcciNRjG18z98BOswy2UTFr+G6iaTSAyZ+e9+72ymKNVGc115aEt1TNmP7zRm9dsR3NUpz
LMtZSWEngin2dP9X0+yp3GEgy5eTI3wIwQT804WmPBGBmk+4q3vABHqeazGdS4hUrAkkwOaq78FV
4/uP0lvPzIN2KcmEdJ3jVbnM2p3FowbHasHmQk9o565MWf2INOL878K/temEL1vYr+FvEH1fU4dH
6WPzeXriEnR0DqeLSgGxV74yvo8xHJSxzh/ThHoZzzoKvfaSGkjVPHNOvpAycXTcMArCb0anR6cQ
zi2VaNFlOiU22tCI/XkTsfFn3Zxc+q7qKUINW9L6yYenayZaOzrDt45c5j0myPUfKy66qBKmHPJq
Z4pA67cQnV10BKLh95FYLTi3W1lov/XtFHlKPt+JFLRoNES0NFqsQ7vSgI+JxvF+SwkyAhlE3s/v
zTkJvsZnpHUarfrmGVD1/hvlZL7IVgFgGtD8mNXMfktkZeIY8VxQm260v9SBPXgr3QMKMiZ6sY+l
tCH0u0V0l/3Naq0hG4iqsFBL+9nVFTJBXP8gH6RFKF5m/fd/J5Z4mlBXs9yVXgUHgIMPDQVdu5AR
Aui1hI/7b1PSr7iJCQKbkNwQRIWyrf3dIrEAcDctsIqlepyTHZOX5b6r2lPyjdqIsLPKFxc69D1s
Bbo7bQsTZ++TTAsYkU8HsrYW/MtEDQpEMaQvKaVIF2oDT9fh18Q+e/Rb0f3etirBuC67bpOusX9W
loc99BSrbM4HGGPQYg9WqhkNq5F6DfB637bOhX5XTPtP0VrgVMB3ZSnxKz7+PCQQAPxDopzqfWst
Fnmu/sS95hxgty1vlO4siZcmxjhzq8b0dTmP207Y7zWQnr1cLiJESugV9EU+GxrZUlIAU+UczOpE
dPuQNYOoANF7a7deI5RZbHxiOnqqlz4eo1C3PH+l1/KJhYhWU6VIdrC+xV7YgXapDuj6qdBdGbvg
/bJ3+STfMDxwYN+ctRTSvlwuz1cqVv23kuGwXbdDqtZPpX9VqfhiAX3LYlx2T84F3j38j4DNmmuX
n7LO4tBAz1SwAy1vzcrlzc4F6K3wa8ZzvDtpteuRLDRRHvlzRFYLifrt0gu8+Dc5GGDz3wK7gGjF
cRshtlA6q3mfUBk8RI4uRpAh6bh2H3dsqFPK8eEjNVOz0PyuHt//SmvselAn8cc7gozdFdG8v8/o
bzSbq0QgEb7TLBoLn5tkNUgrG7VibYoFziJCyVBvi825ZQ/udOB4oeYRxMXeBpee+MtQFFvZKTyO
gdgpLzM9xn9uJ5/V5D2vK0D4lYun3AzTQ2F0b6r/Chvz2+kXlAEDiG4wdhqmmvGpqTt8ARVnunAj
jkAR0NNTR2vqEf3Kv2/riR9kxj8/XvvorJCwfSUeVZEoSu67euyB7KTFPR9MGgRhi3fmYs8z/64z
3RMl6m/Qu7Pi3nhOu2i3EeQszes0xZw92fRzUujDFCJXTyE8r29Zv1H6nYNhJpXY/Cmxhw5cGWHW
zII33zw8eZ5YY/gO3eMPLxGrJqEeLQKj4zKLdlmrr9UdW/UMOZuf3EN79AjdPMk3CLyVDtsNYAnz
Se+TovT5aW6J2gEaEaxcsqr82DNBZA/NpRgbwJJiajXdmv3Lqm0nFEgHsmOC7/ode2f3ejNYY2TW
jwU1RXCdno41XNVSkDAPKF0Sv36TEcqZriey9+4jjQuNk7AfJ7w5xL2LfvvNRy45QBtOZgw4JHQ/
oWSNFIp/MnUlES81/K1wUGNII0dDWAwTjMmfooydxXIwi+qPkfVNVhgpjRsMRA8nFHIiIQKIa7NG
BViIXB/pFLRBuV/goNjpWhVD1rIfQrrnIppH1pnd2mPzvFWfml2UEIrP9nbdZS+X9bSslvqGgWN0
EcBhCU2MTRwPLAJeYxJ3vBwFT3CaRXn/Yulsor8flfsLWaCkDSyldYMNCK5Z4gRFwY40EwLCwpsZ
Em/u6vL3KPaTmQLQDdNyvUqRB6OgBeFzD6oRGa5tcP5NH5TIAvY1RNwULZ5ks/zainUCPrj9KhRr
a6daYMxqDFYT3fcFWcoaKkZDHU4w19yI3M3BcHV4z9tm4/lYwkYRyqXwAJwiEsqotcw42e77gwXJ
UFFMxHHiYTOc03nDCqiQLYHMMCq36JSFPCn+Tn+vZR6mEy1AUtgpOt5FS4JwlDA6AZ0ua7G5zjCY
vqYTAq6DklC+Dxs2SnF1Y3WDIrzGACt9bT9MdrsG/19prlL+8Mksxyc74pk/wU/q6uoLqkko0+Zc
4J1VwMBIhXO3EXIrOvX8x7CNwglZm6c6EjQSRC9969fIVllzOT33ESpU8keO/nYvZIFEATulJaZt
w80BderJrcx5y2imSVBAhx9wKl2nxD8gEOd3ov3ydNwL6mr21PKbh+iyypEMAnsQMPsx5M4JaPAf
UPusBkhXxk7oFCrdQM9EESti9I0shYUxeYBlZMn+x03TlOVafrRoyiu6iLNYf+ZFWI8HSs+osiOx
bXRNDq7fzr7UWark8u0MFPtmdmFZhZTqVqkkO42Ew+eEdycNslSjSdbe2eyHZilhTFb+56b9ZVvY
jPuQhxU0kEB+S9PwOPpEF5of6Pe+/lJHBvAGlmz+bpwXR0RhNlI/TwoEJhgINlWQMBPB2Mi3pH4F
qHdi5DIUragn4oetHNEQSZWv8cvkKmVb75cu/T9ARz2kSHU9Ytrn12n1/rDKd4wpTf6WcMvo6Wts
pXu2XBPG+SqlYGtf06oLiffSittyhPzfRWVjWYfBlvx5spBHBrQS97hyr7fdLR2t9OeAS2rw8nsR
6+3MRSS2j09pJw6Ycov+mQofBL0kPwJcf/YdecFK/nOQJOCzdHpiilLzsk+QogfNWk37Lleczf4u
Wsrq87u9CwEem1AJ73YDINfUD8ntkm8UrBZjUPzc205Vht569g/vQx8dXWRGgMapCHNFs11MlDxs
NPe09VAK6Wy6F5Qr4J1DVKsjIStCwmu49PyUEJvJTE0dmkWgE5I+siMpkPky+O+MplwfrDY7e2wN
GZVfa9sN37vWWbX8Kkv5jPLNCbKK/Lyq1jn9ibL00y5wS9ltFoIp/vFSRI832wtv87sic1scftf8
LVeKVK1w4cnZwj60BsfyUUza8gzrG3jT4ygGCC2Tc5k/GAPa5VO7fojNYFE5Y+5mCizk2A9Qtc0I
0hhw4dV0pbpFu51I9gbSjaBnnmLfyrD0ws/swkDj/5ziYIj0FwRn3DaL72a5gKaG2GVPhDjRcBS+
gjV84siAacmUGk70qMVROXHNmt9SeNTeBhuLvMgGtOUquYvhIk6kc/iN2tQsaR9nzqwOQUkp0y75
T0JJ9AicDVo1Dy2kJ6vPxZtl/FU+ofBgrtXvPJB8lQligGNbtOCWbZsJz1D1JzwgGFAzLkzfHsko
qrX/nyPaWaBos6V+5iwQNsPT+ura8M95n85vaokCl2Ntx86ftmdgOzGTMyEAF5qo5P4vgDS2EEy5
O5GXMLdwLUR2y4sSa/jqb32Ijq7Aeh1ha+KPj3DwuFz+GH1Yq5gGIzC/JdWNVdqYdmH8rx9luKT/
4cJm9vIPNW1FWJ3hXJ0jCHDKcHV/3m+rnfd8oHE6Tp8qJRUcH5u6cDziqc75Lz/h1NJIrMtUiPya
tyd++A4JHwkMYznEwclj5P3lqVIh+sT/QhCISr3NDbpaQnwye5eBd/lFgzJDK6c6VuCK+G6JJkwx
RzJIzpIgr7LixtPqTPXYuxZNhmmCmKJQIKqOQt8o3b0t9EB6jRUXh221XcC9gcKQlhTPOmmIi5hO
VvgU0NfEJVL6AS5xbm5+Epz16h+VALCsLow6VXLSU73Yj8cU3nmdIJxkt9qCgSxwkWYhYwKeevTs
5/upsL1SOCQNmqDCJct0XdV1HS8KQCtfcjovjnw4BXGx6tL5UnmJRfhj8Z9gOBlPFM77KX/h9vXl
24nXDX8NfgKzpx/7F7Crw9lZwVouuIiG8jDRaCA0dqAcV+gKqpdp/t9tPuyZceTo0cmotnSPdYDd
YN55DqlceEMNQmduzrJl3n5aQPDkg1Q2ICaLUcvwpwNFvc3TAQQUwjRZNwo1eU3n2LtdPHBgl2QD
U6zwTocqQD5zuvygv34kfbYwALNezgPomZWdpssi5fKeF5Rzb2BAyYDIqSodjwaU/LcEIoIyU1IZ
m+2XpZwRR2Qpe7vPg0WmZqutdmK4d5dqAbRi94wV8LYVpX4PWSFzfd0q3G+IwqNBtQG5qZDxGB62
qruzou6j9sBQmnk0Sn5DM4B6XwC16l/l3wlDE2VV1vnOVet7XoNOBSYOp66gTX+0tkvb6e2hmeJz
NzodY45dwcZmgCVmSE45Sv3JLlRKLhlMH9pay2Hue/1rVp9pGPB8wTcyrn8MDEM1zUM9L5aPeE6l
zm8PC8rP6wD0m0cLXBXiaCXGxL11xrQbTduz33ucLElG58L923WpT2e/3XSeLxdDjMY1r8NW2OsO
y6HFsUoi8KSttY86BNHVM2cLrTZP0NoT5Zq6xVx5KSVcZeTPP6KfrJQzHRbyQ2iT2Ud0/EPRmlGy
xuotUNytTYG0u+0AANsp0eSjAJFpXWnRbaT8+v/ZPnOHlpkTjaeUZeDlWcQWusJudwQAH+hL6Lmu
KLdSeopLbHf5iOy7FHUsJTt+AUkUvBMnmcq5PZtljPJFdQKBbuZppp5MjEqO5p0HNIWtIdbfJpy5
qJIg81qH7t830gvxr7FTCnqZYmDQcc9O166KAaI1cMUVaaaud8G87yOlKExGf2VXKgh98qVjtgiK
ZCcZIv9+Y+qX+M1oqsZsLzn8VlMMZvm6G+pKZ/an271xboIuwmq3TjoLGSx2+IgQOuTqitqRMWAY
e3jrRWrGE1zua2XeTfS0L2QTjyIumsFPxPv/ZAc0Lic2r4lh3kmFLsOAjxdtrC0HzTg/kDUBO2to
ExUcJZy7OlFkraRM+NyStPqE0/iYJorenqhJpPnnuiFEV+eP/Ip/xUFN0Ys36jlhLG5zz76zRe+P
7jUKr9qzKae4dK/Cy8P0MKe8WdGElGPds9D8KxGpPzGLnMOG1w4Jm5TphwPlt9ghDYsRnkVdBlAR
agIwGUTFcD5sQIgwnfWnHw/ss7epkkIb28KkkyfCk/uyO+LJkt4pBZv25LUblrbjnArkgynvHSQ5
HLeMUlxB5qxtBBUqSt4BgKP5FRLFwbUD+DmVUeCHsTni3/UIYATLUqnWqUH3JfHY39BndatyuRhx
9DrUE5ST9cVlwYEYdOILLbKwjyt266r/xckcHFYipWCoLbKQmkcj2ycnCN2e54jw+NCkBQDEtasM
8rl7XkFBRjbIMlEffxF3wucg0lTVu+tMrvsoLkvXVImptUTSyX0Q/i4fr1flGkxjzTSlPIz5aRwQ
6kIBuuRrAuXlIU5/qCMZ9rsHFA/Cp+G0mrt/4602AMd7M+3mLZdmZuFN6IZw4HBsjAF+7UAgQIcs
eYxZE1Gf63Kzur7ZcrUEFajh1WrCENHNv4gKegWSbDrlTDXZcMKr5gMeBtK7v0TVx2U+zl9b2QYv
j7JL7e2prPTBNBH9kNEHJ41qzclj7q7Xe2DOUKcP5kaTxTi4BSWdNA6wfRDRWRDklD6Yd4X6K3xn
16K/rWVqm5yUjp2dI3gfOSPVJb7iwnSJItTgPbQg54fMSu0gzrEQ+Wyq0tuf5bAQiqIhpnODZiBa
fEsuG7HqJa7wvgXLltn8DtS6C6fQeCaZzMInxZZfPrrcRg7S0uwyBAyTyEG+xk9i7eqohLRrEmfx
t3HOpKZpHtamBvlxFI3hzvYS5oVlBzB294UH3fLitODqR84khCFUPWgahOpLC4L28dxDSK4tBlo1
5a6DZtzjGm6Sq7K1z4lbcZ8KwvNoquq/8Vm/FnN/nGgKkhc831Opex5I+IIY27mGNlYp+9pKpY2N
S08Q/hE6SFZQkDJxAZh5iL/SlawNg7M+QKiKBYAMebhUmgphfM6CLALn0WEchBBsDCB0bWAmp2Wp
a4w5VFoIWDVKQPjckjOfB6acI7nCtLt4LQx7oJuEltDzBw4jLYzllV6NvOURTQoIF9m529hGr/ac
7t/lM7CubQkXbMppV9463DzXyLDNw09NpQtWc8fo4IFB+mcR4QizEinpu9zlEZaGIG6QkrZb3UQX
rmolkhS4hkxgDUruBlbtmdeV38T1WxHh4xZEDZiPW6hlRPtnF756o+NFUPMR/ahJzIqS6WqJnxBD
DcUfQJM4cs54yxMAtHN5zTPWvbutApJiZLUhvR5u4Rv/M16+3dPkC4QPA8JDPf0aP1Z2UV1D70G/
VdZmzUP6TSRo7xOfXE9UTIBkiCfjfhfw1rhZLXAC6QwOtmWI17LTe7GEr7DE+y15VMD+24uI5J6H
FfVRi+IManysYdY2cm2Ugy3lL0xWadGkpLhEfw2FQVIYe9cLMaz3jhEXx1KIeSclFoxmoi4MmKj1
Rr54Pib4TC+eEQNLHUdGlzOsK3ws/0N3XwWMX71u9oRl7fClakSCWrQP/H15xFfFGFZ0Xygno4CO
qLzaGCdzDHsOiSRXBirfDe2GXIs2lYzNtt7LAp91FB/SAKckwq8PCI5rtjO4p2p192SwhqpZXArd
2VlA4O8mSBn/8I778bpu28tvfuE2yKnUTC+KT1Tu7kpSJDnPm1QpKcA9CPgtzQbLqRXyMiMUChL1
M1LnUo7BwvtE7eL4MRYzcE91L4uDjm+ZaxiqRX2y+LgglcjO7yEIW/VDNEXmvTCTodw1B9LWpgDk
hjoO+LfmyfRv5mSMH218qpFvW5+IUnzqoZy82qjF90Vhc2BAIHSkGcfNMhOC7JOTnPCvyakod7rj
hgCL8jeVmPxRS5ZMaSSOTwDY6jpmyr4cLoYRXzJdb3zuF56r+bTCnEEoPJJ8VSzCwMrSwrIzxX1A
gsMbKzgTIm2UzSHseP8WZKXiOTJeIIQf0LYzAlQiOzfMzHuxlA1uYb2WeeZsLSW0csFTOqkN3jhc
bQsAeL0HESXVgi/O7qTVC0Oe/BbWSzbaFO+dTwEKSlilFIqpn4iepS3VJye8pbzwwlokE/vft2DO
u4bFNQYiYFo12FuouEP1Wj7NhEiem6C9q0oXSX8d3cUkkGefBTuq3wtcq9muwokDoIhLaZDkegiT
G3WkAKwnVOxpBEI+RGEfUbmHEn6m9YtdmdPPPuq7fncY/c7Hk9vHKrD60+BylbjUiKKQpWN9ZU7Z
6UGg904Vc0taNZ6jjHuLIkm34h6gsgSnpEokoiZwKdcoWQ4kqhtS705TCujTi492Y8wXmzlf7qEI
Q2fkXBpViwZni0qEWz5i/EXKUoF3ExyaypGbTKjRvpNNTPxmnLTr3z2HW9+Xl1NcPVfVIjn6/Z/z
ga6S8HtvV2VQyX663DWsNPADy2jIx8Jqno5TFkrtNFCIitx5v4uVU7Zm48E8u0w3GOjqDj8YOv9j
dxB8Gx2kOw6V8oxHP9QRMXfGZQSvebZSSo9srQHSrd6ehnCSPxn0XyOXR6rsfVrJrGQUDGvR9AlW
5PdH6B/pVUkRjVLRNQl5O2tsJuJLohMHxchBKQX4xYxwkbjo1Evt72B40s6z5G7xNSyZ8lGk//6Z
gkIfZ984G/nBums6q2+WmFMOhkGko2cEh5GplLm1mt6UkoUw0C1UHESNt1ESqGSzCUoE00iHk9xO
CxMQATezSUzuYudig2S5feyfwQmr3XJqRA6GaAhmYtUL4xizQMnFO+Nba+IIBWjqfRvh+XgLWNjq
diKOIJGr6q8IlXRpsEPT6fhb3FOG6QcYyG68oDMNw72uNGXZUANBCS9HxB6a9s5iDkAWK4j7rKHg
ibmmq0xwSBWaE2omwVHJHKqg+bhxObgqMshFjQd1nQc0xIG1WdXbqtoRLahlmm4+B+dNfqdhnFtl
CVUL663CJtTeI8JyuzG23tOPA0YBVeqMKhDVAlv1zO4/4cBUeB8TTwRytiJIrbRfVz4/uEkcu7y1
f6Y1AC7gaktBDiJkxIo2RN8Ev5aYyQXc69PEcs18h2+aD0CrYGnv1lWbcHcS5La8su0K04VXB2fx
91Ia44WPMwRVeD9Bxpq6Y4Y8npp+5HwjZ29FnaFKVXMcjoJ4IaOnaEjsBB6BzFaIPR/WCncv1AMc
ov8L3VphmYhpSt7K65+vAM+5e6HzEeWZIunB5fwxT3Xxbl6m/Yros+yNI+MaadieMLCk+s+gnkFB
jImf/YtLusyzDLIcerW/+m55YdJfst0HiIz/MSOxsjKwT/x/3Y5QX3+9dzuEDdyVPA95N5D2MlJN
TP8fZbVqhpb9Pw/pfGH3wE7NOETjA80HafORGxknkXmnBmb7VDXwtxvPADNhDUXtb6JtUePT+csP
ooBoZVdTl0Is8KlBxw8pZeqLBLEsqkqNBJNJX+E6ap0D97rEqvZTTlMoMn7U3PWE2NnKI5qNb1o+
7u8wgkJJbFbPUpwjxMor3+RAVatj2zqllJ2vDGVhQEIfCZuOWJS2vGmXk7vn0r7CEEqlK4v6enkd
DpU8PgkR7HnDU1ui0oP3QlNX7Ki0YR0NnbB/SNZ1ryBanhxoywb7R05DQWCAw5d8GDyzF644Pr6M
uvvPFYVkLg33WXwuZSOOe+uldOgJxi35p9oAODPqq26hswCjF/Q+QX36Z4HBePr4fS48VqsHiwXu
6Z/wTj+sawVMGjptPJ11kThfhLoseNP+2MXQk0m8nzNYN7hGLpKghBENWNWzuMDVcn1Jp35KqMcK
RUR9plX+TpLQKRD72hGC1HNvs6KMYxi7UVz9hxBvsA9xrKsKYmQr56oXWpLxn1IBWkud3eT9MaXX
IFS8KLsXvE6MuKYdtX9HuSK/v6+7inhC3vMco48tRzNe1wM1MkbsE/tJKlbIqY5Ud8cAQov3OEFs
VWWAHLbtyZx/EcK9mWWceuWOp2uO90UArrT6cCEcNylvv+Rp6lenkRcnI5VRAUbZDcoJyMmY96pN
yl6lGVMbFU3vhQfWbfezZPRvzxZpDYBv0mRiplgmOB15PPjXny3AHx4JiVDVDixnoD2sOymJDRi1
TR0crn3L6EfNNrI8GYrdSXX+VFpFkcq6TM6p6ot0LpBMxnGgkd+u3fy4S1mmH0YlVemvH72ZlfZZ
HAFwDI5Sgn3KrpJLVnn30Qz6SAmNHXtJVvYC7Gi7SbkWBnjZLsqPG3G3xZCJxoCMj8ghjVQSOAyW
2v8NVn9l2C/EWNvZYYpkngpOwclA3J/cLLNDs0xDx4ic9U+ZS7BwBRTXEbL56Vcqrcq5R5o72oJE
RT8M0E5bbmMMckMmjRhDXKzMjphMUVkx+45Y4fo/0S1UjngITnyzdH8lI68Bnj7jyNAssun3SYLv
17PhwqT/zOgWYUobOQqFM+ED1n5MzEKVd5XDfmjXVulC62IhHM0zPZd+g9EVHNQrt8o4iOVec9Tg
THaIIpich2vWD8TfhtAtfa3H5SSzfW44fHTZvLshxFzMJ5P2f8snkMouVX9Ksk6RFGGibUa14xI6
FGmFUT9/4tpe20s/hZXy+2Lh08SWoepvCh8MDadlYnWCe/ZBMAH8on/8yxD6f5vxdJ9dIHEt11rC
I9GA+AYb7QSxVC/M4ZYuGIv/w/TVaN9VWf1TVN1lYYDiovTDVNDWaUKwu5O5Kd6hhjpWDvT46aUo
kHaGYEhgA7s9n5p0bvRdxq4SVYdL74K3Fklv9zji4sdooyi+KnK/PDPWKo6qVAZDihF+iWZqu4dr
pXLjWd9xyWss8s8NNhuRQkCZUSnnt2gTuxoUIaDMx+8KJbtHw3H6mtOrJe+bclm1vw99v29X98TC
kCR8y1BaLgtRazO9eA+SyMdlP/DSUTOv4K5i4RQSPx73ed/6vQiduD2JgCzv6jrShoDDvS6MSgho
8KFCUMXSD3jkqsWG00pwFMppXXed9hIF5bWyZNxSoSh7F0t/iiW5Dm8ek25TnLNZqTPsbBh1ICNL
0SEuobwmvecfW3NJo6ulkdUaucT7zaeVgSQB+O+y7gF6QwI2NtIAMK7YieniW/pmtUwHNakqB4Dz
yjxeEY/e+o3ntvnnCqhk5+wUfpTHWEmnmhp4b/DkC4kB1iT6gqUtWCMPh3qhaq7NwidbpdTmlR+g
//fbkDSgS+x5vFjanNBGerDmYVo6w78pk3TRvO5DLTXy+DfZxQ43KkppiB2qeB8MgQTO5MID5EfH
aJb4TmqeObA48GZAIEcrfZFV7yepscwoCcRmOm1mr/TfdSVs4dBcDXZLS6KOiY1oCl6JQiVCPk7N
GPFucB9HRCY3VdJGRC+oDECKGJbQULf0meeRb2fM/GVEw7U16Hh2JK2iIJemkLZ5X3+SXwtDMr4t
UqDAl6RXB2+GiSeEs4Qm1JOJK3CX8KCuJo0DosUg2FsE/jCXVfAys4ZtSWo4WCMSEXRmRQ65WXNF
pVc0GRixUVDwSytlTQYRMXGt4ziMGDMcn4UMRDoVFdopLqFZk93noiDF2rJBj9iISZUzl7WXYPKO
SQG3twwcVfrwK+C2BKb0BkneLAfPwd/95JHt0aV/6b6Hb7oI+1EyXvdumpUOgxpb0YvPmaY/OtEt
pccXmfXLxKk22lTswzy64fUfwYOYgGvu+0Gfcre8XiOFj1+vXWKzdtdtJ/s/MGuk8xLc19vBZsGl
gyar0eGLGpMk0oOLyxpSvtlmveMWMGA5kQynqRWnP0rAtc11fJFC1sn0wS8d2de4EdivpQisDnsb
N07aRCIgCE6VkDXHTPTH/gHqmcMV41dVc3sL0ZZuFkZluvoFHZ9JIZYNOAFsGTmZG4Djg0Fuzuh4
R2ahIQW7cSbWqOUI1Wk2qM3GZ6hPqqxtGEq0fh/ItUSjkg0r2Azs3CIy1fztKYHOPlBCvQBmYomK
eR/qwifqA/btwFusQHyy/XHvlQeA/o9Xb0Cb7XYEUgR9NWzCXyZ4XU1pmOGDeloRai4Ws87Wb9BW
Vt3kOk2tEZWMLk4rDqBFEZYqmIYnWFl/0OdwT6F5SxTOf3x9YAKGcKj2qsDqd1NfuqBHq/pnJuN7
XrCXXvFqUumWpswLjWJhjdxIfevaDJQQgPidzJz7DEm9N9ZaSzVu18Hjs2gHXwCZIuaxeHQkqkvJ
pg+2L9wEqDI/wW+QeoVgW57w1tQMJn38Z3VT1CR2SnifY2Z0igQhBYmxXfRSCZW436YFh8K3eLFe
y0QYimiHJA4tgdjXaC5bdzdoujWr2elJ8WNVOmNako0BwIxFl2WDXQzmtXf7zVRRbYU3vogeqYHU
bQ1w8UhwKDy1XXX1ot9ByRPE29xi9bZ4Mg7dUGuY/FEFlUluD+L4dT+Wh3oV0QPwCh7AJbcDRzq7
uFj7CGembRSARy30sH3dX1AoRyY6xaI0ba1DqVsxEhg/smOJsuVdVIppCgn1A1FmClgGrCANaVlH
hhicXOC4jhBjomQ8ZzAWlbdnr8x4q+soqkj7hf/FPDbwK1rjxTOz3cfTcWWkG99qenaKgPfQ/K6u
+Z0kE5LPn7bk0xWSa8pJkAjduqHykCLJB/qDRJYMGRMmnLL19VPibcGsaEZY1mJ1pTbrzZL5B3Mg
+QeW9c/SwPT3Eoi2xWq3TGZUCKpCNKTMEnC5cWlJXukSi51ez3HWvW3lhwABKVOCL/6VYdnitvJn
uLXHIP7JxBlOjgXAVaEk9hGMJmEhxPnZtNyS+bh4QlEywSvU7k9jgcuGcDMt2zBxKqnI/JWals/v
9mH/JSEdGKfQ90EeQTE06YPPcB5YmtZ/8ttPbytRlKDyHH8m317Y1XUQSMVNDsKN6atIqQDOi9uk
nuDeXbcQnu0l1xn1hmeH87FJ2WtA3y/Jw7aDjy8tBKJT/n28YAOODyC5ypTMviBtJKv8vGce9xBk
8Pnbd8zXvDsBJIkssKcAcw7clo/RMfTCf+Ht6ufJI2qCeFD7ZgQ4nffr5u+sKiDjGLLR0sKUQSPN
qA3YS+6Nkz0BtcAjBzjfn4744ailvAN9pmm22wCTbJvGhARcb9dgjOCmTmd4s3PDRGAi17jCmOvP
lg6tJEx44DSMoKcMLiyvdYQ2gNMw/+5nGcjLlXg73edxszsmwq3suV7i7jEzV1+k29Ml0JBvQka4
f6GAJxIl6rXSEJCjuFb1bzG67Z5QMUmZ9gHn29Ig2Rf0ht2GXC3Ne3QtJrPA19kPK+2mkK0u/tem
USnzeX/x5WqYQnD5YuCW0Jg6OTnx0WXvHujw2Am61ldhvo05VLijl8ouxR3gp7IISKH25aDEcMUg
chlY3MH2sHIT/jU6iTsm2h/5g8yBZQ9YkGgBLMgV+ALe/0n89Jklvcx+oT+3E0SYzjsTvbX8gfNO
x6EoG6U/Jne/cvXlquLg+hnTIQRcuwvuFZVDQlll1qtqWC9WezobTops3fX+tOk6ZvIvSsvlQUV1
ZWcQucf+Dz5BcWyYZgU0PxIBvH7NaIh3+TVx0+K1PPQdNTk4PBIAn4SSSzwIbt7TlLAFl8WAPD8U
d/Q7dNbBST+Yk4MrKSblgkkKxrD+dqUi0muJXl/qqd5uRBjhbUjsKm7hXACvxh22WXSyMDX7JQ6t
QzTgBA92sPdLEyyuevhfPXTZDVPdOWG37Rnuw1bsm3cQittAExlnCKlXElhvqnqEIE8hcO1hTCaR
bp/NL1Hv8SkvOjyLdwyxlP8NTzHvvMuIVpjMQR7IObEL+9FnLfcCY2DTwEatR9rjmI1lahQXbPaD
ZJq3sQkNGv83Zl7yiEvSRI6fX/Hh7LJ21270C9R7zsKNhPu91f8rVscDPJ+9Lh3ohcu16VF9g+r/
DIR4DD5/JFxspVMxcWixd8WovGnDby5pMj5A0a+fZkP0jkaI9iECZZwavUxFSAbWN2Uuyz4hP7Si
p8NUYsmw2zBCwcC0f7Jlpm+WA4dCkj0JbiPR0n/PL0Se4A0TiYZ1nSovxHohXUEOgpZF4jhKA3Ir
/GDEii6N4HWoCvrltv+VqPZ0strY1VqItTxGhppxahWYePhs+PuSCpAFvtsTWQoEhqXIxcVsNDnr
tsApJM1/y8gXbPH4i4YQ52JYcmz9gfR9+m0XPq9g/9YHKIf4oo1rfW9KEyTILLWo1obSRIpwP0sX
4/219khzVP3OmXI1JURzXiwvyW2z17qiw+m80qOQzVPcoZmodwd5+2nhIoaOImkbIKaoFG+eQcmo
/9xJvkzpwpgPYt3zx4djxbzYXnw0Jk5vv2vyDpe9MjqsW9VwgWBRrvJ7q8rGhupvBOLs+4xZOxZb
W1GLalTZyY8ljLkWK/r2BxVE9tBdpVuHiluBgFy3SptIww1RFougHFGXxwPQNyxUhsdwP5Z8vbED
YAWrteP2RrJ1UbJpTMV1ADvhI0yXGEfSigcs8TbCmVmSxF5lgYBCTXwx1ZlONDGxUKoRTP3/WqFZ
yVnRazfxjJkEeuF2k1Kiyckxmw1F98eJmne51+8saDNOHpOCljVAgr1Wn5lUJVzZ8Ss/lWS08QKt
S8HGrO5mJVT+PMBd9ruGyXtDA6J2BDX2Cwh2A0IsLBvrigFKfU33F9P3iICs+tCAStaAkVkXMY9d
0YYPGJj0qrk2y3N8KEUU4wePpDPa6RGlUhRejqRidlq2/w3X3b48K6VYb8pf6n/Y1b+WIFeVAj7o
Ru3fWdOgBgFa3SuVNAqW7jBWrYNxhqT37WqKiiJD0PQPecTU7mtshtVenPx6gGEhUQqg+HOWOMcq
WCkjWILtI+eUBvxVvRX01Vrot1x7EtmYpvKlo0ohZTayhOCMFrJfGsaxvkBSr17H+DpjDQUurqRl
Q7pg4pLn0Zn/uCIR4CwllRBXf+6RDbFKeGq2XGTXknzZ/luUicSoKxNyBw449eGyfMN/FgCvhAM6
AYWtIQBPDg/TYiht82we8ZeF1whGk9zaAddP7lMDMaLD+0TzUGcJh4FxP2D5Yax2WrwkeURGGpuA
jkkR7J3Oibkk7DwWD+CTxk67FgosKBWRvSXc0I4/5IRJDGXf4c5IpODjjLbiAMLaHXA23r+Fy4yI
3mlVjTy158Lm3xz+lddWOzZzIt70/AwFByu7dutkYn/j2dfkluz5XESXstEaKbDxjuEh3Ggy4DQg
wXeQi1zndh6DSSVd07dwLu9Myj/LpqPlcuM7iYt2y+w+Mq1jeOuU3OUn6eu4bab857O81jIviSSh
Ng8xhYGn3S2VR+BJmDhhCTyj6OVhTHyWHAKDprPE03pPm/kG9UoN+DnRMdn7o9/j46v8duWmbQsh
QJB7A6wGpO097kO3/+aA+wAowQuS/m1kelBl6JaAQQlDZ0z+s9cy8DfpPZMYZtjLxh1KyCM/kVo7
sGBDKOUd/QbDOLNb1tbJ/sWkwH2nTzru6LXSjrf3bAIpDluzBcsNQ2/hZUCyTHcr2uXxUhxKJ0pU
48x86KZodkett9VEyM/zmAPhWEJRyNvx2d5f2N2grjPEDxAU0BIOR6SIurvHHNHlv2NSY6/k6qfa
PwTMy3dShryudHMTkLIV9/zz4rjAgY5hsapN7NxpFmdDWYdZ5d8AROjAopEvsU2OIRTebhNmbfoW
iUZZlSx0I+sNS/i94uW/dNygnu90IkhTselKGh099dtfDGxeNRUuBwTy4Bx8tp6/KP06OqCA5Amj
1JOE/8vAl1S1bhO46UR4TIuZYZ6rX4cuPC8QVHSLjIznY3Khv0+x5rBs43KYNwJSKTNu/zXj0/Ag
mPqkDO3z8t8Inw0O9vv1wXb8usnGpQ2JY4qelAsyw0hGeyWZxCitRTx8PDs2ReW4DTbxwYxg5Cxd
oWbbY/WALSLlgPft5qwh+Xnt0VGyQLeVncIAtW5NkunTtYAPbRIMP827FQbq5ErM+ALUzxIRfsmr
l16M2dLPg5ZNremobCUuyHp6EbQPwGjpDpBrdiXLNGjfaeot9NrxRbpW2errr3C7YZrEmFW9E53R
CfcQquUgbsp/Q0zMn0xt0UUaovBGdm4oti7c4qpNIMREiwszTfbT+jBvIWurTITB0aSrDVe2S7yG
K+IqKzlZfgYHvjjGPSJk1FOAROvn+VioHWooDJNHZnYgop3uRwGIQG8o4A0MyDIBFPbOe9RZeIcu
+2aHb1nP1uq9S9SOkdItYSeu8t+sTm82XK9oeonyTmhsIQGQsAaXYBkEqu3gP4G97P8vb7/jY+Ly
Dw2y1Kmd2GKy3cJdA0hpu+xxgzowNj+6lZ/j3eog6pn0cx2Ylj3eRPZ03rwiKX26ulfQmKXu4hEm
KJR+sHlKbxCoOvF9FwvapIsb+37N/MuJmAm//oDPZBx1Gmx01cA1MuoZfvfEK4ATkWiOfWrTOet8
OA6uCLkd0x17G5FZuP2OEI/LYeqwd1uBGGMAKo1vpSTGYz3parECpqXYvfOkLrHoqXmaHEEoLnvC
/SmG1nQXIKq0LXWXXV69yoYc/o0KdTleY2Blpm+HXM6xuT6iEZQoHMT1yIaF8LKUqXUODQ6+yVyl
L9EXDdEDLVYOGzcGNfE3pm9wpoJ8Z5ohbwRr6kNFLy6bdhx+/hyAX22M9r+taDQhCADQpQh3rwoG
/F3T3lMN0/S3+hA6cYzGn7oxsP8kI4p6GF6UrSjatd7iUZtoh/nqalQg+DLdWZ2JXbC2KQpsok6I
y8j9wxsKMbPURwVQR4qSDXfUCM531hhjIQExtxi6bOcEOEIYMZNxxLcezRs6djFAYgrw57WlKAFn
E8HOICFM/GY05t1oTs8soi6uofnjvECXUzffk/z11uFFH6oq0HyKzzY+h2U9s5oywMSpg7ew+nmX
ECiegOG5dRlxhWw6usXS9YWgfrdkPrOz9lMCnUf9L8AOA3sou9sFqG3Dl2Egf3FR0RsVNKmVpZ4g
v7mz8arxEZ/bMHICzAwcrcFCNXKCYIQViQK3ff9szp5BorCKntKab0yJtDHEucMD93+nopmymXmh
ZoTL/UtIvPQMek2nOJhdoSL/Qow/dZ71v6jkwtmaNLjoQ8gRllsPh0ZaEWR9jruh72ilaaqMMyZa
SUBK439k9lI8CUlxGTEPy7dh0QvVtKuARO1FdLVeKX4a1fk8/LVVPRD3+IaqyTg5N/aQWQ8/zmfp
N6gRRD3cAu8PdwJDoKYQ7CbK/OBcagDAX/ZZiqjVXsF1PPHVJBGX82+47v+I9ssECcqMKO9hlaTc
lciRCHugrfjIknrayfVFUc/M8tD3bYhd/wzRZtA9JvI0Q2vm4o0tHBklyc5Xeawl1fHYlJlq/LVo
rWnzIUtsugUfG+B/H+Lf+yleQI3DXdk1alqCFaQpurmdo52Ol6fQrRbhDiStZDHj2LBrBDs26KeN
1F+7hY4GyexqJMKLB8mlGU9MevbJyM5SUjAtwI10DByLkjdd3kTalNhHwaii166CBfT7K6ljIpDn
N9vbbrPDlcws0Ppki9Zoc8gD61scdydex4L3wUfG1zfoslMvCZHboacUWKszZnbS7/bnMRDSKHhi
TPrwMWmwHFCfSl7kcJLBKQpSCDvP+uRwBGjDINv7tOuXLYAnN1lKYh+Cx4EqfaDyPotqywU5TnxM
nvrL2L0k6kbuMjF0ZWcRuFzBUsgoIi5gUwhQBIzWcc1dOUrkATwOh2LKK2r0c1R2N4m5cyowCgp3
5OQvJP4cJyB7mTpWBb0dimyi56Uzmw5q7de4QYrFzThTFnTXFVPj7CO/x5pHJbWX1InYVEma10Ps
j+x2U6K3NQdS+0uRfZp9YQpFsv64qz/C6Kmn7d3gKifvBi9cITm3mWRnZFjnrJk4qA5h+RVxmHGl
RqjPpWPICsQKrFwrSwV+IKNxRnMfe7la81fR4ijfU9P64VrM2VQ+VKwHhYfDgnCLStFgSpwWxAqd
0usAsVVzbMu9jjRqhrzw3CWf7FOb+hsWN7JMbg4fnYiHeW5Jmv0Sew+a7uVglNElARk1T+vTnZtl
MuFEqIqzrqSNZmUKmTkfDYF+bhE7UqMh9CVshYhz+l1yWAI0GzEqiRjTG/uacOrB4S9FnR2p8J6a
F36tDGhRHtopU4inERgQr06ByqhTFvkJJyml4W3FvjkpvBnQ4iIcCF0Yly+M8j0gSw5azGXAu/MT
W4UHfhEx9QW77yo/pWdO0GhKFOalJuEPHjE2ZTwLnRnSV+s9MfhgvNKeLRk/rYeciAvjibCRB09R
0PE8AEoCowk+3lonJ2UQCtj6Z6Putd6IFBf8K5LaIxZzvt2FWa1UMnRhK6XUc+NwxYY31XyVLrJN
YvGEU/bG/n4V0uPYHbD3wk2BcO9cQhw5VsX5muDKhi+lrIKZvX2neqYqID0qtKGMgVDaC6y34faW
Lf/41C5cYxInp0JYH5b+X5cUPpylvg9gwecSBOz/HVxW6QtNioKBF2e89c9QgOeAOl2ALcICU0ZS
s3gdYMfQsduPcpHtJK6EbhiPOCgNy2iJdKpPsY8jUSPM4Qf3juQx1NahDyesLQs/CclPciaNwtg4
1FxLtt5fpuvcxv/Hu8Tn9BeqMOxESB5P77rSOV4kJdTVNh89ySpCvQUZwJq4iNXFt76KkvCxKBSv
cEWCZ3UgNjF/46L5ioUG+PP/4/vVrdnXXbAIi9CYIBTbZL4NSvP3WPUMeYwGOSve+U0DOFgNcxOo
tthaX4ygxuAGM4NIwwZn1nOIx9JEQ7AUernjXkkA0u3bjbxFo5iEe0d758wi0sfX7m/4StK/pvUK
eFk+nbg8OjcEUsiZfPDxrwNMAFLvzljqYZV7jKlkxLtIqe3zASmT5ZOOB+wzRxFIFWs6gefwI0Br
VYu8F/RteccfPlI2d/PY6TrwcRTF7jwTNm78MyXKHUd6JOUmnvhiOMX85W2yzSvxEjEZs39Jx1pX
c6zIsfhI3D8rRR6/1BAf9V6J8gT1UMekcbImCN5d0ZwhB2F8Fm1cwGmD8+ARlFcffhC/5RVjxKmZ
nUAfB3/9aP5Iz8ZUIJEylbCb0WOFXpb0QwxLnaah6JG9kgYxCcQ+R/zrtXb7AKxnCygrzhlCsGmG
mDpJuLTs3X5UqpaIqjj3Xgu0PlrOzHcI+R6makPYxbmf6mNQpJsyaYyaQKGf6TyYb0e4IvjkCs4i
eF+tGzSVElSykBxHReFaXnPSr2UF+pY2JKpZjzXCTbXzfSC2sG89mqgsIp2aqfiYYlBJ8cFETGK4
p+xS82PGtVrFuzjjvr1SsTBGqZQdXihS/OeFjIAfoxyTAjVKM1u2x3r50ZI1fYUJwQzKvwbXXlMb
B752Mn404zWHThBUSx4fKxtCPAoZBvbMbXMY4+Tr1ezhegDv/v4dMKI8z2gdpfFvtSlVknHV3sNk
1RGry0KzsbHaiEeGXvkjnOcf5jLjnKWc2aPtPUdfaHOkHn+wrqoVGaHZIZSN1SxnKQ/w1kEL/oJU
pD6GHxspPMjtu4mLlgPK5s+J1PoNFGK1aL+sOI8Gdq7uzFUOIqJvqFq8q+JlhOJUbg6kMwpvL9fE
gD2Emqe+SFL+D415odY4EZibseNhJwoiWkKsfXnZ2Va1PrnappiQGDk/QJ1Dz5HRQTpB2UigQG++
+wC06xO86KFwzUhVsFjic9JY7AH2tWiGUTLVGo6CKWYkI4G+cBMYScRDWeeT6xpSJVIkOlCVwQp7
qAr182osB18HhE579+gQCL+cFqJLT2fTLJTm1JkbiftB4267yQ6EBfF1Bcy2IBbaYXv9g79t7UiQ
C5BNRAynHYbDPJ8oFEINa0TtzTIxOTo8uWAWylAd54ldUl7ZlTt+audw2PmFYmwRYU7oHJuyPiYU
5c97k6mCiy/fPbXbJVu0gX+9gxbB1gqSKgkT5Yjfz6rPZm3Z/w1KPGQH8dLNS0MAWNk01rMLtE7y
XsG0xbEcPu5Dm9c7YD9W2r/rY+JyRu70kKxxdr0e7gGp+eDvLrpm/HYC/n/St91Nrlydz0fjSlCm
wVHvKrA1OPfAV4nNqcqyxW86a+KSbvqzh9tY1iF3RAWpD2KeYBWwEQ2uUTPVEjxP8DNF0DJv4rmn
gz2T1LvZhuhDVcxD30qiMcFD5xGYbvM/WeJ8SRXS7m7gQx70n07JnC+Woxk3auwnJeSoGqdrE5Fj
WsAt9Km+EWFIlHGghu8an8KCGqFWOrXA/VUrXdWS4X5EGHOXFvqOPAhdSDXFcWRNDRMn+ybMAGfh
lrsYKdRSjxmOGJIqdX4ysCvePD64ZHY2ur9e1xChUvyIgxUR2imJ1WhxnEERq6FWk9b4o7YVAAJQ
UqOzJ7OSnN4wzLysn3W/aOZXrTVf/vVgHcvf5ZP2axzlUP0M+mQ6niB03msUh2wMiY6A4lyJUUW2
rYyiZBTDmP6SxTD3ykRz+wuLlOU6UBax31b+h2qoDvO3DoTnZbxqhBmN36sbVm+30QoCNfuHdyp8
dTvUCc6ZCVgVtYPZsZqGTL6J516ZcOfn1nqq2yT4SW8hMoWTVgvQnAeW6ZWxwjEzFbzpstKmPPWj
kKPQZl1pvFobZHAvBeqQAGk1vwTIB/BskVCl/oVPsU1Wm3xUE1VC5rkLQdiBniq0RrfKL12uwREA
jEw63vqvZkQskHQOodWhqBv1nrgYr7QlehKhLl4CJVc7XKP2boWEaQpnxDEN1mh71G+VdaQyPQhe
sqQa1O30kpbM8y715OHBmkOSIewbdu8RzH8SMqyM2/pKXd14g+IslF/Q12h+q4+o7jroWPo5AESb
qgSQGPQWDV2B6/IsKMT857GKV1farECHcKnB8CEqArBH8G8x/Ndmeclb3KYtJ/MZFBEy64iOhOya
hrljB0hXSBNspAKYpDOFip+Wg4qMVmktOJVqSSBMJyE10svfeH5JMrBXloBkoNiC6zny1JTwetdw
+e6TavhdwKuhlYRzcbG2AXWkQWb39d20MCl/wEdjf5OhSn9+RF1jFeEPTMkpND41ZuxPGXHTMY7f
Nums7rgK8hi7zuK6aeij6kNxOAVuA6MMo/fIDOeZag/4OiN3bs3kVe0zrtCrGq21G9HFtilwQ5Ys
u9s0vn5O2WOvv+b05sZecAeWjnKX9JnLPHTYFErnGIrHBp52yD6T51idSmrchfh9LlDrRpd6OKqq
mrrgRmeKSB5C9ihLSlpg2TWIO52C54o9cvFRmqCgc5qEDPTE83T2Q6sH6aUssQOi5ymr9L0QwxgN
LqdqzdAWcyR/VeXLk9mas7FEN37nzeMEABtifDfniCowviiD+TEpdlYwwHSlcTmoyB1pXYSvblpM
wpqlRmIPgvuBiZwA2hYZzXPWipYHKGeTuNi5iK6P486kQJdRaNuvQQUTCebkcVtF6cW9UPm3O5Nj
ueNr1ul8toa+8s3dpH5Uwo9S/8jdRVTRm2jP42ocraWTx6q6WTo4zjXLqcLv9jDsnMG5Ti4nXgID
7Mm7rj9ncgZ7SyMybqatFpIrDV0gP16UFjvoTWMU5oX0T9WrJlLm0U2NQgERaYnh0tAo/5cD9B11
1TR7aVlRCgxmjeAV1M0mwBGSuG3SYolMnOHtasLUAcbjPGpEd7OH7nFq1hJnOtkZ5JA7Usq3Yqv7
4gq2ZyWJH2BItGLf+mKOxqp73JUaFpo7hC0jTsoNURq+vu4YmWIeInjjw6DNiHeAReG5xN/hvZzw
bSM7O5Shr/Kixb9G8FsHknKURb9zbkgbxd4jpXfO+F/tg2e2UmOF4UXkLZrDqNnAAWfUD+E1hWUH
V2uI/AClpi42RnRL/QbjUwHfURUformKPWCeEPexwr1h+O2gBpTwGPtcI5FzeI9ORkbOj07NA9wk
hzogSXK9dq5zCWod3Y0uavSXgR+7mRq4+xsJtUd9cE8EelkEBe5ZRQ6YppMTLrrTq6W7IhQwuiwp
YVvOFV/Ou7RVpyOSFW0oLPX8KFL+ghi/YagFUxOV0bm6rTzPWkh70Y1DLH6R8Agz9fbTd+NpYmuh
/xwZZgz+SoR6CbcGC4ywmZOfHaGQub+X4gogi70d0ZaF65WInQWM6spfsm+4zou81I2a1Aj/d1ZA
X98Gmv/8iw0YlB2j1Vt+ouvs4DGEni2N0BBNslPoHjDq02hZuMi6RphthDpEDSR1BYlOzedGNCab
+N9ZaiaSHBUJUnOiaX7uyt7NgkyBWoKzR19kj1+a9hi8w55ZUDPoId3gKo12RDTybjfNCUm9ZNgx
+7vr14GDIwENMm95o1F4n294u0sKGl4FxB235ue+lKUkiI+PqIROfep5ZAlX9+ULWfoN+nHtPvEu
b4X2YWGFz4OQUOeic/WeU967g3tTPOMHEfP01QCgHe7rh5njCP++t3p+yAv4yJLKzS4v0Z7x8M9C
Z6wPQFTCsEgSgjZGMFpVzinuTB7T2NbTYID1ZZQhxwn5izq1L1ZZJfRXbGUvHh8RH5oIYkLRv1cL
bsrISfAgToZVFWWLGJYWHfM3DuQOnU+jnC91cpCiN8ZsUl5ZJDZyLswJ4ID/B/RDrnQJD27FXbMx
qej4D2h8LRBuipM9HWQHvwdg0PkkmKptm9BcTuK08xXIMSpOXX+BdIlCJakHis9BxCMwLXwSZKhP
G/7J12gqBMlOR/gsb6x+WbC3VIYotk6wCHIPPNcL+qAn63RW7JQQB+nLHAHIbkpiJV40zx2/1ZtY
mMkOWP3XrxYKwLmg6f0C0bD5CojqWYwiCFlnWkghWdSp2Jpz2TrCq8+UMxdRVGZ/9r82g8FZGkwQ
VcAycIWXwmFs/MVDcZvEAbp0aFJiU8Kp4mlmVQa5hKS8E1ZYBsYgV1UJ+EwfSkIJCanLpn4T0/q2
4gCe+pJ8esyheRJTloiIkOu/WGAzJdo/q5Nan/bRT2jz0N4uhsQqJgqA8UTvdpDbhkFiIFpDjSY6
zHl1UjS4TB7kh9ujI4rnB6Fjb+tEOBjacJykuhUJASBtLnXURnvoINF2fCoYSzGuei5Rv50KF9iq
1qJ2zScD+L4gG1xzJjYZ0icuRzWpbANNJn/SD7RAgs2j26b0TRJ7aeQJsez7egB1ib6GL4MHuVR9
qpbnND87EaZqG/FTigrjEpdEG1VJQA83Qh2hIoEhqyURXgWdr3VxZgAWOk0KynNgRsFXS2oy+n6U
sxQ0iVFQaUiWiKDdWam/eSlDzW8D5kDYRE1YmdtXXq+WHUqW2b6VK0Zhu/HqrheMLJINc+CbloPa
PVGsB2uMKzdQSguUAgCu4JDsJ8+1wOp0iKsZ+5fc3MS2XaorBeAt07mC8PtbSSEFqg4Yn59yTyJ4
rB7imzeGpxwmkArHee54rUl0OAPaqwC6vyZ6Oa0aKuw07cOxL2KFgI9A/9sOJJ9F4J5EaIZfssbp
s2bRpImh4F+QMePgl2JOzP9xlclpAgXxOpNf03dMR5jHtIGvXDddHnstSYzOhwUbX82euP1nsisw
+Vu5uDRt9hVdydpQeiHl0yuvVWIZ1Vs917PKiEGOpXeT74bBY7eYuM/5vlHh6oEqpVd9DsnBJi9T
Xkq8AASOuTCrLz3hTLzMwbkO3Y02PVHQTybjFBzwmx/T4WNrSL7Y5Vvruiz8BdqwRV2EfPnEnsQh
0RzkAu6DtxHkLKCQKCYDSNsZTxrGrq4Foon0Iibx9sMZuG9nAgkS1Q2tqYWlyo/PgQx7YbnHS1gl
NWWwP3xVaXyMLYZbqlJgjBe3xd0s8MYaNI+DnIZO+RUoBtjCX1Wqtn4l4wVHP6CI+/uc5qPflGBC
bXwmTI9xy+a49ZjDfM3LykN/+xlA9avmxOkZ9VO2O8C+k1svg5ACyv6HIVLIcFqbAUFAZIJ5kA/H
dnzM0QfjWf7ge9RMvvoYHsV5V3UnskadpS7wDETXif9XFqklC9PCZWYPLSym0Cl+F/qRkuq3KMim
fRGCqhw3lKZMQsERTkuEhVmJrfDdir7p9FoTSDYE89uMD7f+QH6yasGELL9xhimLV5cAfjXceBcn
tl7sV2SvmvGm3ZBlDg17dChd+B+hGV0kBmY5c6GjWl1zqJV3ttHnq6etQyFE4rYMkPwXVInr49cO
70+qeMLW/hUaEmnoAxhc1psLZEBBEZI6EAINOvUg0jTpCD4Gmgc8bXLAxZ2528kYj05961oIKs5i
MX23uOefzVAsMcG/mxxZCn7n3jVVZkSeOEXCWsgFAwBmKEWVoVExuTyy4o8TrOU4YP0u2Jbduh7+
GMb9zbjCdlPdSRQwjrqJltOyu+vY4O7gdXNnsndSUK6a0/B15h0ac64vOsYWnZhBrz90S8FNFUCK
nLldAFoaROWAfkwObFnZAdgVhxPcrvDwU8Ak62Fp4rXZ/zo5WHlGS/ZbAbi4h3E1tvGaTR8PKrCU
HayPY2y3IJSl9iNx06TsmRSrqiZKvE/cPoE7t/Uq8sC4vgVfjkYCsqwVp892lvLhFLb+eq0bpyyB
UghLBc92V/Yx/4imKKY2EHxiyH7r+UB51hpcQpsuET5bOL1YHJHhfblA3Kb4IVfBDhkFB4EP41bF
vOWc2Ufx3Z8dNAV+L/0MyCpZOTb+lSkpwQKgT9BQeY/wXqBLaLD24p/tCzkq/en2LIGHUgDDnL4K
seFfZwXnnbmbXTL6dAy+SL/wSqw9DuUYIIsBUvE0vZlPG6OVrJK0CXErXHGg6pBEkZ76w7VdwbQ2
STda4b3YRKbt8g/UX0fKqbsEbEUV4UyFMwmeRL3v9/+o/mxo0lrWBeXpKyej9/xO/wOz4QRiDptR
mfygEcBtL2EFzOCg9zzMKHuQ7QhYqEKtQ/nb88e3t0J+elcOMwL8496qN8bY5WtFquYIP++TdmiA
7NRT70NLEvRu+5JWPvhkWhz4B629NXshAtB767jt5//Mc2V1hSnNAJZyQLu4BzO1p+wyeLFw0C4c
vBmKmBllklYDS9ikVVKOPG78677mtHgSIHYbXHbg0VjElu127bhZMbqiLRqj2MqzUXtgr2PkJWFM
dpO2bW90AgC2cVPIUEVkxv4JynCrNjLmoXg+FJ0ngI+iLQnJWSMpC8eZchofk7HSdnex0SxJt2Dr
n61mH0lCOcKhwAvgjyuUxnaAoReJDOyUPjJv8MyGIJHQgpSGb9fh2kgBnrfUmCCpOIk5LtXwrjfC
VWTCZZZ0CrAbnsL5ZZwisLG1gacbiMSjrrVdSY76XlmMjZIB3BL0HC7dHwW0oUJ4Ja9e4hBoHk5R
ZxqAVqVoxeAXnOtA+7rjd4We8lkQQKwiG9YxrwZGgMTkc3AmsEGgcxe4+kSiDiHbmPP2bBWNq9m6
oO4nbB2hXhldEBk3FEkd6RNDwLBvyz/STEJEXPMovUlC7W1F+Ak1bfGorypWjg+7ab4UwtHTcJU3
uDc9071j4nAdPTkogmr9YjyfS0yEuCKyBA/YjpMe+kMsYJIMtd7numCgfnYEOOE5bfHTW3BYRsCO
4GSobicNgTrRW4lsL4sQ0USD2oFNW2KAAHJ2EL3ZXDgIxicf0PrDfZvVWssOtthBLlepQxafk8nB
VtkFjsw41pWqNDkqZSZG92y7CmNT6vhNwwtVMVOXZKFimr/q7dVdNi/uFc8gkRi5I68p1I7Hns60
vjqp92LN86Ck+J3ibUZDr2pkKL4DAXSvZUN1qf18FDj/tf1APLWU9oSyUtQHF+Gi6836vA5lUAPj
REbIdVw9mvTHdFTxDCg3CyUZNTYUWzdaOYPGmVslin4nxkti1pafbQeXA4U3u137OliP2jXMFg2k
ATf6hYa3woh4vfOsIqrFsxGp6f7Ncz8iime8seB9NUxMk+xCzEgTTEpoHlV8XwNNqQ2bL6IOFRXd
udNnpbCifKV5vPYTsaQUC9AM3MJlNsn1RtyE1MWx+J8DpZ1obhSeW7zTeXloCx3vp0YfThZKIWTO
6kP3bk9kg7aPs4/gLj8fP6X+3YMkUohOBzJBt1uRwDHGrPY3VnkH1uIxB0xoRVt6H+WEzNCcY3F5
o9rBCKYaAsaViIQ4bVVL6w5X+RrtGSF0KNWBC7I0SiIQ4E34OAHrzOuE9OC0UIzv++OqeDJifXDx
7LKWB+Vuqso/OWJ5AiXd4nTQJwBtyKkM46QtQAHH2TnPPQGp9Xrpj4VVSLQUEyGGkgisvx91VwSd
/46q1ZfcY7qdJyvbClLs27Hu/opZyiggl55JUljStjWd9FQDmGyFFGEROH1+57G+zS3nVu0VIKyO
VmmiOWVuFR3lpnAvShRoPkGdJPvmNAOk6xsApRKyDYh+6pVIxQZjZUuCIHrTE15tSwfPYfDhNWwu
Dl2gRcL2sxjM1SzJJ1vqmbWo9t0DEz5KK7qgHXemAz+x2wZGVQHSyKmz2eG7bVIvSheI+gRy3Xn3
wS9X2oJnVDYSj8uWAizeFUJN3WZBme5CpIfW7uw908OgiNQ4f09vONAgTkOhqRup2c9wm1IDlRd2
7UqtJ81ponda+ZhfCLXhEhBpVcO0fQHBMZXV+ZI2OD9Vj+GSy5DsXuRWqbGBaq+CT+9n5i4ePWac
F12MCTIUoSTE4+VeHhHkjYQD7C3zc80MtJ5JuTiqRVeC9xVIOZ4GBTDxjubSgzRuWDTjx9UU2+kl
ctO+JzO1kqvAVMUPnVxU0BKFeRgorWkY/8L4PKXux4e5kjpu3PPzKNc+jV5cVYkNQ2+dh3p+4DHZ
2xLHaxzYl91hBuD929Fd55ACzHczd94hR5E2+umm2hsi0XzTk05a0eM0E32f3zmTQrKkUpoNxH9z
MEt/0ruOxieqTdvDDR633RtkdK8dGSY9lNz9CUM6hbrGJZM1ov7hJWMoBtnw0XpYQD6phcGJKXox
zkzodOjkjXC/1Z8WNuCZtoeHh2I/Fnd00k2Tw5ARg8VwUo/U2v7TFD6hLmQ/bLtW/Bru+e4I+uLr
uy/ERCmegcyriwaAyAIqFlud+s5Skvl8dyi7TjIFF6cZ05rpT5TdA3MEpnnz0XCdMiO19Cz+wV0L
tpHl0p/rM41ey+6sPKqAvKMU7kRAxRjecceuIdNGwplSukSPW5DX13XyMC+tDiZh1/ZpZmG9WKoQ
snTAYEviOIlzAK/gGBpgr+WDYTsv2nE+QufWWOF+LQSEFvNZsmf/LN65TSVV8SZm7/twx+X6zs1m
bXJvOhzZyR19zP+L5Jj/HN3WElFtFC/RsHpmGcpC5wt9JHh9xuwEqLILyQvcBPOhTzjaquErvwBj
CEgfBP1FDYqarM31DlxizobInamsGTMjTWZYk+lRpyQAUpuWUuzrkwJFaWiNN7dp6i8TkFtaJsiH
ZXnIYh/FRlDBTLnYSiiMBwq3ZAPgQ4vzmKYnH3IL2UFw1eRcR/k2zxfgyHZUD7mciUFdp4cZGYgt
rgne6CoFXXBfHw3Qk4ZhLsUQGmjWLPQ/OCUDK1IlUugKsnc8wjMjP563AYhsUw4uzqtSLNmS/Unk
11RkVNj06Pm7xbi35V5hYXdVCK+JoeWyqeobmv8fGELlW8RGbnoAyvYrKLjCnsqZcTO9MYKHRxBy
t5pgMc351Xp32Y+IHGCIsZg1SoDWo1fGOiUZC4d9xww2gauJlZZkhYJUOeoKVAkCD8YzJHcPY0LJ
KFOCjMmUHY25FyDmBvnXtSk6/GaeQBubgHwTwaITKADy6qLXaFFIpkgLDe0VMKFmEehO2ljFGK7t
KsIkzBBA1InL3AVy7nExT33aFwUi1wPPoCT3ivhHvnxrcO3eng4Oob4jH/qiKUp/jKkVdyfc9v5R
Wn9ANKR1qPgjxryweHdFxtgc2ZN9nrXOreuaIW/5/WHvyT1ybBHFaQMXAEbrKxkEXUpKGiBi8Mrx
jcy6RPEul52cngZHuz4u5ZO8nfkfw3f1p0z8V1bHd/o+HX7Vm1fqPnhaKGJtfsugNY4+EwmSGkqd
6EjCYrS94n4MRUxawRNKC39fpo4P4J1qPT991wCBWrQ/9zB7vEQK4q1KwjP96zU86l8vKYdBRFb7
zR1WX/+ghCdYsX4797MgU5DOcdjrfEjgT5m1rhblNIZ8Nfg3XwoyQGeLX8gy5foHtQ6Gdv0FUE7y
3S1yvcBGrVzICu1pSlt7/AuOaNXBG5tQLjviCxC43UxRH5I1cuUeQlp6IH/5IIP8/WR+v9WgFB9Z
I3t1LmPka6rZSRyd4Kb45PN/r56IEG2c3dojPqenZWPYPq4hTENujR2qb3IbFl7CnSX1MR1xDw8U
gbwwWR13FsrLaHVCU7yfJrtkggV22LZS3bACi04QXkK9s/d/tz3mIps/07Y3TIk2ZWQLwf6D0ECu
W3k4XT+yz9IWpf2Yyiwcmu0lHDm/5zTzL/lqvrOetsdpDZoX1/CWnfTURGb7EykEjqXmLEH58c9M
BMC/h6JLQZHK1PogL1r9+lQvT/d0LpJ7DCkqP7WfX64gBp/vJgCU+Ktb9hOi0SyBmt1lJbwTqkO/
J2Zd2PiccnICxdZ/9ZCogbgzP3DGa30ggMpXcct07PNlCj/BRlGpmCbHoXgqidTlpHbH7jDCIRji
YXPOAet4I4jqS5Kh92gEUrM8uFqnTyjax3OzwYcauCYEVNo6fbWrXfiS13LCDRmPtsY/ggftEUjQ
rd3FUuFavnKNxCIdBh03SfQP7hgwbP7kJijpRt4ZErUWHCHXPTPc9ys9E7+Hf23+X0MDycLBKboX
LacUsVV4EWwTeMnzxZ0hmonevlPAQyVU0xq5JEAVwNceCi1QEIWC3TvXqc0zFaA176Bda8j7RLUW
r4UQfugNspVUUFwfHd5CkFB5YG/Ee2lfD8zPRiTmPFvO7qnaS4siSCRnWFSmbRjC2o8BMlI3sMRY
Ws6wxQp6sNS58P3UzrwbYfGNb667fct1IaxIHPPSC/eKnN2Z6Mb78qZUtETvTg5gpkwzVqgNESjo
UI7nkO4rJz44sKy4/xHrlS5B3+e/7tDaDVW4vKWCuuJMnBnrei3Y7H1/raM70Op82ibshTjb9PRm
xHfjEGJMpRVJHrLj7RA+QsFiz0PX4BLq9f8L/xx22YyBw3JY1savd4j30nFyprWeMzVTsbTQj3D+
K+VL0uuD/pzRy22DZCnTyYuLQy/4rNVKqJ2YjFyP0K7MgYorxApOP99AlcL7NIVNYRI40756Wab9
mNzolCSMOIwJndJ21NbhDtQf6SKaDruKp+6AET8lGFfUcBj33nVtE391YaHfyL3Tx8Zu36lfYJ7Q
v5rbouPXKdx3zwg9OIQg2kLP70OIKdfPkq1hUdIC5mBqndpESLVeS1wWQNdOx4bw2FPDgrBh2aRi
Zx2xIGKAYEWhm1lWpKWmN11qLIN1YgnuMdi8D9DwD/h35yQ46xHSeTFlAgtKeqkqg++V+dlLxNXI
rmbTjVL3XbM6VoxWe2wi/06Ik+ZAnCzjBkIE1ALugTU3hQ7SeD0szxWc0yAYeqxABBr457C5nW9H
XvO53WTPa0lJPYoE29jN7QcQTaCeg4b7DFfhzmLktG7PghTdC6zmytSNWoBKrZAq4Dthrj6inXLf
JgPnOdNOc0S3FhiTFX+YLjt7HDrPMmAXhnot1yHBeeM1gIcLZmQ5R8Oo5ChpqmEOJiqXMpQWkS7L
f47ShkXA1LMMa9R8L+5qyTjzqjGZ2e+A7Tx13DJ4TDIj3o83JoeObEAtU6jgxllD0SfsIr4LVm0V
+R62VJChr8gcjeKvnrMU7hV7SVL0VsySmzvh8WZqZlD6M3otcMx6BQOBC/xnQTTnuBNHM4n7qz9+
BHKX7F8iefJC4e2oTFDePy1BrMnK4c0gZPNbqj0EYxI9ZucXsHr0Jmw28tLf3WC2a454TxYR0p6s
YIY9gZAfAUSflaKQKYTjeoEkasfpQnSvJvx7vLUPDO/wVTUI1hx8QnE9uXP74z7f98Q1tpaai3md
5BYMwXjVIjhAMahhWU9xhKOR52T+M9SpIs8q/MPENKBTi64m6UohgyEyzj8OLAlnYjoX0Q0GZZpk
qJj2airdGT0es/ueyOE/+x5mN0uQPgRKf/kvxHFFJ3Qg/FE46+b+EjyBZQgK5E30cCtxA35IL7xL
YlOsV8b5/yRmMhP2CBhExPEw8cIVPSA5/lR56YwmPK9MZ6SIx3k75J0+wX/tBaOSYQdc+SPIxOpl
U9TP30mzAmUc9ec08ZPcbqj286LHk6p8od1sINWPkxEn9GPopgYEvY0QmNCdUAu5nrZnl3Nm7fxO
uwu/Sl7YwksIAt8EXyFMnYg+wZD1qyRHuZtnK6xzj9uwQB0c3vRMVblMFd9oPaglAGEyn+np+mMI
EHqGytHfbGY6Oc/p8VmmRrEcHMLCxq9c7CSXHrxKo9eTly67wYQR145Cjx1AxWHclFTomIho128C
PUsfI1Frh9j4y9t7FAPIncI2VsKsvEsNqqd76NSvX63FIFgzuqzcFtZvbRX6ncKbN4wG9wPVUeI8
8c5ULkn49GJ5Jpnsht5RO6yLm2bzb4i7Mz7G6gxGPaE13RTJyjbzn08MAGL9uwxeMk0WvnT8Bg0H
gt73oGRwGnpIBCQT2KO932Rr2iqAVUEx4/80+xIYuhdbMjzuCm1AL5qkmQz6WQDeKc+8i9WH8jeK
jT6/wv8UgJB5VjCegl/YzObA37SAszl2WliJ9WwpPdE5dVEHbdMIdDBOu+tph3bZqkAM8v51+liD
mSQBupwDqbYx7iDet/PM8Fs4BJDdcux/PNXCQCsnocCVcV93t+ICPI7DS9wu+HsuuWwOl2cr+ZTs
CjhELxnyGV2V5au+2AvcyahieuFGOWIyYpDglkeihw7xoy3QaYhVsagpAApO7vKN+mIb3KXmkF0J
OwsP8uT7+F4E2Sut2ZVHPdpCI6GPBUGZJ9N4941LoTS7Qc5zoTCqLpIwi3CuOLqBxiQH+ua4CFWQ
UcwSNc8PXR/0lYb7shHXVzDndgcIqaaG9+W+hKucrCV3M8aFQQpz/hS8LmeQL87JtcYVxK8UKXd+
SZXq119DDoNquqWku/nTw8VPj+M7uGp27wB5uVin1Izg7JsLtW/Mxg2OnQWY9mB4/4nRujmqYgBB
t5J72wrMXZE00fUOPjb22kXdfHVIRNTxWKXEZ5GRz7zxRaOIaZQ5ilGilheTQWq9/0Zui8drKaTS
0Cl00wclinMqz00IFyIheiqO7OrZS/56s/wg1zFsZNiCuadDDy/G4n/WunZuRTh+TW9ZBHkBf6tl
hLsJujl4S5MWoS6fY3fb41bWepT22wEclVr8oDDBFtmCPw6IRswnHCxM7vSTZ2EOmZB+0c78qkjH
lqG/QKtBrgH5BTtRL7/w9mSdSeITXTe6XzRD3riyUGHjWUZPyIiL6a7fwiqs4/HOcYXgLLsPl2X9
n+YVR+Ew8Uf5NMslNEhOb1tn2shI0WSVpR0dOQjtmMkQGuoQ/EV3crWixQAB/dxQOQMQyLny/hd0
0poa/g3w/Wsea7zQf/4p9Pr50O9xhLOQ/IJEGPWdyshtGgQU4+mqmkDGDEKVzoAD61SQnCQK15si
lKq7GwpIbK8COLcgWkScUq+puWbPAmaBlQoMqK7A/iS6IdsVp7azH8/totewqe/6Gp7IO1HxMFr4
q+oljarEmDcEJ2YlUeVWA5fQ0oEitx5Urw+8EsKXiUWkLsKZp9dawlgNy65LLZBH8eWj9rYCTEZq
oIlVQU9+k9vV11O7wN/OQ73bMiwvOFJudsW16zTb9urNbMJyau85uczrPFa1mQkYDTmhZQjaMLu6
cv7okxJ3d2eY3zoAg12JNcLsiBQ+ie4Aab4c/ufUPBXT6am3XAra3Y0TH5ND79SG7tEfcfQCWlEZ
/RziMD+VoltyQbv2LVeIHTZdXDIM80SADPg8DSEybtlLPaSZZosR7PuuSgUZmeN8Fdl0vqUYYQgw
9Cnu3k6CF30vwbbT8csrXd2nivtiw4J00o9vUmnr11c/BlNfA6t0ZZz9r5QeXE/OIZR9RDZ01gQl
4LxWGYRwVdfZeZRmAm5W48hTa6SaLmC8R0aAlcLbLcFoqMpTDnWllsHygHdW1Y2KajZtgfPSTu6t
6HukWYb8U4A3NGJsEguXwNMbBS1mN7QLuS8iVQze8CqaD4zmlMzCyqtQoJgP3MaXbKWUOk3znwN5
GL5Va2PXT64tvCCotZwh8uUymZySeHi4n4EZ5WN8+FmF4NgmyHhze+COXHBYTCLZCKnyteX95jCV
pox+crW81eptNdgu3lTFMnsI6hsaP9XM8U4ooF0Zb3iIYcRE1J/3B9IPyDkKIWOKs5iPZXqAcd/T
WKrU4OOarHo6QIXjIw2XtoFkzudp/P+764X2UzXJkCbihnILBQNa5enrhmGrzM/dBayu0DkBOuTu
6Y9PcSDui5+XDQ4p0SGeOwUVc8n2ECas8a32y00gNRnvNxz2ZrYC+M5OUrIn6QIc2FP7oxMHdxvm
PU0CgKj8EPrjHGVG3jolQkBY9dE67oShiMsMWLBOe8TA5rU3kZYPUDPsSGfMRaNSz0ODtFCBLUYC
x5ywkcYh50iLaRidcdNbIwDcv1vVqOnD/Kz41CUZrjSF1iVtMGeGVGWaZu5FeqlKuZ73ud2Civkp
T+yBy2Cd3JCLlzy/a52SbHAoNiHJPa5hLsVPoRaVvMZKG43YzuiK/OATYsKKDCcSH2CkO04h2ciy
cxsaRCtUdN0PPvmIUteJ6oR32rbAakaXmUGIbg9AeH5M2vTAwk2/lWZFVMo3jgowP8JN2ZYwxtOm
1ouM40eTa7MAqWbWwU2gkCeSs66jCk4+RkQI2cQlLxvttFU/eu6xQhqr6lEf3o+Rq/izbvPV2Dit
CCw2lIxnBrvwzjdWfGXABW9IEy8Wf0uma/YScMbJHimSBFKC/2PBwY6k8iAcTOiZtmorskg3pmOW
4yzHllJqcoM6Zq8HAZJNv1P0slHT4bxkbF146vi68dhWvZNfNQQX1dzlFWIGe6+c0aHkO8xMcsS2
465F5ebZ4Wchd+oL/a5RtrmCIzY0hNXyRIojocOWlWcd0a1Q8llQcmPMtUmSCqVbsZVsHOzQygPC
ycNvjPwjsNG3km+0UX4IoLbpHk1fRtscnDeSVVNLWeM93CpDVNQ3SKypIGVgEheUTt2PRUmsQN08
rzbuptFr4000S4PYPr7Yzz3f/7RbUj97xFrPH8Hv9E8/yNCFaz7bgTZlOTBFr0PdLelAHDVz7n+T
mSlXbfX3d+dBUMbYtO58zP6waZcdn0tmxqOmyZr05R2i04pQzhpH/fvoM8Guin03cm0rVcJRthaU
6Q4grsKXwnoLZ1aF07I6HJ8O98htBjlq5dffONPBCZSy8KK166kL1KQaI998uwpbjrndETBbiykS
uRxbE/Ey96AfFE8Xus/6SqXomi5RAEOh2+icaDO5EatJfQEc8xd7onR6bB8SHMF7i0HmRVF6lJre
xnCtPnGeiPYbH4YTucNbslHRIcYItuMw+rFUXgWcVYgq58JZNH0QE821C12mT2YSD48e0uHMf4SF
h33ZpgVaeWtuZ/qFlSrhMFmXhwk2COopYP02r1r6cjvGT+y3Uk2nHSO0ejpWplA1Ic1RqWeNqirT
SvKXsHq7ImH3A0CyG8z+fDeUQFg+9ZBcmyGrfB6rUcPtWi8sAYZ1qfpTxucrf8OFogE4OEAEDqfp
YTazfjqZxEieiICTABpOEmvalNTUW4KpxSH6fz3ZF8+XznptLh0Hv/Ea0/OwvkhziBZIAQbHOvMT
s7p47celxLqAwaxmMp3KAV0pJnnbKL4iqhATSNlIk5N1wlQJlKs0kMx068v2JPrwdwWxe0HH5yvt
rZl+Y/ILyFG5fAG10ZbKFHL2642HKw6RZF9JJJZOLN3FU6Z+Px2PQAZe3Jl9lqtMSheB+r8RgMjV
1lfixpTjeXhJTWBXIBhvnBrhXW1w8W9tpyVUnNwW30TxR0PHM6zkFwIEizX2DAC7pE2UMhj91Qfn
hC/3/4IQQA37Omm1KgkWjnLGnCCfzz/otWozOGiMKac5KlariAHDFas1ULWQzwST0U4VRg8v52Ic
wE1fzUYjg8UTh/i3BpWuVQ4GQFugi749USdkTZ/WqWhSNiPwKKpzL7Pny66rGOXm4mAQnm8SN46T
rxYCxojFiUjJitg5FVqd9vKt/zCcQoPhW7DWp23AhUZaRZvVvBGknYNYSXq8xlyyboCJfuAjNNWJ
XH7Q0P7fozTi+hMhH+9fKRToKsxbZNHIeeFwyONYRaR8F2AMyKBijt00eabAX7Q4vR1N24CHY8on
TtyfQdRdEOP/+k0/cx5wX9RcWWpdzwrkVAmBj/rhxnOBsaEykJzvUJ37+3EiCUaahKgk88JmbiRr
H/RLVIREQgl0r3MR8hT9hvF9cKxMRQhGHbhy2Wzv62okeUwKMSg3//Q0gMEi9QrDSJLPs8Vo/47l
WapJ4WyxaQBlimaKA94AqZ7GpSQkFA97l2LN+WhfaskFAYwUqtJIDbH3zs3AeL4AYdHREnYWLfPI
doCZSZtDBuneckixp3g8XKk1ZmiCsCh5d07WkRPh/OxgETMmstMO2PfiTyUv7q89oPk76g02c9RM
NLBpSZQ25nmksdPF6cKNFdT0lsEcHZchbzQh9KDk1dh5svz1WfMaoJffrtTSGVCS46Uo9sPEbyxs
tDE+uCRLBTloMCJw1HJKVPXhGLgXFsXMSsT7cklpE7SUMKDKwYWwuHOH7ksfQnjgqQndpxpE9fZb
PlfqEPaw3GPGmQGrUni9nP4di3aWs6YDGqh/pGtEQn46tQW/tt9j7vi2KW6o6WZGHV4ZgcjprDfI
tUlC1owvxSaSBBV1RKYRAmMDnR6+OfMjQ5Qqdvr0tz5y0wCj852ZRdzqR9d709co9aCrmIhVgbJF
hXy9wK/Fu19fUUufOO71a3rYv2ug7CpsKXWrnXUHF66Pd1+fZRQkbBxK4DgM/YS7+hXnVh0aOXTw
n1Kal5NU06sIHAn/eOE1AcQBm99nI/aqmW+hejtI2pjQgYeDzUXNxb6t7llAWLR0s8HIZQ/5Lc7q
7HoUTiMhQ0818384O0YOkKmY0PKZNfOJUAOPVCP1j/viVFknFyeOG9Nwvdfli1D0IlFWDHdZRIa/
Ogx05t0EaJ4Qk4UK5SwW0AdCyKp5+79nZcnSLfeKPspL2cE+qf6IL5xE+2UChXLivkxzaTWvaD4k
qmIAo8wh+213/KqcVIZz7XaeWsV+MHWXwNxbvb2JM5NPVztVJc10+OerDr1Btnnb/HfvV2K4AuPK
AwiXn1TD7XXPSHX7d7IdiYqT04wTr+Pq2/r0Yvw70wSkPN/AAMxD+WXuzkK0tB3O26s1Y8pfUqJI
pxFtDkWazTgULas5bWU6CBWxszUYaYOqWVdNNHBxynmgVgYDHqcUUF9Qi8r0McanUR4kDVEPDFwM
2ae4hfFf2pXQSxYUpNxTMg23W+ZeN5dWljHEArynMkykMReYadJEZNsQBctub280n7Dqpr71aLVR
VAt5eNmQXbqy3hIMsjpX08T1+bPnwx7ALbaKb/VenUP8OC92NhDxinmfrQWh0cxDgeCblFOsUYyO
ubZ/0iiw3489suxzhg3RhemhxRPctlN/RQSX499qm2JT7h0ZvX5dA0Wnh+jfFSF968e74lJyvAIL
ZAxmENI6CIYcgvryB5C6J/0rv6oNwFqkzxxGirPbDAVbDbc0u7s9S9MkMHbU3Ufrpc2CUtrEgoLE
brIA8FBkgfNsVci5IDE4XmhyYurUSkh0zh2z6yA2iQIiT3+MORmZ1XKBBHPr5UtUVs04sm0XBTLd
kU34TcgrZlO1s0VVRmRUZsbbey73xKrZCm6doMBsLUWFxUTqTR2sgBqAfTkRt0CFglC/y2n1ORci
hXb8nNyF53Ti4xF64wJheKvcLO8kU10uavs3fA884sgtWFxb78dKYwNadK4JCDiSV4lHOnnwDtzQ
yZEuL2FN6dS6o4/st9s4wzfES9hBRjTsDkKczI9t44bnAUmL6sYeUbK2bB43c7xXiMJJk/lGTYS9
J+NjrPSjvtaIGCid5CBq2aTMAJ66oW6Wr1a89C8Owtofo8YkW39mrEeG5kKf7zRojPvkpa/1XUP/
CMnEYVpwY0py8bXETdsUV0fKyFNeZXJHOFVV7xjoMsnxKNWqXTZiWPLNDGGZPL1TDykNp8PyimGO
RMWX0FUkSacxf7O/CvvqG+UVlOxMj46+shnVqdNNPtsY+3iG1MPNhyv5/xDWWPNyHbLjH7g3bAfm
DuOx+63AXLr5sxScmheG1fhT8ni3YXjIz4Rr2+KzO14rVxWeLWkgqcZ2elV6G/3vQwVnk8mA8BUe
+PVDCwOxXrgxFuwDx/LdfOYHUTuZbHMYNFhYL+XTZrpZGQzzps+/eZQ95MZ/Fe5M2R34JaXL1v7E
DmiUreqG+WYngUWt3UM8wClj1OC7fKsH2nWMfKHo/l7cT//BQebIN7mY2u80jxSwnWw/BUq2e3AJ
PE2hDbP6j/A3zGcQJe0zKU3SVbdmbGrvPlUMm6sKoui9NRtsWZiFzywjDnG7fIT4DkcLrZWE4V9n
l/XSu2N50/zDXg2vD0/leGzM1BvTSf+ekijVgJ+3BVJnyvYkBKbs5vYSUrcGxficssgBnKAziqfY
CoQ37nHQefoyxGh6dTKJTTcFVvapyXMSxf4wxR6QmEdTAOyhsqsuL3HiFLRPgnA8HzD6ziNnkOJz
U9xooCz8biFMbwq6DaaMTgGT6l9ruuw7QLZGDr18vNs93cf9HrytNcLxCCD0RFzV4nKKfUxG8sJy
X9n4sN2Gq9MJr7heL1lzVeyeB1YK94vKfzKh9I+iTieRESnmn5r5r3NESV8Drhc/Bw5uwElx0umZ
qGnqLprc8dtnSd4CYIsvNT9n3D6/lUNlhdW5YZZqz3PWeHFHjRyhhzdXm+b4WvQmW/loTldo8ffz
i/Igz+V4WMLovONCkPHDDkJWL+3oYp4V40Z8ADj6kjAW6WYptbHmLt11SiLNIy8Fw37WfWbeiYhe
12cioHhYnB7YnPa83LeIZCB8ArXw1TqUgNkWHzznRrm0ZaS2rzEqfavuP5WkuHiCu1LGHdnIhnWb
/TswW2PWLkketFnwQkxXC2ezKFyYOyxybaaIDefiGSUZqpV69J6elHcTeso7r6ZDUQ/2wWaYcy8H
hvUqYUci6dPbaBSq2ZQQAnxYZN9X6RIaoa5lmKqUnHqUH+H3gVujs73LDTJ2CHsBixXMs7aGFD0c
xwO+qi1GpPxxW7W0MSVn91zayvu/PELJJSpU4auIfp8nAdVh4MVaLIQYpcWcSgqVMeBQRER4l2Bl
WEdWt7eTR5XWwBxjRuTwaIdLYZMQ22/3tvExmpdsq0mmTfF/m2efWIFTXAQr9Nm+VKB74pKpSq4c
HI6NfYNFTZNi/YE8BSp1PEch/z9fY2DdbF4iKmGKia2+KYSsd90ynoOWDP1dNX0YU4gsKZr9aA+B
2gB63Zbyc5+pV0s/B0GPFEjNQ7uB7z6f21iXN3/+2Li7bjXEBrRd6n0+ijBWpbSNvKbc4ACLzeDa
jfVAH6MCBdIWvk6a6/TZOfoD2pNzk50XJhO8G0aibas6SjdGr7I/gjlS3ArhKqe6J7AONEqdotHP
Sya2RaxFuhUGv1YZyWCS+yZ5WzY7lHaO6tWuUwm7mRwNuccSGGhJQM+LirRL8IZvj/L+oLVYlkwY
gO61DZ/zfW8MRXcyv2fqTdgjT5TcZ323JN9LraAggWNDienlfeIu++GlUcklIxlGYZ/Q5mh7a5qd
+EIhdgJrMyDcKUNFvuTltu0ckq3XFpGrf7RgoW0TRE7utTO/yXv/o9C6pZTEej/K3IOsPzN/7rA+
X9jFT36BhXHh8XoqVWVfI27L8M8FU5jABRkGZoNabbfrCVJNu7p4ntCL/KWoNdpICPg3pNVkcBc/
zLG0V/V0LvYPVzQy0Ke+I3+U85wMB9dMnUPdAeSOtv/SW/kfT72d7gL3swnNj4hMm7uqQjA8eskl
lkOSsQKP1TQExZkkfug9QXsV/nnxiiPRiStbiY9o9lhw9aGvyreVU7PplRtIAtchMzwoytH9LSLd
zAFQjuGXU24wuFi9LNupIPhZgVBtUC7zEiNJ464N0dG6Cd4hmkkuocnVRtUopp6DJKQeqH5iRLnN
B2fmvwQs/pLGGyOrGBHPQVFwiD+WLCO2joWvJuYWGUEgGcb6JmGAY2HQbkATTsRfRj0WYl+2BSTp
s+vfyJ+Vd9v+Ws/u4axO++ec31zIfMpJhvnnm+Np+RtmrzxtpRj4+SOSCEJedRScARvWSJq7FG2g
W7VZFJvmrYFYA3bHvMoNFJ83LYgXqeQ9447u7w3eH2XeVCru3focQRLuEXMHXn3xXlscTd1qy4xj
Mm2eOMqUnA7MdVcqTKD/10tiQqfMKqe/ELXEXQKF75RehSPb+bdscVHw9dcrwedHjcJ07YD1vO7/
yhbvT+t3ogVQv0vs9QsOSkkIg0lYD3PyCGEg6XhXcGDUDDWmDN745tb+GoelkpxjXLRVkTTGQj+N
VLfHDrOO132kdWkx30Uz/revGojUOXSG8gOPa+zK6i5+/YtcbFqWIwuYnO7wbhIX4b7T9zj2pu+2
BGo0vB+zVmPaHVi8VMImH20nCm+vtmmgE88qzTRjLXC/EoBMRRiX/SEFP8QnpAyln95jHAR0CE/I
pt7jphWI25gulUC49D8hCwcsi4pIzpss4xXU19FsTYqPnEdKjgeIPmkDY+ksyYQZIAoUVIjVer/3
keK7oQhNiHIRP+hONOc2JlixcFzwNjZ9WxMZyHlvr63ekY4Bed7p9WhSUf3ZXRCRksKzh68m3GqG
1E7JZa20Y07jlVvMZwZmTWo6o+N+AADCxV6VWu6WjZ6sShNiBGqARjtiSbHAG3Juoj31y+7E6hMT
NhdmCfPIQAVFUy72wqzIkZqbscjzHaSy8mA7UuYengJdoym+6hJi5CTXp9c60/NfFus0gDZ8/luU
eG/iM3dSu0oEkMIURQTwJ2YnhPMpX7KkV5BsgMfUPme/fU5Sq6on5iAwNUmTqwLc9Df4V5w/Qptr
X3z6cDDM71JVphbJYefd/dv5+PESefrhR8uDndQSVqhJjlmQQMZU9ljzS/mZxlzrmh89tQkJIuKZ
J5vA1W+54Mhzyg/j43MpeGI1YYbyF3TodLkzvgmzuC0++7OP7/kolIgdqbYWwS7XYQY50kaJVQ5a
hG2zQ75sP9kIKuJiNnpiupWDove6L+S+qO6k83rOKBQe7XGfMREt7q2BSR2OwE4OdEbi4gmhbw6S
W0RoBXemw4hZrntt1QlBvKclG5oMwAoeKcUHh9h1Jd6Bd4fFaB+koOh7mj0yf9mRWDmP6uV/Tpsv
9lK+nzKtEjIE0SXbGjS6RrsWJUW/G+RyAJ48eQy39T3AOYvOmY/s2pTm4pv0iN7zq0yhAjuJwrUf
lLZIIp+whiqvU0tX6xvnOzm/s68fOMCcidALseh3ARyD+YKKZ6L7BkOfMwbgFv0Nqtdl9jTipMnM
T5tNkvdmi8gPa1dYJAX4qA5qxRhtapJ1jyWsK+mtuATGezfb9XlPQI6fqxOrv+DhQbe0TDDKPlf1
u1X+u5tPqtYaoHpZNBGRCMB55BRvo7/dVmgPa5Y8OVEdWf1D33/nhmYLxdcuy4okRSVMbGe4toUn
gXJYPELA5ASTLRoGmj2xYGJNPjXFyfZRZ7DzKlUsqd2maWJvWqEes4DesxQkKexjMXrrQ+F6XUqi
lOzyVS77tj/hQrLv5fKK8tuGpA5SAlAR9IoNPgp/hHVu0UkxeY1Yq8JqJ+TkXvKqGe68tci/14Tq
j1cpUKVoqF+X/TvDzd5o79fgI4OToS0O9g2KD2Ka7p9QDuoqK6J0aiabMMQpawaFSBskBoOLagwO
3q3ULhbBCm+oOoUdx9oxov46wnAKTWEIYWxjuVoJl9vIwnPrTuQA3kvRRdHtH5148ODRGnbvSBC5
ulMJrrgdzc3i0wu6bBcjTY1mNvIOpsW8cbL7UMd/IjZxvys0rnpH1v2zMF7yO95zlgGtM8lIKA/h
sT48abN2hmTfZ/qZb9iWU1L0iiSmF9QXfapcZFAcDq0eOZSSey6UnNFFJWYyTawhIIrwo8GzUXds
ZYXdmV+gLecrAcxG/aFusmKwjznNlKtgRR8vVUMNILpLagZZrm6W4Gkczb2BZPgYbuM5GxPfP+xX
w0qWYPfPGbEwmNEetxxUn2ClBiq7M/fAwYWgNft1qPxHaS8Xx7scUFAmUnwBJs21/fSi+o74Rue7
44PCME/T7URGRTS6tL+uMt2KO0A2fiHpi7EQYyiC7K/hf8KVHBPJMFmokcxTRluYNfNJmuBgFfD7
hb2kFnnVQsct72vsusdQ0swkDZknHDLRIEQpQs+oj1OPqs5GNEU9jVtORoCHY36RikvmciApvfu5
TQqQhJVBnGD8gu+KQeNYpCAw8HEI72gPFMSsoEBrYXArruuicsibQBj4CiDbS8DspvWK29SJp7VD
zTdx4Bh7Y9eWfELfGMby3OW0JNRug3FkEOcMaNOFBW3l3bIGsTXl4Qkq6DAa7xN+gbzISKwLP2aR
ms77MH0/9GqwgfBBqd0Ny2fxQfET1WKALYJ9mep5VI7Fe97pMAqvdmQDYOCUaNgzknzu++I3FYjl
5cBKjJfVJVNH0+pNTT7aBnJpZWY3r9IBHdgdB6XCd9kUqIZt7qO17nA1hLFv0nbNPpJAQYDEl4qY
vJ1LIIm4VdqCEGUtE7Z80OOU+WpU/GpDaixgKeQ0Omv15W+7+ZPk2faeQr2sEAJVGQZCii6Uol7p
bg7mASmBpucslmeLrpBJ9R6P61mclv/mME9rpWwCabTBJgQ7bpSgez1DwjaFGobbstIDwwbZFqVx
zB9AxDPm7yphRCExOO0xV3PU9QlgrXt3ThOK9bpRobgWiNLGEV++orAvh7TQ4VAb53TVdd4rCM44
YX4Sw2tQe3kTdol+3uQM5MNllbjlt83ZUAa0qLwr+z24eMGXJ5ncKYtA+tPTFI14T2BDDvJ1qRjV
UiDNMSt6IhOvzQq21Tx9oVWgv1q+4/eTBWf1UYjsqS58sX6nAQdKS2dxLoxzuadVnRyCvzHvjqeK
sj2YwdkVvaf166tB4AE7FiE1KIf8X5TFC95BSXGZ3vXhvjCcCCK+G1parXV0KXVPqTaRyD+amWcc
NVmNWH6HOUYHx+p7aD6uN6LP9VcOYpA+MshBl4dubi5LBZ8W3DF/KPjXpW5m+JLDjSRsFqazumbH
T8LvhWXCt1kPyN/jBrdNS3vjMlJWRhmU8HRK4mnp8m1X54xS5yTU+NvYW3zOQu02Zo4wl4XkKqjO
tSVSaoFJltfSjnEDG6sjfY6PO5/W6yKsdmp38AzUc/YRR6sCAvhgMcWB05SllgJraDr6wRq916jT
PdaVUbj80puM6xtNMVIxXKJ55Wus7w8fb46fSneZFSwggJ2MdeP9rK4aoj0/6DHhnsyniw0dwE6v
FMBCjySH2aeZ4PYs0QBpo29wr9qLAic//Q1jl18lGyTYxZbFoUBaNhP1ChgFj0Ux9Mt2G7rR9R/x
DtUkIqMaQ9ytjYCnfJ6HFG6E0a2zYyqxc19EL6pV2MGuJa+3hGIYcLjqz5bEeA8nwc5JswavyG5t
Ei/COUuIsghhvYL3/HtUxomOd/4pI6LR0L+h6/qXGoUggnm85LRsh2uIMYIjU67W8PF6RaiOZZkB
N/rCxyHZDT4myel6JQXPTLfENHFP6FbvPIlr0GErCC/JQlQJxVKaFCWFx4YBNWMuFmKz/ZppX41c
3Vqw6SObtEvs6TJ5zo16h8KMchEzc5a0UcqFMmGTM+HotS6G82OwtovSSLzCHWIB2XjiVPHjgQbA
atiYneUqCfNm459V9xXliSmifadf9gn3ustC8cndMP2MzQAeXujUXZogfvg4NIg8Hqxj2WGZaHlr
ZM5JpZXZuBy61KOyo4s71vB2Y7M2Lmb6e2qACV4BtVVZWoIjkkXU9TF8PUA/leNrT8a0vxYp1ooI
AJTSOHuNK849c3mNPBL1ubTeYqTmUcLIJO6aOr+pflq//+QoxvXnNq5tvOPb9jweBMZszyJ6y3va
kEJxA3+Fx53FdQbXrwVOX9rNS+eRNzWE6YXKqr5LsUdArUrq/TCRascnQGGt8fS15IPU/w/ucpsG
BEz3la6pYAJf5g4B2pL2t5lUXc80gie3f7ZIQSSjWSeq2QJndN1rZMNSFVM1PcGkwUegh12afLPh
PAauR6yTs0iID31h7ompyryD6lhUTI/KplBi53rtdMctl1JpmW2JphX+Ujt92cBCiILAlNTmaMWG
lrwTA/j1ccn2ruhBYptI1SbddG3hwljBeuGhO0qPq5TP3Ruyz3Xw6jboTuDUcsuj6Vl/LVBlL2cR
2Uw/ehbs51LcGR3fxXRODbpcptb1TAtwjKJZHY7lUfWqdKbM03sGulJRYFnA6Gkc6DYYwRb/paxW
bOW+m0jvhdgB1BSRnKNdzPxzzMiTnoApOu2uXGp8EgbRgWghG8Tt2JU0iAdQpE2EER2Q/0AsDiIv
gPPgq6ovPKiYz4wVh2OtYu1NTS3cfQmQLrWY9ArIRVUBIgiDEJWjhE/+5HR+eLPGa8vARNpcBpo4
X/8VYyJzoiTIpYRaMSnYdEP2ypYTZKVbDA4AYK/ZXZp0TmJVefYgNBJEkMBiGPLepcH999DBZEF5
xcm8iR61MDE+xPj+tQbbDppkSk0jYzy2wS2iybE/Sn9fSPCH0SE8IwaloR6n9cFSk2FoZdPYKmTl
gd9mSIV8IHfsX9MFOlSHd0U0thNkzo3qtxg3wGyL0MKDva046Mmg5Cj007112nyDATEsjgj5RqED
BrQekCxoc4fN7KKpX/GgNLYOltnpz6sQSFL7n4SrI7MhIgYRE4s27fQ557F9EVP9NzKRMLfr0S4T
ciPlXiJ4Q9XFkkotM9QfBckgTOKZG6an4AdZsLZ697R3RD7eFB1HRL+WFXNJ4/xRrFDNVh3Dw07t
A1Hzlyj3xDoqintQB+8V1z19ULutJmIMEV4WdOCpGrr1bYYPDdGQ5vkRrxDL4+cB8joqct57CtPP
DpIlDPN2RGU5fF6BqOASI7XgwunwgsZc/AwcBpc4Gg9P0gAjmUAS3b6jD0N+T/A05rHafLtOHrTu
2AtmrY+LI6xMR0Fh8WowVpm9AOoPQhn2HvxE+ykgzRf3sIhFG/dRaQDZe+U4Dtb9vmOHS5m0ETX0
rTtDd5/HKOFME/6nlzj2ZpeH+g0cpyiatkgIEIGbyrQx+A2Y50/UgCvnsi4Ez2dPYHvGTeG7K5dw
/ZFmFKalSjCeVjRkYbz2dmFbmD0fRWOQtO1b7pcCfv/DgaN6qimvuLuH3zl3yicEZJxtocNnWKZF
v5Ag6ASqH/3fdSkHdTy4n+9QIvWqcT65qCyylvmJGd9RTXMHUZlC5+bzKqHBxM5kpgnUJXeCk/CJ
L0XciTybFGW/Z43C82umK+b4CbCm0AytF28O/zZWZvOaHo95A0nKtR0fzyp/oB8msyS+fuXdu81s
BigGDKnux1hXFxTYY+fOOFUxi6tHsLtwAxXdRyl+bw0+WNNJTmqt4MF67AdrDIP6umk4N7apb9L5
DJEqQ1DTGujRw2hy/UtJ2/3Z3H+/C2NQ4b4/Y/J5cPzYV+9C9wfKsbRJ+ly75swMaQmNjoFUhPAa
vBEQaakscVUfUWlbI9Ufc/D/spCUG6yWFgoA9Q3MyoWvqEtkCLAdamk74wY6WqnYnkiNFqAhpmxA
qvuf83jLQtpO59LMAoxnC6MFmRRXygKiIYzohMi4lj2qyzrwmrlyV/lUx+5j9Outxvp3DLPEIlb9
QoLCIfQPajicTvFipYLMuQF8/ueusANxkCGqvlRQpDJXBvO9cPh3odooYSyIwH/2iLvJkdT8Dyon
BWqsW7yI/gkJK7lDAQvfPQQhA7au6xibBh90E1vVLokaJfQ2wJbG87zmDUAR3ILs5IwB0vzwPoZY
2ecMFQRrIaQAFDPVju/DzKd853wK4hubkwHanH9gRbclB34FrKLXCvixwnpO8hmFQtpsJAojim2x
eWViyEMLNSjd31PNq672xPSOHzbUO3PwNH/ncylNkdX0wfZSlMxOUhnX7nGjRUpWP18FqzEWIfJ+
VK8MIcsFGKjhDy/3yJKSTTMlmBhd7KdQJCZ1+PuUEZWtjra2WKwjS4/XXtQGD1WszmfyXaFD9oZy
gh0UP+DDqziYlTelvMOlbhMw9zph4c1DLTYWIoh1rFXDYkF15mgAHZnDauI5NtC2l4MjyxXz+Cyf
nN9ruPHcKfySW+8kF2Hb+N5BKDjUaYfbWfyZMm8WnaJAgUXQiC3vS+EKV6j2Qy0LGgY59Dz6kLMt
vRjSTykgezcIAG2lqJgiK4iGbTC6LDvS/i+lz/6LghdmcYKpFqjNafGaY1qySTg0bm7G3sGuYOBv
Zd1hay0DF++9KwcDi/0TNNJbngHJ0RTeAqSGAA/jzPfGCKahMbD9BhDQwE/JLeXhIsyMWqrxp+5p
+NxK1XMsy0/+6zlOGiyNELCP3QxlUvqyH1j7Uhmm0Rre3y8dY2MXzaslA9yi7devUN2m2lGdAq4u
ejg5sgPhdHUUf7UiuhjGWFsX0sdYPuN5ZWcqIadKmBiuBCrr3uTGuVxVtg+QWaAN9xYYvD0tcH9G
UBOg99nX5kukrrfpHqmlMngRWy8lfMTZ+0wdBe629YsmZYXbLCvFm2pYkLyrPXMJoW+m2K+gRZEe
wYQKldXcaN9icE9jRC8EXRaiCn7tuJIjIruu+Tna0R/oZOkT+TNHOLIFvC3jIQ6F2D/+0VVPpGbG
hMTZOzAwZkXsn3m6lognNDfYPG8CPeURnsWCQAN78w0YP9RiAGX1pZ/OhQB77XjIQcsC1+u1X/0l
dtDYHuOpjULcoPlcyhqsiHrv2UX9H8ks6GLJiBlCHmeML82m/z+wBSxFd/wWWgNlJ6sGVtTSWuD2
kUhI/5pvJOZ3As8+5EnrUpo5f6+OSRwZKEvq7P7IA899r2W34PtLsXMduYst0w1XJcNIirk1ml02
q7+cHyy7C21oTHaqBZMfH6VwGDB7aehTj/GXWOSfie5yXexa9KW2iksA8Ts0ZJaGYoymvquzUwrl
se2F9bpR4Atn4Snjdci32XiK9N5lx1aeYGyBDGe4LxNggkfOZPH1+Gw7//r4QQX9dvYW1Jl3O/19
VU8YmLZncfqbs+UqGYYuQfGwz+2u6POQMj0/kBtTv8uRflIaUX89a9x6htpy+PG0p/tGMT1vUfkf
J5/3qJYggW7comsA1fJqvRuKoEChvMkcm8J0+T7eBz8rew/ERhbZDz49DlljsN8qUJ5Rsh/IbcBJ
C/aUZ0E8DvmF1HB/XAuT6I7Picc907qQEN6xPk48RZVZ3MxwJc69h3ET0dnfNqK/3Uv227HeQYmA
YrkVzK1aijo8haMJPNX/RjZvg7FOljiZfjWMmpYi1EBdo6EubgjTFLRq1cDlRIH9v/BcnSV4VU+6
eJYesSTWaRQKYhu+l/TOJgRmCffNKZjX75ifTqvFG+rQgmUPWLmqu6K0RrprzqmfzN/3DVZbmoBN
L3E+BhtGElZCMMtIFXqpLdK0wMTdNAxU6H2m4f1p+T6WNmK1cItXMuq75kl1xWT5hWygICAV5m10
Yvq+wMrKOILFNB6vo0hFaRvg6JyxNzoCWhU2Njs6DXFLdsaQkVKruqZLfBjP7O6k1rWxk9LHKjIA
y+Oj2/j3FYDJ9ut4UqYv0La+pD2YCORuqOhHJRhK01jREipI/Tf1lfrsFFSVuWoD2fumEBtX9vu1
rKg5/wYDc0Fv9MDNiU211Yg3P/Yq/UX5dt8axU/y3NF7C62HeyVIvB20IvdwhbIIgGT9PFpW627/
vEf/E70ckF4yyREizEjEJpDy8Z274lvfirnMMpXbPgOagEu5Xvlw4nQ4seyp4OS95lj2SUft65IL
7+mEcBVjKiy/WJMryuRFjq4zGtuvCF8Nvf0Vu1kHJ+5xh9QLSMtsnipERFLW3KbOvhic6/FPPbbA
ZD6bjKC95d1KLIraB+LmnO98zjvO3n5iLMCNaW+tPhWI1mifFKFIbLNa1jvaIMtCh8QRh9N0HRZx
ef3elmPilq2qmSW7eqAHumZfxqEs0JeCe/wSh1Gvb9g8Fzdp1T3XW9SyMLxqEsNLSLFSD2jwflG/
Yz32zwRO77EhxRD4A6QfNH6hHa4FwUoRbWdgS7l+6u32QWaVhUNLYkKo2a8fwp4RwNqzCX97LxYH
gGNsBA66AdEigf0IhmWK+m5TSCT7KA7/GvEYRPXKGjARDWr5w4CA1c97L4QYbCu5uSQFi20r5wa1
EBxA13mfdtC63MkgBRYhqsfnu66OCSHtEjOFzQESx9Tuak6Nsv9WzXiLCRhNt8KrllGF44pcWaKa
qhUR1TfX5M+7o+4pVHvSxoq6ICdFg5c9L7EL5ZrA037kgz2HV/x7IV+GLiBafIxkPty4owCeuMnS
4bNYemim1MwTGKJxFtNKlKv5wUDYvVzRh0HEPZSvUhyXfDWMKrSt44fdRjQRfkCXEodulg+y4o25
wcc0LI3Rc8E2lZ76TmSrnwm6ltFX4XGFlnYlX0I4m+0+gqC82gQBdu85ryDKf+Pm2jGbE8kbjnjf
CwMYn/7Zz3wFqu3v04FN8X7spMg34tpc0sE1+c7lic2Dc743fpzhnRBNpbYvuyTuRVxGuWobX+/g
xdTqDEeFZTJHxY34FWh5hLp5TB0VeXXsw+WPxgeMNUrS6ghJ3sugf2356ZVz1UQX22Bl03nUY2mt
rO7nN6/7sYz/ndMa/AfiybGZuiQAM4fBd1KGIZEKfNvkDNHCRmTL3EoINeSzMuSVsVgybOicqS/u
L4hmfAiIQZaOT6OL7ca+g1xcZbBqvG1nyEbbYuYRB7+Rodn0KRv3Aed767nrjKPDaN9JOfjoRfD6
nrgiR8I9Ka5pDvimoqlAGvYVdNL7/qna6kqFKIObYUhlFS5WxJ4EEyeVnGH3PUtU1b9Q/VM6TTVA
2eATHxMIKk9lVC/isqSBYScw4e86hMUKoopuw5DRBj7KXXDAQzgL6kz1+8E9j7nbrOcSSG6Kf+WV
faesXR5QpOzo6zOmfOp7wzK42nlTaddk3oY5qrMEH5QSB0JZ19YtrMBamouDVtBUHd1HnpoY5wgm
pnir8WggohOAV4QfJaCSBQcYOoIs2ajFAI1pst6cR2luX4WPbeSRnokMMG1LzcgHLMPdJEp5Emvw
n/8wvAce3fqoQaTc2l9V15/2rtPUnCvdGO5fMKEg9tRkJ2BI2Er6f4A67X1CwMbYFhWV9tQ0MCfm
aw0C4hYX2Om6LRBjAxcpgXU3An1n19AtonCxYQWVrWP25UGNhAsEPPdIR8iNS4lM1puiHC/X29o/
LLjMeXR4Ngv2wQOEYNOaEDWd6FYo1mcwjTGJy4DVwpTqQLL2Gm22wZn4kayWU9Ld2dWkcHoEgaWE
xoyn4SKrzGfFzU5v40PhP3jr5B7NbZRKW0iigbSMBeArEnlIpP27D8b/AWgZ6awGorCGs5NHjfrH
9vrJ5VIWhp/VSNpWj3s3olPBbHEaE4BLgil9DSV4p0LjGnCKhxQSE8UsCND4JEBW2gQ2j8ovS9nG
e0EKOrelbbSwBN9vp5NU3xbMipz7/tPV3wnTm1szX2mHAY35HY8PDj3YS9H5EHvPDyic1fvMcrai
kI2lg43AsPgqi3VqDZ5jCLqYXqC1aVzYoHCy2FoozFZKlno/1hTja6/vQQm2aV+GsqXB1NzOE6pF
RyeyJtYXR64GjxXOL8NSnRNLaz3KTr3RMMjHDhuUzc9SZNkEbvBsGugMvT3If+sqOIrI8bZM5EPV
BqRkXp2vTnpO9zBvjZpoUx9W3hjEr1ohm5PLTrWCiecMQlkpyIHImA93i9J51aej+XpkhX33CU4C
g56+T7Nu6xeLJOSIBLt6Fh2J7SrmCU2KJg5McQ2dtR5iVJo/9Lb1kozoN/dTlvPL/L3IdPJ5Pz1T
mHf/4kEjWd7Fre6f8l2Wns5SNOCx9OpsQrJ1cFNLEW4dzG9fq7hH4xlW4NSa6UMOK2nB7Xc/dp9f
xpCPEqBo0iSXNauoR+5mNb44eSEwhlzHherKNlYMqimvAfCdJITBGcUk1ovYrovwvBpLepHn5olW
vP5U32/o4RKuKeJEKxziX0PrzG30UYoBAomc+LxQxTlZn14zcpKvHgasyuS3Bwm+r773zWZE6Ueh
SMKT5W+qOaa5e/l7mbfI6xpcE2w8wmgP5N+rVtGTAjFfInrNeBEAWcwyZMMEydQvsjgsKEfM7Bky
I64LR6Qdpf7SHW4fsiMq4Oh+9lf2m2Opibquv4+OY8Us4WZJ57ZyfWu1JrNOustIbfXesl+pz+Pd
kbKQSz5jWk384u/160arArcioZ1hZlgglgse33JJ9A8sf88GyIvUAwr9dGzupoH28jaUMyYO2/0S
qyUwkroaH+h48UAZQRnfwg23i3lr+nl/aic33gHwYufdGB8a8jhi9mltZ+6iB+nsc87e7h6EcpjL
3EkKHozkqBTDyYjPGUocw23vTQksT6oAepQXDIbUoVxBaOnACFBfw4CjCXesIWd59On5bG6wqmY1
z6SutDYa8Igd9+TZhYI3VTIFo5L3GMmtAtYmTXcjgrpmntKZqSTehJzP7epppYpUcQ3EL0p5aE1M
OHZNgbgHJQlISLWkNVs/Od4x3RWVxVkU02wSCz31z3ljIFebc1lyHX0Pz6GZ1lTT0NyEqTY//L49
7hcUA7qACzieNxbT2m5InoR9Bn6JThHmJJFUdf+/5hqkuEMiZae1JKK4jMYvg8ohBj7iU5GKY659
gLJwBZSqw8TLpOmQfuOESkvSLD1FihIZ5b6Rx/tlq6jQpyBErDcwpwYCp56v1lkUWm16cvV2yoH+
6JbfsV5sM4ph5bxBsF3KIgSZTzEiHkGfAR3spv4F+xykPO2sKVz54wKe2V9rfR2+4V3Go02BQIEn
19FO7rgmkZXGDcW9wQeRgsOtXVY+i4/hGdCaA4xkwyxoJgJH9KiUSZp+9nxW2n45f6knkKdPqpz6
2ihTqeUTmsCaN7xoLaEUg4nERwdyEvcA1f5RRdQMIuDuZsFI5rxurEUakaSQ2JC0ULqRQrRwLPS9
44JY/979GH7M/57w8fzuFUspp5eDC5vlWpkToFDtL7TZWhnRy1E1CtfemZXBAjoYsvT1LuB4ZI3r
Mrgigaqh3/CfhlV6dkbKJCTQfyKQZkDOiIylf6Mr5/f5bYLPIDB7CpudusPcgffMWVFZraC/ghyV
g54IWnyEOEBFBQoPfxAQ4nWsj59arbw6QUJP6xiUF5BbS0+pje+OHXywBgDl73/aDnDSjYwsKCP+
R3oET289pj9BbDi4VdW6jkA90DM8KJxWT74qSRRYpUE4IxZuAJ9K+QwdkHR0J2iRrew9Mvpjw+wa
hk3AsR9ZYcRFsyvwaD/qrDIk2sz0gcLAh2lGacPvLPrKMp/HJYn5NpDfXD42T12O2GO3Y1dwhotA
3KO8ChtvvuHwTO4G1gyG+jos40V48nVDNEizOxxJ0UDgoPZw5E+OlzQxcGbUSa8bYy6mgDFOiS0U
PXEopJo/bGYABoQyj93KI2GsW3EJhbTcNzIQZwfXgm5KhCQi7S/iQi3Xbkxt4ZIuidK+tUiADjKN
FpZooRJbXfIpRYbJhANu1SmDOq5Lq305DPybxE3UaRckS/WxJTR/8uPFbIgv+bCPHaWPgkcSh9Ig
IjQgXGfeLSa6jq2G21BLIB0WyezLnvxeVuxOQ4qib80kWuCYVSrVMYkfZ3lKh2bD892k1e6euMfe
inUM5Sd9i14tPwFhplelmt7RsBbmLIP5lkmbUCynphIjsqqJIJJjYLt2fLqnaHz0dff+p7K/xBLa
6hDBt1loxL25RIpQbWc4s8nIyzyXvLEzFiZx+1ATMaZEsOP8rVg6aO8D6jHQQTYWi8hBwgQ28BVF
I7sUF3wUE9cZlkS2a9sQC/NOtgsMMEdr03LwgEPy9WUjKvQaX5hXU74Bma26aZUtmGPQgJJhwElw
+ces2w6sPo8JlsH7C7XFpXsQLM51/SDk1xhNxsUuEkNP1u+CbdiMPLi38hgTAu0VavzdseLYRL/P
WZ51npxLmSdq7NJ/ZazTA9h9pQM+iFLahtSGgiO5x7FmeBS03sQTKNNYtYaiZDjMht2PKI03iQ8k
csrZ3agATH9ATJGmufIOY5+9w4LieRsqSi782gt3xT/FpGJ6dWgIksz/guTjd9d2WjPKDmj93XrT
wzJijpmDwqgHhAsK1OxMH65PuM/yZ+q1djo2jMsSxNmqKm/+kIc3qol3aaPot3y5SkaPb8yB0chh
Kxay1ZcZQwOYH9VHehVLUExBYcHv8uBVAdEYPKIB40/flF6cZ6I/7HDFUbNYyBfGCtpb5EOSJ8AI
+HDWzlsH4v8bdyvb183Hx03H6dQYB080434nkzj0Gz6vJg/cV2g06yEARy3c0Fc+dwmjwld+C8C0
869pQP3GFGtlx5BQI2GrtSDKBk0bR0uTQ2ir0MNBt2jVOdNSveoyzkehlGLIaw/o4hpxX+qf4Gfi
u4mkt0nFpleOIP8xhUNPfKDqKy+a0DtmOGFcMw4/QE7Mj7srmdqNy+OjqWMmhMHFWhKjmSkuzBVv
kmEkT+HkmJPVcrVjxuFb/ya7U+ihCVQZUuszOY17uzc9Lov2ryRRc22DUx5G7PyQACbpAIXzeh8g
BZU4sclr0u1OxcK6AclIeBugfTtjdOOQb/CsdXKaayjytty0T0o7aTH8ui5oSyA3QSVFGIoBLKWL
VZ2lomyE3h2Y3pglr375+D2bgokrrsIxosQj8tKJmtJtXPs0BFPT4CiVCUuQB3gHmodkJHX/HB9o
DEB/yyEDYmjIIwBx/xgofrtnkvir5LqxANFfnpmpgjQ7cGwEiEgoaRnmf7/0ScSnAIChxcA5BfsU
DFIwPlQy6DksxXjmggwnU+P3fCUwE0mXSEAoYZXK97cAcDdJO0zxXl4sRqLL7z5VgsUWb26UsCex
Mh4jP3urvZ8daIZbd81uheEeApBQdcWCjpF3EO8fLzJAUy0jNOmY6ZxSZLO37HEcneS77YzOpeJT
4ncHXjaR2/mQ+h/Fh1ICd3GAg3yq0UC25wnDwM9cZfoniARZZd7DZELciXG5spQaHoyGyc1kD0sh
dqn22yL0q1yas0t7lUBgEvWeT7yUEPjAo5XNz+gARcNOoLe/P+Tw6Wq6JofjesMPjDM8dO7jZ6R+
Ck01m0o08Hm/iQEDa9A4JK2xYtJKzvMTHm09KUeEWPNLys9dG/glAYnZQFV67wfMRBDFF/9/7gKe
YmvcE5WyZWjOlDlpGlu944q9dlpEPSMs5K+3Cj0N/GOmyahTEwV44g7c4zVZUnu5ogVvh2K9oG5I
3lA0YVUTmiqX/zEX24e29iCPvDQjvL6ID7tlExQqLc+lnxD18NcWnJ2N2tEtiHSWkqcTrlCA7Rca
kWlY4Ia7UrTbKobIVD6EuVD29SW44BY5pnmh3RHbG3NT8VmiDOGAoMiRuV0j1zWdOHGjSzzjzz+l
OmEAl8rPbOmRBxrYpt9K3fBthr4nXeO+FLE19oB6rsI3/0sg8RqP7tz+F5y1UwinuLIhybGOMcuC
9JSdi66lzrM01tnhwPiniZqIB+RzRRGIyCUFMITG+3Fvb0gyLjOtaXT09kQmbhsS+CH6wfQ9rJ24
Q3hC8Tvh+Htr2PepElT8dM6dEdq3o3Q6/lOExASlGs7LfTRUAzei0eyU7eVTQcwyNU8wmhnoUWnD
TO0DwW9rVyI2vTZ0srs/ArRcD7ZuVcweaWUMM1aXhroI7SKpzSnUAsTTONE2xICULdwNOZRcDd27
UIdCLX9mTBFrEQt0addzkzw9BwnZ50GncDAg5aqBo2bSFrDALt8NhJvOWCAR2+pTqNw53QLpnxzF
vcxoMpgzA3lF/z1fabewo80wMztRb7bccgmqfjyQoCkqUey8sJetWzmU41QUtc+mxUMaPA/BzapN
z3xtLRr1/I39ML3Kvg1c/4NSRK4ov7Ud9feSDGn7+GEJhjtJu3NKhKtgrcOELE+umzLvEJV+JPdl
NSboX6CPOE0d13SzR54ldzle4CCByT7Jy0qEf7Eg/e5oeKryfgjdDA2lyVtPYceudT4v5qVtBxDg
TjnofjFNBWAvJ3/rNw9lX3MVFMSRGkWfUGIF2BWjBYUhUDzTdC9LDb8plfO8HqxXQa2quXGe0SQZ
tjYCLZbr8dw1Z5UlBe5LmqZ+RXZs9rbmJ1N7tFYljRiaZ2R2O7l9/czPnzRyGsYzKMcobJ+ORmY9
Zc9btStTZQ1aVljAMpvwhUcCjY84oPks8vDQBA1ALL5zmg5gYLVB4Hm3TKa5kgxa1TwjScjFyVp6
53E+c0JV0T79zIvhMK073CODj8H+FShYaIuW0WradPiwLiyI1WGvcECXtnJxExrnG/IurRSqiBNh
AIA2sLP85cX4dzlFVrpEoLsqhWzHCdkaQmWgoxnOZdKrqYZATWuY3PHydZ6II9ZD2eUYpps1eSF0
zVcnWMWQY0utmuyV30ebc/qmhYI33xQAnhnzSZJ+WnSRdT/8UPkxVaPxdrkPawv7JB6YHGNsrsKd
C0HxT6cdJBbZZ5NgDI3U7HJu2oCyBvYUA1uyFUL8YEE62ipHZ7ud2yOx7wP+wDzTzd8OcHkS95HZ
2BXfgYbGfS9/jfgVCooJKdLa2mtmOW2OlEDHAgCgwRnu+aOPx3aizFsz34p0GsIBej2ov18v78jC
zA1hgGAJ22rvYfIZ4hgcIcSbD2eIZCwK4hjSTqVaWrQQhWr4eYjLjNcnLhswL2XQPOW6nWbFNnqH
kHB93XIIYl+h87lKbBXoiHBO1q83a6b7UPyLFvFN0zb0X74hjaN/DC+XjYzEGF7vC7dygdV2CS8b
yaXh0HRS1X/tSJZswL8j3nVZnxtUULmyL9AqcziqEKsW/agwIzS7F2x/dGyAFxqz6yVujaehNDAm
mrByk/XeL39eAnALteB+rKFp5BFaptv/9U49vC/dgmPdCGoNzYnc9S9mGEX+PapS4vzPIgepHLDm
U5HQaA815MYCJaIyqztcANnaqQkQuvyDabpjvxXwGrB2xJ1gH6pN9B7ndJp+I5meVf5AJjW9yBWZ
ZiFmkXzT2lsepcpfq8G3fe5Yd3gAPb+BryqTR8IfGvJu/+IOIx5bVztGQ/fMSN/1ZNKNVBK615VA
aWAsZtM5crp5UoqYwDrcWedBZpTmj0ArXuYaTbsf9JS5QlYTLNnpHT+IaoP/7+0JLDXFRK/z54Kf
R+uYoRQsxjYseD5W5wie/2eOCS+areoTkWyuDAgOwvib6pgEJIZNyGBO54etLH/4Hc18FZXjDE75
OcvvvSC641Vu/MqL7Os8N6wcNJWqGA9Ytp8y+RacwrFpZxU1tM1P6hCcFqnrk2ekqTo7AyrQnpjy
L3+m/ee8F9hwLMXpGGnyIWkiUFJF2wszpvpk8NEim6DaJay5xCbNhK/HNAapfdBhz2WBxdNkLfGP
xAV2srzx2qrZGGBzQe8/3U6+ZNmnqehOt3la7BMXYHlqKinEgf+ohJ0vxS2oc/y57qihcBf5ITNn
AKNkMMlrjWF73ufGFvnhQPQGiJP015gCUFGz1D1uOJVP93901uB2yGH8GpIPkxn5IwoSm8OAO6Ey
6NG2rKT8FihSl7Qd0omv77CRbRnK+2skmEVKwl9dLYzycZ71jDNE06fmfEIR4wnA8RQ1c4ZvktW/
3+HpjSgrTsDVNXCUldoWyEF3/eEWNr/msoe8/WJ/8YwPHsf6ABlsZZC+jZAqp9ykenh8Xr009E9y
UmcYhOXzF9fbzMDZcJLQHvqYRMZW+a1IMpcjgP6wzHjs4QWEfaMWsGARVxZxrFkEP9lPiikMwg4Z
270mEY0D6Viqlgi76IG5O//QkHUpBiA1+rtqi1WzXpQtgoqZtlzgbwJ0PVfA0boGbUXOrQ9bszjF
tBkel6NmkYCdV8Zb7RSAXoAnSiayZhzPNjg/ti+Je/gFn5rsSUDhU5AsZmeDW5dj0IcihhIsvHCu
lSS8dC39K/lkZCfyw10zZJqhZ3EOdKuSlIeIP4/45nu8cabEKOHfd08hFumB3NPit7CKoZJQq0ko
nS+pFan6Y+MINJ29HhGdXRbQEo64Auyop9jt4OjIlZ8ZROC3xjfKEwAvXg3sHnt6E9diFh6hJX/A
WKGVIb2TTVJY0Xuf9VGq1PKoYA5OgWrbkKIwSEYiJRe9u6xt/hjhxlFPvmMsTQYXyMMhh0Zd8lAQ
tdBLsZDGVJw7PX7y3JMGQ0MxU3KGx5DFePY94FN6QOyCY4iVKkmApSc9ZQclcNXyeBsUXREU9EL6
pCZz8miPuMvrjN7PHpwX0h0YMC47jEvTBLOdff5yKgr4xBfwoTgb1zqcOHKOPCZNBvSRpd7n2V0I
QTrpXecHK9F20cS1R5RTramgv1cmy7HNn8JOamj1VWgS1ZRHoIlGMiZnHV+5Iiwi+qjwAm7WlHdx
bFljsRBwHOljCjUDV574sDf7VAsAgNIpJvC+ixe5yjL9PvnnG+vz6jgp6Krlb++WHaUX7m+VAK0K
weGz5W7J6VMaPlo3UhPaarhn4qRcnMhjUtLVZ3uFp1WjNGzSMgylmV2GIwX0VN1vuQxYZpoT2C4U
bqWaEsaD9DdpEaFIIblsUK07di8POJYjQ4UZXqu1rW/Q1FCasgnbBkj3lcDzFZCy5wGd/CJRSdO6
GSMADmUlLaB1nGX7AjAk8LZltwwSzxU+fzS9C4SVJH4Yephx/wYJCra9vWILVelZKdUFb205si9i
vtnfPRkROS46qzeQUwVeWuIA0+GF8IIhyli0Onsu9xcRfFGiHljYQb9rN1NxUbzk9+A1Q2pHjNiR
35xY9TFgwOUvnZpqaTyTsErkGI+Ht4uretDpJW+z6IMYG1gF2QRULFS4vkIuiguXtu2TNkjm5xMq
46dPUYxZl1P/gl1ULrzn9PTGduassyLP2/K3VmBRHgd6Pxt6gmRD5Kx4a3X3YL9386LGubTMCx5D
/FY5XUYL68jd2e5x+LNBBM/WoW1+P/3T1mYKYR0kLQQ3K4rmJdmO0ORXgEG+0fnmsxxGDgwewmwR
X9dOJcBDJ9VQ/uBuWkZfo4WoMMMgN4kdHNniEL2nYAwsMnzeV/8DedjOtoH7JQzZXPK42z108WJl
hR4qTjpnYev/RA+BWnONTG4QfhxUcRjc0YKTOX0zJ6eIoEpmU0u1C2XaDJYXWhrtZk7QaEG+ANwS
FPFgf0QeKiGNY+w7hMB7Yjss9N9Y9FJjF9YVKOa9c1ZbrJ5T8yAGH9rrd9WKxqtzaDsP3lIAvSsW
3EVxDsZympec6kxvCQ+j8vuXuUIssPQGtntSohCM7vIBKqWN2udobC3GWI6CnyRTknHLgZ/egYTx
ysKQ/FjqLejrvVFA34sKc3L8ea3Y7lb4m/69ON0+ZFjOL2nHfDl5vJ1uyPdB2z2Du4mDgS+WxRGa
sF86HhV1Mn5KV3G+8mso9uF/+OV4MuDLEgJTw1b/6bwShsaa+l9aymkVA5+WrgsGQ9TzLlhXRS4G
jcRWFtWYepCzig7f5R1nJWZAelngzN5QUDJAzeiO1QOjPVvYyj2S+TVRdwNU0f9pwJakcM6chCMt
XtKLjMrJQ3Hl21X8ZkD6+7Zjcd+carQNE8K9SWSRXRsT1xpwy5JQ3kiWweXsTgN9KnlQlBinOE2e
Q+ceDd+dns+QkGb4JaoYfF+ngQmC6tUJW0H5oHEzZXVWc+sgY6+5XlmX/KESRu+gK3hmATmOvgjF
yMPcQDLbHSwtosov9/v+oVNnQArwAuRMEWLiAewoGt4LQV8G7fCtErmH/jXEjbwkYsC/lSIEuPnH
47e+bZj5uslrac9roNvEX3Hn6ecB4plEjA6W3kElh3s0zT8m0wwCOOevGs7xj6DQLQsIksek2np7
OppwEXnlLzzUjGllN9w7SP2eCehVKCDZ7OFCXUf/WnewDDvNzzddekuSppnDJtrZM9CANda+hNrW
50RO+j+KKZMfdwPh87/ItdjCkXKmE0lCsNzxNst/uMj+VOLjDA1kSoy7d/M2vQoGD+c3I0ZOPqXi
7mCsPGFPuyq1zsKNuN8ptod9Js4n56lm+Ud8l7gf74qgRqxrYubuRWGwkaTTjgHdbYbGJi164u+3
MfLKV0QO6oNu2Lx498mJQ6kUN5ObNykV5Rfmy+kuzAmBezc9rTWg7BT92uRfhRbeWDpRdonycK9M
fuijBXm1GDfJzY0cV1ygVVZvwebKukYKtDgrNn8p9mPRrkc1yNCGrjg9Jcj3b2FAPFl9rOpAlTPA
0GTfnJ2+9oWg5hb3yoW6PxEDnW6uamN0mNQKFIVYZQic3oAb4LkX4343m1w0Ilz46QUj2olnAzjS
rmHj0LqbM/Qr8rB7gKIvDXQ8PKef+xbgI0GZbDrHJtRYlJ0B5HaDNPiATumkiHx0A1v8x7yOZ0mZ
DDmne/rzFKS8PQgdCWDd/hcZcCLs5EtN77nkEihZyx0dEru0z/0s+zG79S3Ay3MjIZBXUb2qqDiB
M5C6F46IJXIEovMIRYu6+IoPTWe1SWDezECRiYTDfqgJ0U5SnRoFNQTOfjs4igSXXl3+hBdUXxg7
K3dfqBqe8f17gZL2fM18FhWgWIqkMD4xpa4Zp7b9bf6cW4uaIkcNhdAULzks7VK22NUSM+F03JaU
5LyeP1Cg4DxnA/jjHSO1gytRUcVCSFDCdv7JhDnyPj3wjLVU46y6Dji4ONSVHWZCrQ0EascbZTPt
TaIt1fWPwo7Qy1qmjxh8eSxYKzLdUdOcQw1EEG2O5VTwSaK0cgnIHzsuAoGzn2CWuJLiKl9OkgiQ
cl+QqnaZ69/6sWPdAbx1fS+1Y4VPvG9lvVCn/h3B9QkEu17K3DF+/TOuG/2kvzuj0TkNuXulSOGA
NhsuFN1oXL0aBKGfPllAZS2ug0g7SBRVNev97h9KirNXCoUI6FZ16O5fkQfEWf3bi6upYhata9HC
Y2NkqgNyhGZo4QxoPH5POqEHOjAinRsunTpmFLu1GK/XaSuBAgHlbiAUwli5TsLDaXc4DzklkmXh
MQfysh8nzdR6H1tPHOe+vop/IDJJttqAoHIC8Cn7v8KOnrheGMV3o06VJ949y+g+vl774e/+d62E
jS+heaT4vD5HBREjVC0XsVFHoNVUil9u7+CqnqBoRgk6VSYTQ9Tu33BpQ1wxXaBtRSTl73nusJb8
ZIpOdSnsh3IAu7i/iX03sRiTBZXmulWDGIMSKRUgskzFIViIVaGKh0oV0WLpTwTjwycQsjOZo0+4
ftHrY+EzxF0Q4bRKBiodX1B5mZopO1018hZUk+uo+98b7WS5bFFtDULV4OFQ52YUNgZMRtvEoau2
8iFH5MTBcfYQgwhbgmbGipzUX0dAWH3Prtk6W1H8q84c8wknbF6W4q0ep+/hxL40Ml2lQIza6U9y
7jUnqJuknHbGexvnNR8iNLVN+Q1dDicVcBFgGzgXxLdH0YMcSxy1DGF/V5NONTu3SBYBr7eAFckr
YWc3Vb1U1MuDM6qCGJu94rsgKntKQVzSupj8fezqLjCYeLvrUmVWmAYOZJi2ASbNlEEGp3KKmDYS
M+gJdKZPddI5NE3xNoc6N4Y+2ECUiLeMMKZ4e5WUh+ZtqV/ZeeIjjTIsHOd/TydmBWTzPl2W92p0
MrV96ndMRoa9KojWGs9OhQZ+I2JnitPxMjqgeYxczP1T5/WN15ULJtDx0EM3+dUQNcwcedPTzVFP
sPfdMkVm+UlWLtyfW6pp0KWRnwZsEwEexA/fsQzRzfkN+VZ+ivWbkOa2PxUxtLi5QuDwfOnaa28b
lgRPK9nlOMrxeLg7ny5cX8sZVsSl2xhFX6NJUx8Ed6varOTfwXhclVByD1Ipq+c8U0Hkb6rGCgv9
g6HLxZP2R7Lgv3STnqdPNMZyXIJKpo6ihTOUclENF/jzlQBS6b2lBTd0Y5g71BMl4b4tMAfzxwQl
U+yGRG7WOrC9Uo2ZeeBv2tW62rW8LcOqUsZzaarqgYJlBpn9ZlMccOpxgp6WQtYTjCnGqtW9DPPg
EnAxXxzuuejUUmvEGVrBVbkQLhTu4VAzS4PES2yqaLOJHKWWm4mf8M1FeNdtHf9vm6gtwbWUX0xJ
dfL5n6UFw8hvSler0TwHtmSyVrK/HzKErjHuAmfXX20RxA/aOsx0U90WHWjkTbmSycZqiHNMOi3S
UUS410v3BJ5QGhM4gggt6aXYyesJQfNkmtzOBm9pOKOzn8OypuVZHXXoDiOmi5sJbCV+m0w3r5PU
Sj6wcfLfivCPN+iMGmy3U0EkK+3F2jWeCdV3Qj3U/gLj4heL9+rcUmKmlET1nGA3iWL6JwUD27D/
JZdMvq5SGjmrwgQ0qnFDr7Mc/+m4Yh1+8Ft9ItMf/Piat7+X83sOIP4xGQ9uSgsuD0GdTbZJUbcJ
MRjf/ualkfS+p9oo6dn2umEX2SOdADWQL+uYleiwhf0QSx7frK5mCgC1Ko2pjgixA+2YnS8pOmZt
j7g7nvvCWUGaoMlgryxJ7JLQSE7qDxA/iKReP89jDe6UQi/13sA3t6Q1SUF5LC4RHag6ZdiyHZa2
mruioPYjb1vQsMueaG2haBiTAZblK3sT8iI9J/Ys84WfS9QTiFsCEN4ztLv5Tz99dsDO++iAnNJb
biB1LQsoWdHBp1lNR2UN80XWFTQwCzjpkef160uBghKBb8vHxwpvQvAalXvibOxhjiO8Xt5pbTqc
ozWrK7AsAQF/L+CFNQGTHJ3lG+WDCka4KtmBgsaz1H1hnfucMjyeE3dBT6kZQNu0BxyUPvtRmvnL
WdmIXwhkDRx6ub0+BANuwXoc60LMex6Yxq1zb8TwIlC+LIWlY5a81CBFuPAWuqdpFfGdehdLj6QA
mlnpakSWJc4XWSvC2Tw4u4cmoQ0wjqm9s3lj9L5owuuRfucrIQKakewrILEK6GWDxgg22g1DKAcJ
bBBYmQr/ZuPFAakCny1O5W6i2v5H7kTqi+dV8Rgv28VFKbdm5T7l31YokyqdEwE71VP1cCyzhB4U
jW0JNCVQKa+fZ9G40SVXBt9lVyEShnEUYnbRc8Mb13vXYZMn7m2tyNOkSLoRvhgm6V1qh/FXsTCt
F7Pp1+JRaB9obfA/tWo7IdOk5+bCco4vaJ1I4sYM1oYRqGOHt7laV/beC1Z34eRi/gnYKOBRZQHI
qYz6ncthU3IWRP7jHKd6nQsYzc9+42MGwB6UHXW4aGG+YSOCQ3ZBoO4qKFc0GEXk6pXhQz+4lAql
mZ6mXuwn92ivNGniLRDaPxurE9IC6/MuNZOT4kvK3NPrnj2jSpUhJADXVSJmstnLX3p++d0HrlRA
L2D40JXDnaIi3XxrKD19DVXp8mnCr+0tdpLNYg7RZJQQmeb4eVbljQXqHuxmxnPCVTy3Yeu4I4Eq
etf6Z/im/+YmoDIyOhL/2jFQzUB+fdddcRewmW+x5Q6Tf0IX6CAcmqSanxySwWWScColbmg5wFW6
PYQL/CmC0FTHpqmg1g922v1kFraeI/Mdf03sSsjXBkv3JBLnF0az05v+gTGZA/oXtRndfFUMaWbF
JIOv16mdAEVRj0UOFowZyybha1+8Kf7VTd2SqS+KI1NgGTuSWqnrDDjGdx6icU+Nn2LKVakX6Cai
lJ4nwZTZDAnHbijYWfSqc6tHmPUcrYgf8wtOoAL5pHLthz1jTm14vP1OOLEXtxwWZfB3Atks5mBo
vrplNjLfWSnwFuQxhSbVLoS1LMskDPOZmdygTn/1C1AalJXL+i/20PCHsoNxMkAaZlBscVhVA32k
epUN9iMy+GBx9EBzMBUzg8Qc8dpvFTbT+uhjJEd+6d/usNqj/5rLvIOOJ+MkSgf2x3+430loBxUI
LYc9zKZPhCNYIBmnjdJbry042ZFf9VeFYDttiCVzcKKiaJu/7HKwoRbppGQHaeUk2btl1PbTls9P
Qlq/72rMor9sKcL5PxR4ZRe2TZepkPMt5VzDAd4/RVZdCrc3sixBvbVV6utwSjKlvtigeyTfaIMY
ExwU8zXTlGMj9Ppt4EeYG0Zuo4no8gwoBhRUuvTv2c6urT4z76Or2IhwG4ZtjnDXODBm02iqQfeQ
tRnnzTa2HGN/eNNnSr5wr2n+X2v6UQ80uGmFc9Uz5YN2pRooySly8NDuFX+DSLtE67gbW8CNTGMA
CIesH8nbqqlRuRyR3dstMPcP8OHIoxC/bckUNN41AKwpQJ5Ab39RyAWYVsRGFPgXbqd7HPwRhLf+
alLsF8WWMxO3i5uSuGeMRlH6WmZce/PtqMUEbXr+sDkt7D18p+vk8k9D9h3v+lfpaK7Txd4T5Ab/
1jp7zIZ41quQcw4L3j5uKAP9mzHKLcDVi2EiVtqwDfM1IX0lYTYAc1/BRW7N626NEIMQ9KDvB43u
N4pSHQ/z412vELABCBGNmJFEmmTGBuz64LfNj5vBPmQFil0mF6hW9MaMCL0p/bAXNk5S+s9SDVnq
rHIEH0pMpYDixinwvjDwMA8JmwRDMQ6dw33r+WU2mvON1WqbzW/q9DKdsTuoNM76PZGBEVjg0gxJ
FmZ5D/DkMTs3s7tMu7uxS4NUMzdIfu8bZg7SaFe1XERWwmQ0qlWwUOtmIhX1FI92lCdxBknjntfp
7RgmxYTy0hNSUtL4puEWotI1XPPzRG65tq/8f/TCByuY8DVkF/AbFre3TfXBDX3Ri11Pn26H93OS
DNGH5vQcKRLdOSyJ5KoX8Qpga7sy6hZAm1z682gWcvGAktjHo3BBzCSAPUKl8oukO7vOYne3kPhu
de9vDg9FOoEi7D5fanJVvqPuXGus8zKoEc/WyuZwEXHRlGnjCpJ16/5ju0ieRxC4tjNBn6fzQAO/
RQTRFONojJQnxl2aNSfRL4cCF9HDeAoI7plNmJtS3k098mDGv8s1R8RpSXtzHmIUZAVyW3Cla/9F
68wKeCqKwikjMyL/q5HC0Bk9GWUwHt3VVnEanATCvz/gVVqkW1TS0Xyqb9RjToOerHdONH8CFZHB
QEiXO7C27I6sV2UZW1HiXG/bXt1f6aHnPvKWUyCK8wuwCV+O9c3XZSN3OJIFrytcIKC/kHzHxfMf
UJt3BwYqVxxe5rFcPLrf0mIFjTppdZG2uDhnNmz2kY0qylPdRMB4pFyv8AF41fZMtIsDdP3jsXNH
P8gCWjrY92e/9nB5A/66B3UHzPW/jTE6Uv/lVvNEkCqfYRCIPq7ScgtQz46Zy7uR7zcARjFcis/z
3HvRdjPcgsZJ8gecxkSKxyp/nZ5E8NHEE5+qLm7s204xxo/IhytFstQWnHFbGmu0HQaHM583A0Np
U5vXCQpsSa0nf76v7M02kk9DC2CpjKxT+EfLpy26L16+96GNX3L1VIrGNwGzc8Ug4pKTlxQO+fVz
WKYAfBGLNHVsZiaACDt0u6GEkbvFqWpaxmCDUERHaKigaJGD8hoIUsNfGkJKLmA9S79PhdPvX+CV
odYhcDlgBrHEi2lNpm+9/RQvZi9eAlnxQ9EqAfigwwzWQi+GPFYeYz24oO16hk64owfccReWSZe2
OzzQbAhhGNDGPK97yXlq/KuBzQ00e7ils6s7QGBtPx5mKOgVDboNbarKLmpYFgFNuzNFNZRcH1Bu
N12MyJW2CaDpXXGJid2JJ6b7fbs93OZj+xL7LlGGiMHkRogBLrDCe5IApq7nG1jHl0/VZCjlG07f
oPZMKSc2MVouUcUz2Pwe/BtxckThyynXwSAj3b56dHdwsoXwFeon2IdSB8VYKtqYogTz1pR9ylIN
GteZk3xoEAsO7cnVtXpmPZ2e//wWNqh/l7soauEDKvYQtscK+u7g60I2IPRovF/IyEKfkZuWL38E
GQebjpebsre7ixQvRpcRplthV31VBftzKXBnqsBy0wcnLcF9gAV3lzSQN0GWGiUac+MoNH+4DCRW
zVg2+QyGySfOU6Dmah1sGhbOunqzPsOYJTwmFASQVs+smwENsgn7LuBznxgaLyPNhG6fT1BThR79
otWT2/hzLQCIx67T55/fvI9xDXECCZl6aXXlPrFnjuQvKie0HEfWbCUMviS0b2k8rbc10IJ2ZWPN
xoUfH/3IhbZaI1PWn109lb5eg5AAaRSU0BMMI6Q1mpTB4KcnbVWt+N8lNmuLubjE+spQ4Jp5rLXi
O6KtzNwSlchlmvjro2HSe6DceAiZpvf1IpBOrDLKGdaRstCzlnE760cqdmMQtZ+vXo9qr/h865PS
ZuUOPI/Y0+BIEV63Nsn88/XdOCqMTVkIhaAmsln0dHXJbwECiWZp8UXvhTPN4D3rYJ4gNITrsw33
sqiil8GjmYaNX9TKYI7zpRA69zpdULuiZqIUfECyOZa9BwuKZyESBi0xadCTBfUzzBnduHvxbrCW
cR/i9lI2BnrxX2A/3UXG1lCGQ0KCWL6pHOa60ca79zIfbjRR8pTk42S/Z7M6IYA/co5LkxN22KHv
r1ndGg6x43pex4FI/umAeetfu4lII4afR7EcXzIxBQYpC1y8V4a/o1qDT/WU5P8rRHLlLaxBEXJ1
SyprHrsYvqz2rd+Fo1Ut6xqKSHACCK3t/WwW0uj8LqnsOjRrXH3frZe9wVclehYBAq7itig0JIua
zLmWLcaNMnafzFQ1LSTAOEDSVqse7pRSZjosDoDuk5DvaZiuHQnCUagxvlRJQvS13GFPYiAs4uAS
af9JAX1hswMOUBFv5bgkn2HRMd9cFzwiQlNIMuSuCopnSaDqbIvOh5vZr7nXToeK7SunpheX+XAW
iC55ipc2PIWP0yH2kDVvLzTVBssCQejatqqcjnF/ZRZspgrZ/Rxfpu25JUUoJZdB9Wdt9vssee9d
F8QCCCbQBivzBCRulvhLUJ5JZgRQ7xvttUOVzenBoWdS4tS9iQD8erriyjYUeBH4vA6rF0W3EbTN
7ivSm2WWKPTK4IdOPBnrlogjew77E2f7hQw9gI6K8xJzMWFVR77Gyxo5d+Ib+32jHl2Gz7JAw4hE
G9VdiFX3UCJljSxUWg0NIFN9nX58fy5hBmWeCk/Xt8kZugXkpiegGIOeNKD1AscpBxF2dIxmnP/p
xNPxBzepdf5zM76Z+ZQ1QUW4/HMMPvHknYQgdYalpKt93oxMqX0Jv3/BhYE1PQhC2R0HJTJF5PYQ
9lM91R475O1s+a1kIeJzuhGr++OuZSWubRg0m3AQIXXlboU5cwVV3LIOUgqjSXk04UOLs9QYwKb/
PSiiG8zrPyPkjjwwlubp+kBuAI+bXqGlOF8EpvscmloeBLRrblItRcCTCe33SiGG8t07STV2o8kk
n9AzAmysb12EQusaiZNS+REZAwXzgKF94mZuw/xPM1rYDhig3NawIaMl8ZmpH3hMp7sVOdSKPDYK
KEkvM2/XehW3tFYmIzY/NihCvPvt7fUcfxxQ1EJBzzdjw2gfqei08HMmgYbYj6IuZwUEBeCFTspU
2IQWFNxWmYMgbUcA5gsGwb6T1TGN2SUGgDtLnJKJt+Wm1ipuaF7n8DiLQySAHKONgwE0th7L4PK1
4FIsE/76Nlt8e5XD5mMNRG+xP5pcl/wWa6wLmEQFKl70y4yGudkEeFyKNnKkWv2jL9FeH2T+Qdw1
UjjcUO4/c/3K2j0JePO1ZbZNdbJ28c/xORSGoOoWqT7YuMi8txFNi41VtumXGz+1H6V5/OxaTYLg
rMzk7bxWZG9OCgdVsU/7cfiolUbx2FFYw4Qs2uW1LmlBqLR9vCgvS1YjIQ7iOpb0zG5zXh7cCI2N
MfdPvkUePBH0uq5RUihzm6zlEBUh+PwQO9aG7wqK7uB4fx9edmvdg0DweueDo+00SwTpzCQEH2U+
8ZzGtSpSwMg1p1RIyYK1Suq/ELyeBR8Sm7OnyfCjwhXD94dcjKY+67NaLwY7J5d8Na+VmafKO529
y4Roh3B3w7mgHxRR+2rRu4MPLgQBzwDeaDQ0KXWIcOQmK1dKdjp1aWN/i3aRtU2g+mlEcsl2bGSk
Iv74mUU2ckV/GpOMf3yp5vsRWChgZyTfsyfayhE16m4yUFxc8dkXDH3MbEfivBW25s6mhv2+vpr6
Yi5/ZksCPiyBsBLy4cxpO/3P8kSF0sXcAFx5Xr0lDTTwOd0N79wjqbbgE1NAUDNYmbRTxEIxCP3j
PH93a9ATXVO17RctB3QF0MLR6f22eYrxPflKhauGehR3nYFa+NmiGpR3HcVNR9Q0jv0YC/1diM4I
Tq1nB21XoTVo93FzT3OmpFPHX87WDGtR9JKmKbYTPEcD4VpzdRQ2x/zTMjCjrVdSZzZTmSMl1USC
q/mMSTgbenvKoawSneea7m+v90NsbZfENkHJm2zuo3iFmEbLstToXGUUV65pIo4dKB0fnjlkuVz5
Pr+254+yHG4LkSVvp/tHvJk7QUauhqkqxJ8O27qMy6fanNzqrN3nrtPnOUgVDPkgiRUF8lnM80g5
Hr0Sjj4TGdb2KtRRT9mhQcT0u08hSg+9yndqpZctsGnoP0Yar5YTMDk1/DA+x5AWJiAUJhdo2V0h
uSOJ81fUUqF8Xb5B06l5/k5qPwQDlgSy8C5X8kmav5zYlqywnqNxb8eKitEooRPicLrvi0/TSwij
Che4Qew9oVJcXqT2szwy7tSlJrcFnrLtlZm/cMIkEQRqjxPcdZZ5mY30j7+Q2p+8mq51Umh325V9
srpZ1I8ER/Hzbmdh22nbU81rTN8aagEFyYlPReozOD6eqFqhg9j8DlR05TCTdJHmSLBE2uS4cb1S
CDbuA1RIpQWV2X2CPN4MQErXRYgMeCBra4Ckk5c+A3mAo07ZcAu433yQQbPLVF+NJe6onk8TMF0K
U++L/AX6PG03Q3Qf26oDCZaEJuElkPhNOF2mfmbXxrp1ZQQ5IYkGJO7ZHK2FBoxXPqLSbmUNBJFk
UiAyniax5mKiiLB7KLkkPtNhrO0Ikld/3kEcikMaQzVlMeDr1jrH00id4SC5HvKYrizHTUQgE7pd
LVk2DBCd/eOFgidVTAIm2qy8RIBPdVay3D7muhxwBQZWnAakRFPdceYN0r14A0KuDxhczHn6KNZO
czeGCQohGTOt8dBhkyK8/b8U8/rqY1cNNXsyP6+Yk+wz1+RsMO2Ffh4dDFjl8ji/DrqQhsHzHcbN
RsW0AcFG0Vt0a0WkWFucPBz6j3oDJLDf8r4azucyMOnejp0KNEUjcdaGtf4hfqpc3Mm1T12p+ZKi
FEgYmLvd5IDdpeAwNNnTvqn6495vFCxu0sDl4QSMJMSs7p+fP/4C8UKQFmiybDSr/7w3fOy3kZ0S
/NVHNuG28qwM0QNplaMgDRwGTQsSPIO6Ca3T6J9WLrev2XZduMaO9uHN6wPYtZJQtzuC4h4Jljnf
lyugoNiwWweX74bj/eACE3UbUV6tpCZFHPt3ArVoUGJyDa58KGbO4S7fWF/bVJUIuB5+YxlO3Qjo
ZfmKapX3z9XCtP6b2iJAgmPVqPfcmCwrN6yUKwxFY1goM6dGAtIHmhqFIBXta8FoA73n+x1iGtcX
FpCUJwaO6m3TT1FpSr1R+EPUnA2JcnRkzLeHZJpDYi3shXNV4Scw3QaK2apDZzoDVSMLKFNeRvTJ
wtVsj0Licy30GNSTEZIuz9vdNWSdB00LmJ/JAGMtSZrgrPihVN7e9Pr3I/aljB2tSbrWL6ZL+hnQ
WvOFmHadgFzzA5J2oX1lyV1RS/1rrXhZA9msnCRYmc6kw6sXHu9muiRlX+ZpNUVwv6dcZjjJYa+N
jV/ZF5NEbs3WLq2iD91tVmaZPdpCE1fdhXpvbsEo6Dyu0EvPG0azfg0pUsvOxKVTl5HqGYSyG8nM
vw8WkXN/3h3r2z/rB41P6WQLKw7JFc4LuQO3utQ1fLY+j0XU+kacb8AfQnaDsntyZ0CO+vq+ZdEb
DiNl9rhfIhEN+orbGOhyY3YtKLh8R2mQPRbc4s7YDudLrbs/+CJvUaTZc/QsMBje82nV8COkMLYS
dt/kgUZNduxFdxNFzkyKy0ZEg7uqYlUiUHsyRlXZXlL3suqwtRqPOtw16rJe63tfX0x0X5X3AE4E
3av5KDXUX+g96y9L0qvcGDZr+ls/pvNdFHrNUpxzU8d3nGxx2XGRp+eR9+ODM/tS8NR6WTtwRWSN
Hte4+JUKHWk3PT1GOXK2tyvyS/h2uMj7g2NivXWrGZFAelUX5qDU/NLpiHFozGd6x6bdwmIETfCt
wf9XKlTzYB2xU7lIUUh5en6WBHuZlxbMH4XI108VX06o8PfZF8JPzp2NkyKXPx+aXJhx0xye/CBO
hSzawT/VzGc0aSxNUwv/mpmfY8a6cyii43vhb4lOqNxvLKxSkgmn8WDhHBDi/jHEXdei27EjMMhI
Wh3edMLTQqRWKIOnJpYtDj1fJqchN3ZGagHJNs8rWURKY1ryg5obT29OsB0WKMujNQFR+Mi8Ztgd
6GIP5gM6/fyKrIKT6stbDPlNY0CNv2XkzFqF983fAAKPqL45ek7u+CGtiBmkPvPjA2gclMxUdwtl
m2LJMz+gSKTpAgM1ZWJXbHR72+x9Sha9NDEd988soFkoRnnAUXBYih4Lw6WJEd8/H4O+c1oLTQ7D
M2yDLpJSAAcUmYNDBY7MTm8Z82ylIm7SnER1jp+pKA5Cd9tqe4N0kkr/fcELSRpmRhl2h92we7z4
Bhy9MKkuu/EProiBiOo9nU44DXKSbylyGFGzYWAPjrNmLmihM+xovEBFAVHi2pSe4VKKGgZJ5Bic
Xdnrp9SOL7kPteIGGiI58gvKph9CKzCRCkz8fq45ltzRDpSsRmgr1Za+t18XABmHb9i7EqqLxW8h
vtILsUu1tFMQYMigQ/xhwWlHvQPpuBYPxIx0HweVXs4ZVy/70QmBgqdniD1y3exDBgQO1JbqJ7G6
8pnV7HbMXEvDbblvnDOHU4UZDTSFY5c1ozM781XIfQ44Vc++FPzCBI6xEvtpzgZ+ewXKXIFpBcwh
79xXB75dVlsHbHkuJEVWmLn+sjvDvF2DG8SEYUk0//8hB3NpeQ+WSPZp5i1QLvorTWSyLsSMoyfb
LjA6CWpnK+nyincoVEokDkd7KaRpc8gfZzOP0mRIDMbDo/d9s0mvqcDJ5Y70tL09rF++iWbGGb0x
x3bVL9TPyo6gsm9dLTg/KGuMyeg/2HCMSrcMxw3aUq7qPi89Zm0jg1c+Z0XKQNYFvQmNU6IO40gl
p1GJDO/EU0dUSHMzrtv1V2vgw+gqJlDRMtDngC8Ts9bN0OJjOaTQEAu7pRebJPy7xmHJsWNuWh9h
Tci2IlMijCxJC6mNuwqGFFX/qeQ0yUjAL6e1tur/ljsMxKmZS+f9spNM+qYJJiBcVt0GbYjVUuYE
/Qj9USOveirkIujsE8Oh//FMLkWCegXowvMvBu+NSrYLf1RCvQTj0q+eVRJ/Ne8MeNr7wPH71Z9r
NTjZpSYxajCidl/TeDBdXfX8BdoOXHYgiXIgCoZDgUxF4Bal+zJp1BN9ToBWVXDihNNS7e/SQsTb
kLgp+3Ljtw8yDjDb1fYBZ/mreFeG2VbyjiAtpW7jwRxpfi0JNGiK53pXwG10gbnfLbDiMEyVZdcq
VsnWdEZHgeKBgvQ7wEj50RFKXJykJE0qRhyn52zNrhdb6RqE2sSl9vP2fPBFlwDjJZEVZqUqqARg
CRbaXexiAmXFBTD4qjfefjk6lUbs23zZeFbazmuvKoUyGq8C7lr/Btfth0P4oVPJF8NIVY0Altz8
8RJAFpdu34XK9H2/PqRi5YKyGTwUxW6E9xwdeLftJhcD3YcI1sudWDATGqXn9KBO14j98JJA3qFY
RzgtxtpKicqWtGSMwGnU6PZ7QFFfltkqrbMNiiFp45dLYnewVNPCYnP6uhZf6JuFSUbcQmEg/v0d
WPzDZ/Xo5rxLdEivBlzF1KZgIueuazzNLQcZmSWh8M0K7LyjCU94oET8jA9sYKq+bKsgdyWRLgjW
ed8iXAipQO/KFtiPKO3qh+DSuw+K2cs654QW5BHgAdwL8U35w5GlhpSSlQNGp2tDmjHpMbXcwt/8
nPC/YoKdu9Np3OAJEzg3PjiOqrVc7hgm8De8pEPOmmC0vZ0XakV1VnvnZ7WmSYhLejUekGjbdcfS
N4jnMOA2/ZD5ebJQpnK5cuWRFQNKoXpx8IcMti96K4aqTIdE5Memd5S697S6Pyr56czGidOy4WUV
IzfwOid9+FdyOZP3gclKPTlibPJoKNlGyGIkxxyimTHDm3WxUEFwUumBv+1spKZjrweH3pqi1Ntc
dN1GJVmwOTbJBNp5XDv7tv0r0PujRGw1KzfsJUBzuunr7I2L8BseZ0F/HzigWo1aQvKxqQ4kCPxN
Bggh2X0EMwsPQwE7Ui0Gx0cDx679H8fO55t26+jk1PBE/ndLUL+AHpRV3Ly1zIQI02UFcqbQbz97
2XABWWvGwXCRL6ZQdxxLLmjf4pOAmjp0ff0Vm8UWect9T8ISgFEsb3OfhEMFvk+0OQplNPL4GYI6
b3/syxnH0NvbAJ5yGUNm2I+3Kr5i2SYT4DXXOcTEM6QjZCAMjpJL+E3D6Hp5ME6U53gTnMb4sfxU
4zISjHV6T2LnN5aak+KQNDekPlVib0eHrMEO74udVYn+yGDKfeb1HQ9PoUD1BivzXOYW9/cKmtbJ
3Ve6HnGzqVmllX9m0GuU1lx0NyBDX2YLphY3VMnUfAYFpcVkIK0Y6LyV2WSk/zd+9PvfXGU8LQ7F
Aj5VXUrmffs5ABMEUT2blOzJRWZ9t5DOt0ba07Bnv9k30H0ijuMXDQ0I1DgfvvJZKfbc254ROr7g
tW8Py5+lwcjpdg4KmHRBrhRi8tYKlUaRDCmItAvflc8nEbp72FU+xdPCWPAlfIzj+9M12EkKAmjd
n1Y2yeinh2gBRlDSUy9bh2eTgoZ2r0y1cDS+RQMZ0qZ+QTQRwxAIAw96lu2vB9HhBBTbnNQviw6Y
wauLNJSSszzdVP/lT5QEY7Zx3mTsoijCnzD3+cY/HKlCb4PNW5x4wm9Y9h0aq4bGlg+KyUl/EmS8
m/pxTFlTvSRlHGlUcWTVp4iXSl7Ew15EOgmL7z9g5lyrDklqpSB6+3/g1cEyD1daX69ostaWW4X1
0XHRFLU6ZMNe99Z6h5JKdmnqn60E6zQWH2UznShonF/4yVnwNh7egEPB3dxp6w/quM6J+qzR4JVp
AtyUv132su1MMzNbQqzH9C/zFRrRnz8kE8HXj7tvV7ozLpoeblaFaQPVydplU/IhBM3KoOXKtDgO
267gnW9L6S9smH1vEIEZX0zlUmFKAM+7kefwnISmCbTwqcGu1qHqvSHvti0IBZMNceYMta3W7xUV
u6/+J9+Lei43XWIK98fnjl6kFrjLmiZdw9hAvZ1OvNLhSYgaMyb4WL6PNl1/AnMsJhyfPIJHWHs/
g5vEgnEZyDx19DF3dWk/k+BV4rk346v7+P5Tyq3ohakogI07MW5OXgQe9c+h3q5CxaTCWh1bj2ss
iP1nA0ywK5JDl6+De8aFgOD1Z1024jH4DxIWsNYvNvwFMBcvMMVkflf5QvjecRTGfgY/Zm9Ey3Tg
jE0rb2e2CTWDNqces/o6VCqXiAxWNwQRzLdxU4ouj2ZwxwqRlHKHEe0msC/gYPrJz5oGJutf4cO1
ElbrWDMrntt2W29eXLl6j48Eq0zkLbGa/Itl73sDQ+XFdo77DtF8pRXE1h9KV2q8M4/pGfCn3Gk9
zn6N9Nl8CJ2HGwsxFzV8nQohmcEptBSfRov5Z/Jm4TyPhlRd/tRc9o9MBMs7a6CkajvfWehluQRC
9ttDXS9jee8VsP1BWYDmLPjtIhHCC8xMUj2eRO6mc5ecUDyh8y9DhdLrjUM1Gh5DQ8mFCS29rgJS
myUEH1dRK55WYa5sS862/Uo1fJ+jTk6L3sWlcpwQ2oseMLBi9tyOtObKtHeVgpSKwma1so1alpVf
xiKmiJHD4cTHrac4Lc7wKvLuxa6woky+JUCYNUGf0MM4kL0Fz3xxoTsVcOP39wg9UsyKGYhiW4cB
OyuKZX8y1COPLo5m/d7A3VeHdGq3esHakuUUgb5UO7LAFTMIZt6rscpnPnSTd1ILUQVE/5+iLECY
I4MFcCbhjZmAqmR7XIGTY2QwD71owM8CArjILaRZ4BSkBprq5IoMJx9wVe7Wp0DJUhZsivgGjpVB
sxzbiqPMYovPLvzxJf3n3CKhwaHxs3IdVATxswm6KRRsYxdWImpmFEGae09X+K+YMpy8JsOYGJ8Q
pjhnRFUhqCjogL2qQJ+VyHcIfggyU8HwjWJJN/oxQGdY91DTGlVEPAmU7z8KnXnwCatASiYLh0DV
+rH/Ulo9h8UjCPfIvidoPCpOnD7Z3/aCy9r5rU7cpkIkc2wt4rzd0D6/hGvL55Xej1N25ahmIWZu
3SCdD4rPCi9ED63ln2V0SMbj9eQHo+v19JD4eqUNILHZDlw4yO1uKPUPFFku0NAkS8jX6vx6N7ss
uVUIRAE2v6hM89Rxbgj2VocAHSkgnCf38FomMrF232yavHJf+gy6QKq/erVczaCyoIOMBB5Yp4Do
DbPlV+7CYK3zCABgqG7lt79K3YQbL3e4jaItndCZ1XlaQhvAF0S1N8k5XS1HkiBHG34sNImRg1BM
eoSFX3c94LUQSyQ8fjfdGQzdNwi52U0fUQapvZv77JWDQ4al+jsF2udWmjmFFIFEaWzMTPQkW/X1
Wnq3dFmI1XZGIXE891GBA+XcLdvYWdzBfXhzSHmF8yNp57qBgyixpP3Q1qekj2MpQ+6wwpNI99MT
6EOHYZncedHgOlRPNWGpSde8/Fng3qL6QN/d2F0SqdBnCnVSUPxS0tqy5JRy6zLcV5T58d8kV+KX
Zc1j3zd+pbUkuEqEX6YwHRYmo6PdStvQGCA7OevgGTJkjd8eNxAZYSgJU/7jMDHXbgV+T6oYK8hA
tQZjowdYejcmpL3GomHfsYZqJb6v50fJ8DTyyASv92UBQpK+529oaQGICLF6aUqdZnyCBqcLoQOs
x7XgK5sWiGWVSBKQ4jCZDE0SgBK9m/EQbH11qXYBRrMBcWBfKZ92ovSw1brw1c2EXEK0MRCThPMt
jkG8XhxKB0dLUeNCOp8afpRiqQaMaQU7K8zi1o653cDHEl26giuz97F1jl4SD9XbY1KAdssVoiDB
eK4O2kAgl3AadRLTgh8D4lpXo0JbgGseWPVXLAclc4q1UCCxbF9beWC/g9AfjGDUTAZ7a16dm7Jd
UZUkAW97U4r1djh0947skA7qep9ewbnjMVWfc+YIei6bI7x7wDYbSljxSVZsVuLVu+tVssDGzh86
Qm9CmD15zkK/UpmPNEvl0OM6K81pM0bTyf8VEH4IiW90bGRi93EaAz2uP/Xm6LXbVCcpGsX4Fd9z
ErIuev7I5WCemd+m2ZrziN5dzWimP6Ql7nnMGxu4eGfd/KcOwWANDhuInSAunaf654xdaRQsp4vg
1xuK0FsnaywH+ErVMKKvxD+TEzheFbS4EMPCG7lmt3e66xKK8W+yjHqGXMpFMXAGrR+PjtprN6UB
jVtMX3qutU3FZTT/HF/A88NWXgwMUGFAxX6xPRo6xfwIVzvKGxVdS/fi3veIDWbStdpzwD4+eII4
AA11pdV0TnGOWZK5mTEcgmrPsVvqP46JTqkKk4DR3LUYrK66YhEGF4YJQO54pjVMz3BsFRdXpU52
AH86V7xNub1txYyPOqoHNkieeyjo+h5x6EGnov3tXJCjWNvsTxQ5y8NPleAkeGFZxu0YqcOpbYZf
h8yLRU9qjSmMu3D8531asK46ZoUKllLx5E43uzGm/pMG6Qibec8FPxbiOTDYi0WYpQT7CxaOjsfQ
D764JNfPmy11pjib65aLTu+w9Cd9tDLOe+M5XrwO3ZeXD2/NjaJFWSMHc8SmrPk01QbKZM8rl0js
B4NByz3aSGMIfbe/TJ3FzY6jm6LnuKdTbWFxxjPn1ttllSn7XgIisSlCwFnTuw/sQ3A2td3S/XIU
6IdlLwxJESpv31XV+f9xPXvm7id/Nhyn6QJtqjmGkt3suSFAZAEP1in76cCuFwpucNWIZ6RbhgBt
IQFMc4fTOX8mUXXHHIbSx0Ln7Op+mpDQLQm+dCK8Ee6NtI52b95nc81r3YJqjIwv23uE9P4bHKGz
VAwmA7z8uARmcHBVHcNemrW113r61NFV6lZ6JocWpoF1sxLpJREu4JNg+RZ9zncZJfG+lDxxXVwV
yu81suc+SR50xMepxEX9dgVw+04xZRqNxBOIgEFvvZosC4YYFR4wl+A8FovOJM1Hy+TBZjJwsbL4
8lwligg3DPnJdaLyoGub/2i8HXhBP+GOTrUElIahYDnCI/NS7GBtdpfAs9YtUKk2vHA99cFlDKrB
FaOID48hxZK7wjedfaNbWGulaji75fNslqtZgA9dCV3LDTH0mOphyh/P4+hlf6zS5yXwkCDVEhPn
AGInQqx578iZR3BMtqydWLrgfh1MoXNvXuHjiXNaa8d737rXwj4qJK3fmp5WlmkTLc+2yfWsKvdI
JS8G+PwsPN5Cj/OYXgIhC2D4vRr9RIqYzaAua74NQrXidSd+7ryjsAXNa5/1kFChzPlGcHLulqQS
daCvVh/jx+AWujhK3X3dEcaxrPLRpweOXxznaxsZ0QMQ+aMQcQavbKV1XurQgj5Qd+h/4dicSh6p
9cTa9S+x8z/Z8+Tj4UQxe+upVI4NZkM2p2KX1+ZAXbqHhTLH9+HuMpVe9PgRXvbewt3r8ENx3O/v
Qv/Ppe6URmby0z1PzhajJkQjlxTW+OtPZbWrtN1YiquCMcubhH2Mq93kxx3fZh84mvkUOZuNOr+X
KorJpREPMkxMPNeuEwSfwG/6b4+bE99MtLxmzySAFatjqiUPrwOcnNpl+xzYVcU1NLBGU0Vkpew6
jaX9SUHho0uQezWzRupmC852xsL2pDKNaP+F0lsy5wXBVm8LKow7Qxx/46LydsRhpG7YLN6XYShp
xhxy+DE3ayQ8Eh9ZNq9/VcRhVJC/bxkBng0Ku1Tf/Dk3eN/0WGSZtz0sr3VeH4ZKkyv9mWWAJmLd
7s6zi1E3xQ6MhO3h8GQTe31E4fbN4mYcf3Nm8aSDuz3dSc9i5mGc4v+M1j0ggGl0qXVSsh1SxSVG
AM41vteWmw/U0P1HEEj0bssHJRjID+yyNR0hXuc/QxtCaVwF/mY34An5ajlVhI+47yOfRQOUfZH0
2jAalp7BVymvowIrQYFlagGNHyajKh01BRgevAx1hHUALa/K97fNNzbeAKXoSo4bxaEJN3aryqdg
tH4YP2z+menpeDpqO0kZmlJ8p4EdbBppYPvi5guvDJns0iXAdYmSPVhn3kjflpKhxls5qwAMG+Qs
Q5elhvU7eDLAdf3wshg3BMzImef6G6jInRR6pltdk0cK6x4nWoVKMoBcm8CMtQHyenmP7wezXU3A
QkIAMpEkIxhu1hp9vbt/7bhVVDtjgw8DfTBH9nzFxj8w46vH+B6mIL02RwzHK8C8ElDNq0KTCV/g
/BZLR5IE/DHVJnD0Urws5Ss00VZphDiEjM6j3LfQLo292gOrsn4sHOcAk+t980KHTGFMebHOZp1V
rHPz4VVD6wrHMq99z/QUZtu2gw3bZa9xhzaTtEAzs4pKDej/yFhlK3nxyes22Z7WuRHIUSzYYdaX
RbmUTN4yugI4LIMk75ivma0jA2o6RFYD/eN4G90bp4orWoQbrApd6q74e9eUGSRbtXAeBOoqqlaY
L9OnHaGpsty+OM4+iDxGC01eZ0wfEOSsSOWA4Fd4pqdy2xTwtdGaashxQvelxhTryyCjbzfzH9nC
Nykert+kIsUczT7ZfkQZb40IlZxEmZvM5rThOTEcsGHeZ4HZZhiRg44cLpXzsCEcQBTTTwc0zmbW
cYPuGtlIcBw6fkE2t/DScQbOGJrvGfsRdDyPP4WbrcMFw7KVMAPCazszKLlsfogdDW8wU44DVUo3
o0rWVlVgZEoMqksNN/53uIoixXt5ld0cLTCJ/fB3yLmg1q3sruKFoUeQpVywwtwjG4HjDaxpjv7S
JcJMeTvoCuas4bygcI/NRw428faYwQxGOjh7E643PK87zH48U+cx9gvfcVynB8rHAhz8XNU8Ye5W
UJDhINvr8liA3VZFzsRU94I8RE038tKnn9TFu2Z3jueMpv+bwXvSujVlbqm1ikXNZFC6g5zj7Jtx
VL2kD/zjUPWafeIcUupvdHa6IcYEaJOaHA27d6aMFpf/7Ly6ZKJuhtF4ICxPG11/N3uS323swBNJ
Zy86abLlnXv3tjMMeDywa8bJv4OJ9vKtnwwfkRwvzAVU+LaSG6ediUYB0gcJ95SeKR0/vUkHfwjJ
KPCsyx/pK31XUdci97ynLoKftnEZysuOpXagwUlS/Onbyg8ZWfjtmtB6XclNjCrmC3KaDvKoauRG
9GZqyjwSmoyDJ2i8fA8KYKwrgF5/MmSIAjzsp5+Bp2pIQx+5TsWTPN1W7PuIx6gE+MC8Ja7uYflG
1opqNbz4XyVON8xTNC5wx8PRb0NVy4A3LXBVN4hOMYIv7hjHB1aLgD0HscOhApvqIMPt38cIG6i1
4z2jRX7Y6kcNYduK/GV4vKBO/5H8GKtPiPs85ED3aqooP8tnQjoUCnkOt8DGh8pLn1LxQGT+YssO
8+N/davT7Yq+Sa6SO1CbN3Zg1Gy0fSfBsK7JSMwbvMPnPI1tdh+T8gPysGXFA459WjBr1P2QO2Fs
UNM4JcnbEaSgmiJwhRfkq+odlEP1goAklYDIO0h/DnMwhZ2GndnEeCRAgpdLOTNO9feuHToOZp3R
Ff9UNmSNwZYPXylOqlnOJLH0aP3NvwhhbX6sHRSIpIhHJpUlvTyQl3mDHtjNMu6uygdN6UxeeB3W
rdhHeSUg7SfEMqi1ph5P7aiXhNwlSJoBEryaoSoT0KCSVKoFGZ/Ej0mdpU6q0foDqRlUjgVYex38
HhjSMKZtwGjNLzxrMoiIbgkztszD0/0bnvUFlnZEKYCBSUuNbnzSYFhDXUlRANnxl/FxC+St+jUQ
Ps8t1Mggw5O4MV4yhyg1tJ0J2oYhCd54QvoQwwViwtYQqhHNa0ZySRe8NA6uuZIf7oyBWKxZ+07K
CWL9Drt0c5ajXPcn06IJ3xk1p1eLktH29zlxvRZcJvOsExlIVvChROYIRUzw0n2ENRh3rW2FANhG
nfvrseBil2zfpaEep9HMcIHk3TG1WY+YAJDT+FX6IRUzeodj1azpm4hGOURHIHd4uoF8D+gBzAXx
uLaPIkwU5fyD7wNAWM2dw+JnoUbr4mFQ6rgHS1JQMdQyEdhvMzS6FE1HD+fi2hCm7Gpq9DugEShQ
9F8Zbq9cI8+HwSyKBBiOCijGTN9U/2SHkMY9XgqsXvEZx5VJFJbFD+zGuQCynp6NtIw4B+aYirA3
LO1Brv+Rl4HjTJxNjN4kXbdLAAwi/gS0DakUJVZr/K7KQCQr513TgEwVt9/WDTFMmZgUk22Ejnkz
cbcQG3fFHrhN9nggZ9pmyRg4Ej9qfrTa5iQMYpeCR7JR14nCCY3U+Rv+fBJcxipmuIzKme21YuEX
VuadEAFr1QCfl9c+7rzsG6orMi/151NeVJX0mjh8UK5xjubscMCc28NfPfsB9FtIQLMCtZAgZA9l
+MBx5tHr2Cd+tXNyCnFrEsxFchgsFY+kPsqkWGd/81wac+wK1wr6SAR2wQ9CIpEsrQpOcvsc02mc
yoMQPDTCGPrD7qlkr8TsnM1tUY3tQ8JYRwA/5UthU6ocmsNkZvMzUrqCMmg5vlTYV8exbvLqhQAp
6IIIkvHMFuRc25Q7KEFIUiFgmW1l2S+lDdSPGo0ZDbbVeVS2oiM/fuf/xa/qyK0eM7I9fD28JXar
c1aTt+jZQrXIQcpMJhKSbkKZP4dAM5vmk7tZ9eLTYk87bHzaj7j+QOmBnI4Mll1V4y0JPkzQU3J5
pnqzqtfEHDF4qHq18n/5DCTRiwEmr7eqToY8K0c+MMuahtBgoPavQ4c50yOG2+/u88rneDoSeklV
r8c5nI1+jALst2SC+an+zG6nPC758tvnushPKpx4JcbLkI7KTuidXI0+lQ+DYOzeebrLOXok7Atl
NUd1I5ho99dqTsJwcI/UpB0r19gkT1dv24xg/LBhnyvVmDaYPfv7GUT1u05mLG/5IH6LXBhDeP7d
IzZsWEvOY0cHfsFLgdktJ1q/aape49qmSXsMWaS5fI8b7r1Hzs3p7Gq6vajW/D+iCV2nekGMjN9+
oAhTtQw2QJEK7ZbM8RZQvMjp8wJQouulrRe3vMtF/vN20zITLDoyZFXLxTZFfQJOhaDgZDr0K3wY
9E4gG/orFojZEiH4x+rkP/OydgGV1dVJ9AY9dW4oxLsGqApudsamXJqTake2nzHgeujz9vJxXgL+
TMfq3S+9uv09at9IYYIXJsjE4YlOAI1bMwMUOJZDdm4sXrwjS+ZAIUfYGpFXVE1W6YASmKe1wTgu
1H5s1wIOzZCl7mkDkzIYfHQzCsAN8+xTBBQ4rgjLW/lQXQ/9tAc3nXh/gImtMGdrxJzrKRk/nVUV
SX81/M7N0BCV7+IxOYvOoBPjbxjotLlkRvPfT2GyhxThCRBNIqBqlXdpCL0y1XAYl8gc6eDYInd9
o1J7nDW6/RLN55NkQ+VPl7auTcTr/ioiaEH5L1GS0o01nvFueLBR7aC9XKX/LqK6PP7TJ22357iC
RAboXc8I8LgbJ6wPCi42P6+ooDEzUgQMnJSRhJQa+vNFPeHkwqcbVZeNbu17R9SG378tFprUom/v
c80PtLKxJKvwyxdmQYuRflAN6+nd2m2SKTWKHihSDo3W/yqhVDfL7Q+WrhaJYt1tCNGo9IUeSooN
MFlVykXtXWWJlwjvnWiLay/d8WDtWgp88A6QjrhlnABqnHDYqbTY4OG0pJP+0njwR5M/CQk4Y3X+
Lo9dVvyYoIAEiC3bkC2314ICIIl7FVQmbEbRCh38NLMT48aeaK3I7fpsfYAGDrkpBFkymZf3pPzu
nzAOsUfvELX9MmsOYDNZbsBKv+H/Eak0OLhasHZyDykrtxumYqTbOAOtDNRGuC0IQ2gnnwL10Hw6
+CWYQDWM5Z/lwOsp4KJe4l1YZzqlBFb3gJ7rQF7a64sRQHHUXhOwc0q8w4uSF7/hz+MsDHsM6HEW
HmHMZkDO10p9mesL6mkinLXlJGajqN/Eb1QxROr03XiZxnSCNU2wuv38WC99yd2PUOBHltf3RyFV
87mEZlBUXhNq92s5s0LSY8k3tY/XXULUSed97UOGB6p57lGYu+iorsEuXiWhpwBb3n7sTYO1tRPY
mcYt5vXz+A0Tpmgfp954Oocs9aX7PrKMe/zc7HW/6mvfhmNkuPbLmYlI62J1VRSTSzKqVbyhKSnQ
IByPG70lzvUr5893hXru8NBdHc3IfYcC6LiB0F9KBYezKe291+fBVyK9avx6mVHEImrGsdX0Wdho
C0325Exds1M+vsBuGD83cHmYRAHJE2iJjoKLP4N1HgKP4XnRh289oahu6am3TwQIajhWIM061HJK
WQJmUa9cJoAXCRkpnNGqLkooihH/pzcNidavKTUNwgBhajTkj0RG51u9lqPVv2Pmm9eGp1JLZlPp
QODyl1NJGhjxlwRzEXqMvyQlVQRwFR+KoI57WdtV0vxcD7Mawpk99QFJ6R5IKm1t5lrza3xgYu88
lE8Qce4PmxdDFDlaLhgsO9xJCRc+a7BvRFNixa3gT75bcERhJyBofN7vGmZ6l/JP587YkdSeYsJM
9LrIi/YeCjoDoGgE/4mCoMd7wCHCxdeJX1PhFXeGiQ3Nsh8rz84CSJmrXScqmulnkAjOlX0KPcjw
0yDYMgi48uWQwT7CXtzf2FqfGV2PxvFIPeS7PwjV+D2qvrO+Z0D4uLyjqgfetf5t3ojuK6eAza2F
er7h3svcMvyMoMdXz/PHjtO+2v6wr4Q8PmxJYcmccYRV8UQsKF2OHuDynEtS9ww7UwX8pSeToBwC
2bNYlyYgBjtoJ96g9+w16gXhLZrHkJ+KKThrvNA1APkiV+e3Dryi6QU4QX+5dseEjIoHFRwm1M+y
X/RxEypQBY+fucTBoxkrW/+XgWFaH3SWG93qOsAexL5FcQAU5ghmiQpt5UxeglMhcsf2z/61g6bt
V7kg1n73HJvfeg8hBmiD7YQ8AOqRKJYSvM5KIwizdlZHmy2LL+I/f9lXC4x2rDWGxOBBCOR75gzl
VjQE833MrXTWidRaBti4veU6UVSZHW+nxgkGnmWLzQy0A5VLmFM/dxntSHkSZ8bg556RnDmRnf4i
4lzVq1UIvonB/yKnp3FOCIL28mZ9x3nRqaDUEJaHtf6ZoVhYd92KXIqjCTq2EGCrJyne9eWnG9YK
17dn5sc3GwBNd7jXCpK53+6wGN4EpjJ4XxaUZb4GJIYMb6JWdNE2nYPjonEfZrzeONbbLO1Z/N8r
3UvVaCvxwKvZuJPkcAVj7P+NaSU1TYJURutK8C1q3ZBIfWnfjA7VGgODEfLtf8fSbBXGJp5auOM5
UB94KmzY85b+ydGichXDTNFxh7UcWDqmYdfGoM3xa2RpXhbpCQyKghDAGEtpVp9LOgQo0C1X3T/t
pnRH4QvB1fv2FhTsbUo4soh9KVmlvqfymBGy44H9G3qli6UY4LgKqC3X0v8B0nNPbeFsJAf1Ztgh
4dg5jKsyvjsUmiQCtA/HI/qHU5ws7XtypP8U1H5JJ8PXL2a3iCPb/EkU89LAxa7s6P12RE4oy/J1
h6MVjs1VvfiZuquV2hC2diZAw0tgs2Lfu11/KMNqMzx2f2S3/Wdjt+Nb18yI6ZtkaNJhbWhJ8hiC
Y+msFOUA53rB7if3Y3T6KEm9543Ocm9eDR1LhfbwUqrceyocFMGsWZgk+Rhrw+XiT/r3gDCe5T32
4inBRhct6BA4JF53U8O4DWNSTJSN/Q8JGkODsJ3lFLtANIEkq6SZf1aM1cwr2xc+398X4FzcPS5d
GkPzvWqxRLlw/4mfDcd9X8P+LVrDosP5yg9YpotImPZnobrzVef1XCKmST3L2AnGMy6vaamPx340
ugfkS2+nYUN5p1Ccm09XsgpDTbH1hlCw/DJ9O0YPrTylaAOkW6POcPqLSqECX3S0uqhq4umk/FRi
5ovWg8AODxYufQ7Kbw+oa/O1LNcZZTBPGpG3ghz3Ok78/76aWdIhTAPSieHjszEfP3hDsJ9ewWr1
vS9tCSST29kKpMkBMuwcOXYF2S/9JI2uiUk+3HtpDZ1GtaK6t4ElRaTU0OzGNUXjHwjaOPcry2C0
pKLGjTiOQ3UfTsrYmToXbSF8cNuF+ruDe83GN5LaGqLjTiNBV0fh8h8bOkkw20oYOw2NvnAb7+TM
HuZ2JezWlmANJEYQss+QThYBQTTF9DEsm38w+UnxoTkcpe8X3f8Vl68LMixi2yGR42FEJlrFG4Xv
5F4pdSUz4NnpDQ1fgR/cw6jT4iv1VwJf+G3klqVP+8t5VlP5E6uApyL11Rv2NHU9/Ay8T7K+etoM
HqLUMppSz0vgdR+LOo0dUkYMh+VqqGDyid5GeUulvbeT8fXenHZ8gLz7Qm9SLBLqpHjpe1jFoRzP
8Bv5/KVz4AOFqif3CjvUKqqu2u+UPQDAZtoX0n9Pt8z/HYQonkMxrTeLMZEH0UiEXg1qBLuwQO+J
wjMy255oNM5OK/8J71+Wm7KuNqwhY7uXtuax8aOlgldiWuh37Va+xjm/6PWsXIPs1Dt/m0HagCLU
7I8Cn2aq2833SYvsqiRD6k90k1+qfCIALhoQLL0Rsc2wGJB2hXVkCmuVT4WPoT6dJX+EyD9TNYwE
SFKuOBVVCjIEeBYVhLyTwAA+pvzHKXbNl4eIEmgB+obZMZbU4oGWMmznSQ0X8qsw41WwTS65h+fu
BWHfUBP0/wGdDA2q4XeugtkywWZBFNKFFxCfdXWEBRcOSwswKTHuppvq4Jdy4bJsgGPwXpZcmsih
g2hNdKoY0WxypqPhaTc2RgTWCNA7s6KIf7WYgbD4heHMLg3RxrWdLnHgdURE9Vd6QNh62x2lSrHe
RGoACnDCaf+De48obm4YNs53nAnwXY5YiTD/FsGgy9TJHp4//+0FjEtds/wTasgFDsSadoxDuObG
yHM9E7xEEbQXQqly+op+uDhqmch9DLN3VN4eN1MMylP+EBJcA5Jd4W93jLJGF6Lh1Vq1ZMGVRv58
/IyHBvzw456M7MpleWTzICSvK6y/4iFERZ/ZKstlWg04LrcJVZSBZ3Thc/ELNk7Yg/gYOxyoyiOn
jZAcSDcimIdybh7Yi9e/IUpiSf/m7skdJMq5DIo6PsGLILm6m4K+BN1+4DdTFZ7MQHOmtqdPv94+
20W4ApNm97fcuYabNg6PICx1rS7m8Sz69EqTjsuMWzRQnAtVQWooo51mORMd0V/MGvWCOYeC31Xk
lA43K5FXMESMlkKY4OquiZY0MWd0ZM778G4LgbgkzRKmIc9ett6b9O1B2QsJoQHWbes3cFKz0Uh/
l0tZW1FC1TpI3dbDg4cIcS85CqheJtw6rkTkTnZ/bH59jhd1L3hBiRKK62+4+XNoOBshh3Slyy/X
radYGO3q9OWgYt+lgupztTshn+luM3rOUgKQ253xW5W0cmvUbpI73D76+iXhLpHxKO2DT6bivQNY
2eKEwyuRBwieAHLc9f+cwuK5cmIaPDBcbvbKIiX72AnJ68fW50rUg3i9h1hOLmPZr6wd3GXMiesT
rEH+T/7q82MfQOU8C6uXhqsyiZdNt9S80fnREvu+HPwBqB4emwYA0bQKPVpwJ0UA2jB8N0Qk8Q1t
BQ0pKQNaNF0pzF/6GycLbTwNfCiC1cV9/Xx81c/mPVDzuZmg4SDVyqYeTVRzhNs84Alo41Vjuunc
durrDykZyPjvGuW+z7rFuQn7GhmOpXZiwNQBsuU9lTqG4g3SpLnI2dev4WX6fNGJVKFP89bsBUEQ
PiabdrXDexpBSrqQoHMEh9URBVMfD4OpboI/aiKY95thsr+edYShFuUweJpsIkti8ec18iVlJXhJ
PnPj8pVKlVMqcCJCK2I9MrK/lklvCadHyy7K5VfUBSXtczYzOTPMT+rQhZ/qFpGsRlkTfsDqusJK
2/PgfXPQYE3RcBQpwPNPt44l2/ZcKa4S2ubGHgNY8WLA28/BXxFipkMIEfuV4xYeoOxvYIffb/1y
ogxDpDdhSJ2251U32NKDMNIm1A8Y4U/R9lvM2rfK+WskGGYzZzQo9E2KX/STJZTmihQzPpWg1qEs
MJ4xvaL3wb11UBcqqBK4WoIAHdew1qx/Fk5KKKCGbbdNtaghXwzLxkrOjoH1Ii+KXkY5U5x//6dR
qecttdY33kEcztPmsA9OAZBrxpVheZ7QldHFN98X6ZnfA7CfGXPv1UWXs0hpFRgGDCoon57h+Mzg
Q1pebZfyqYReV9xdNggIPEB0EIcyziHLi4WN+8t8DFz3S+CcsOxa3k07p9ouB8NftZXmGOA3hAOI
rLTPAHnV2hbxgotIiB5kstgeQMZILo4uMNnKC7Vlb/o/VlLJKNamB0apuoNol5rVjP8rUM5Bf12x
IcIrSZAKipEee3rJM6HMJx5E+15UlhBG5sTdt/VXx+7qCWc7TbtVZrZ3Ola1Lk9L1FHF9klzXLJj
2j6UX/6CSNMnxaDOMKk9kGm3hGy2eIgHSUCpf/Z9Y1s7Pi2fZ0ENcltgXKdez/0lfvL3XBeMlMfo
amuVBYmeDrKs2mGVezvztMgCCg3Z8cqZ5cf7fW/CzgdRUcKe9PzH/enKTEBPoAeMkPhOV3QdgYhN
bG2d+UKwSPzSQsm8spSgcgI/JywJQ4p9m5OZWO8ZZklpvM7iaZAFin5OHeq75qnAp3ILtmUkgdIp
4Uara5nLnr5zORUCyi/YDUd0Dex5JL059rkcdsLAEzpj/TVPpyELnRSWGD/5z6sXnDX7QVQlLvVU
NrHyyB4jXILFyz1le/ucfhA8HBKRgvubf9FsIWf22Mv+mioqEYuQHZhbtgFORAIhfEzlE9vOwDd6
nrJRRql4CTC4f7W8yAwDkoNXRU2iCpG1d7YUD3Hal1V5UcrA7kntf4n9NASsUA/sgGso+nXUVVYg
3phDNHK+RToqqHNn9J+PE3vE4QnWVhjqmfZUg48tngsbxoUqiukpgtSqqdaOTmVAYIqmQo7tAIzU
9Em5Xk3Sv4ulIuNt+jSPW2ZYJbYdyTO1eRQg42N9qBRATkzeUIIEySO6VBPNsd+firBM/6jvbfM4
boNlu0aFubLz1a8pbmoLM/CkLKsB9qgZrxh0SfPr3GcicX9S5msB/j1re9quDEjX3LysMPrWo8Om
7Y+fxf9Yje7Dckl6mvG+l4AHlLQpmDQ77pFCsN8K77AycZRl2TivQOBNyTbjT979zRGv4AxDjt8Z
dzDFJkSVQvzPsRtnsIabyq1ylpHmOBG2+PeFb2qg95sVz1/HAMulpHgoY5vywlqJHB6NkHRNN0SI
kx+kAC62bLoYqpiCAXNFVb4gWXRtx/srsSWq3c8NRoEIBO3AEi9Gru+mKVZoEN/nh31mH1dnKXzO
SZv66B0JX2r9OH6YI2qvIx338PjoGNHGAy41DMPyWkhsCzIZLl0f21PaS115u8g32c7mrE9oWjSh
x8ssh0kJay2Ytm7MGLJftJQV16/OpevcgmDECjl0LB0lK5ckspzSW41LW1F/VwnDJv953VlQWOGX
i1+Su22n6F+L6wqXKs43G3isqgLRbdx48Lr3J2aXyyORYsevmixbugtirb4wDI/BYENGQTJVpLPg
FqWhsj2NwUVUuFqpDitAFXRqgSb+kVVRHbks9yKJUNVdqJ9ezpBHlfezXkwniprbew1eFaxFHN3S
LoFAdWnL5xojFLFfwWt7u9ac6qP3s31NP1/u8XmShCYigCqgwEjVvHc2UytdoKdB+WVom+u4GYoj
JycEpPEOSRpvgiTaWvgW2UpPz0m3xszRL7WQFc73JE6SGJbLR53vtK7XbHZQd0Xd5bm2hU/8Ewoe
avxoECySafzndZtMQZ/4RH9TVqPSU3ilNqiDm11Neas6AuqEpOBx46wNwo7bIjcutbU8VqwgGDzp
1zJhPXDg8BqDrVtS581RMAKLx2bjG19QkGRafuG5NyN8LwBCU8tNZX4L8qn3/LW5GpLsz4+rg2qa
rYiiJQ5VFjXRSnzh1tkulGOs0oPcd75gaOb76bLcuye1KxvGqVBPnV7KbUAYnOsaFlIVZWRwbS1z
64WLD0/EAhpDSNSYCKN3tc6FxoyFMEvpjNwpijKkGDUfiG4ejUY8vWdDNnuRrD234nAtZ0SXm9/g
YW3/TIRjxDGKoWm7Krh5+04ixD1sFDqc+hmQKM57rnn361zaUQgfs4IPkt9kBpalNhDM9bAMHIqV
wiStJwqDTu/+Zu4vqETGlxuWfsS5ReVHvQ0w1DM4ujKzj6M48fXLHVHsvCsqoyDSMAamMEj7FIU6
YKOQ3aRSaNp/FCmYOc17JxBiwJJFq1FZGeTzZWcclRCppNNc9J8BtXwGcWqi5DdaYuKoaAKAuC26
XxNZ5mztqqMzOBd0c/nS4oiZagMPjYhnzKEKcxQqVn4oiP99dsWN0pIXkBP4/mQSb1XEt3JimIfT
w5IBAxUsm+cW4VaZZ7hHjeYCwF3aQ4yiCvvB3yEM/5ObzVlrb8vbNL0UyRF+r7VcXK0pyMA0Ny13
OeFYY59DwZD3hzl14yDNt1vnu1CjOJo4Gu0E5zEJQqx+KtCiG/CWfZ2nW7ApB74y/z9+zUkftmQv
VE07LToO3X+72maHRfiam7MNw3ZOYKIgqw0lQFZydw+A7JhinIEf+ncVSDLMkWEiW+QPAyz1dAT9
Q9E11FZ7sz9YB1+3uo3d/Ny19kHK0QuRyYNEH2E+FD5uV74PkS9b6QzVttf3TDlOa3HTkw+ZEBzo
TZI14AJKCiruw/XaD+hCUZerP9oLpU2s/681+y50IdnUkKOkmfi8DJpgFWNDQVZX7LjjfgGvnP6p
eGiR3SI5ETRlmghP6OtF39PyeR3UZmucQNZtqCdI2uJ8xIFcG3D1asM+u0e39TT415U/Jdeld+rX
3sDgL0MH/jbArR9KJQM5qqw9vCjrFsB1wo/7YvORMnV6hQ5UFeLqxh563J/GjPbRCEgS457JZBBH
+vdMo2aiVxaM52rQDnIVpT5h9KDdsSAK9LBAp3D5PiwMnH0IPBnp6hDsmBEdDhmeeRRTclDZPEVE
094TSksi42WycpenQCnJ8YjPOHHluSrklUeM7L2KL7o3RhKZj5B54RN2VtW/qT6zqIBRholPu7NL
IA2us2uno2UFOYBH14OgSY81bk1biZqdEfVWjmiL3kuW8SxwUkhPKWl7+r2BIq4hddbwDhAazgKz
K9jntl1Xq7wVEGWCEN7KyjBHfzaknPg8F/V7Z9QFUOWC/zHGY9Zy+l9rleXbo5cByrEx2EasmzBf
NsuqlmDB5BiAGEZII6jxhAh/suDGJOhgdzlvhaB4QEmrYQm+Mh8fnfWwB1qKY2jRjjdILNtlKUmZ
Dn9IN04MghO4MUJQWIiwK0kjcLrGsAb7UME7bkOWxoJrgMhiRUqhI25SgisBHCjxSa2C9zMx7oBh
bI914QA5T+zs+wWuK6XPsNyDdb6eYABpuv+uHZCF2R0ErYxgUUe1VkNcAI8oq+x/5EARxrbdRB8k
0kIISrOPNl1WZV6D+ErlrCleLC6hpU2pNjp5+xRIQk8eHuo6Fn4rJ+IQVaMMMXyu+pCKJqwU6xu/
erkqMheNNg4co6CcTfLXJRdBtUDkeR9zaeNUjlZs8NX4UV3bxe8l0uzeOlXDU2AsfVP49LxaXzM3
env5rKJqR44SIhnRs9ktfwFx2dQ2lfNw8j0/wxJCkWp0p0LO36t/L5eXRelI9SfBxheyD2q9i5Z8
gxUk9/IaioYJxQ40Cy7zDeN0OOa1cbV6Z+INRVJbZoymzSWQHZpZPwMtGZoH8egZWXKllf0UBrIy
mEeY4u27kIV5/NcTS+FE8Z+WEiezKXD3hZPNuES/evTUTASv2WgF09+Alkxko7jI5A1dm3sNxJui
M4cLZUC6xa1ztzowHKJ/QnA7yXF45auA0RoKE21fZZSZugu3Lx+Fc5LcaHDqr0ESjv8+7MYsakdu
jS4bhm3AVnE6idBu+xZwBEKNNnR0uACBjwFg4nW0diKypXq4oSbXC1u5ALOCl6aNeZWxKoAUqUch
tLrGzuHLVE37aUJ68UxHFpwTtoaUbh8ECpHIUR5XkOsG8jZOAm+4o8qp0l7pJKv5DDp0/hbsuCyM
HIXwMXMRcfieG/1KebKUCBWNWddtSPX4thIAR/WjzwAv3J/N2vBTQZUYTI+WhpZkZSdGjjO36TTx
baA5Z7AGnqayXQZAV9Jyj48kXZyrSYzMbj0ZLsWPJygdPBl/b3SU5puMxCUZ34SnNj/HPWHyf/eM
urWrRYdN+XCdVfcvA5hs4HdlAj8mZ5MU+DMb8AKSt4hdDiDNoqRS+W6wIF/OSQ/KHFwuaGGRLqx5
EDN5ckSXH7Oj4dFWJWMm9Y7mah8MkfXHxrP6/ESOQIw5i/IZULVExwnXtUrOBMxeaZJyT5sFDqIE
uOTB7xX0lMIIov+0+b2ixMDS8vTh12GeX8WH/sfFuOSE/yI4ET3E5ukWV1Ey8iIXa62Y3ATca6Wy
1X2uSYUC59lXRV/jnrgT9dobg1go3CrebQl/CHpp0KKs9oAPpQ8VkiqahYNNwtT/bk9RQkBWmFkL
ervXoD5pgvKOrLBM5U6ax0MWeRmCgnB8n0FheRk7tOIwByqqtTpSGxMJeeJMPZkLglzV9dJnkowZ
FHmpZG/Bd3QAL7V4/XbyxL18cZR3/MGLzlDW9PdWa0tCVgBazXS82doouU7fZkdiMwGPcw1OIV9f
Tw07Xws4AJl4JmtptTVPWBInKquDg/NiwPzCb9ggMuduUWqy1+mdNpHCvrewe+XzZyUHR4PR8CtC
jGWMYMngSgMvRExViuFHatc/dpOjB5jv8lsrRci1dUamyvpXfn506Dw+wR4OqWic7ec3dbneSfpp
saSzADqMnpBAhS+WnjsqLxD5F5Y93UY5UzEZiKK3HGsITfHuRK6kZrcB+dhLPP3TR72VYxYTiJIr
iy5OVXfwe+nfEQq9QT/4Nve1W2q6ZsY5wk5Qgl450oVlIh1jMXbEQ8Nq9ExoMifAUtqzY+urrKEm
AzstnSh//timGdYfmLKcMAdObjdclCKt8nxVGjJBambAmx21gI2QJOhE77AGN3SGLZ3Am2mrExxb
ES+2t1bEzaLxAXAbRTsdPlj5Ad5GiBf9juLL6xRn6gpg5p51YvJf3mNn+Xv3Cp+F8FMRB0X3uxgO
id3ggXkrSQCe2WhvP43QWEtgDAmTLOYrdh15MvSPNhFeaQ96OIzUJPc10jkEOTLBTx4W5xtNVThd
CjwfnKhbh0xPsOhzA2M1I0/RQ8Ks37upA1eM4QF+B2JyfeGaB0q/hO6cQnmCokhcB571izKoqSp+
SEQU6G06dA8iNdXv5JCADBTaKWcmZXwkRrep0HOVNs2GKEEG2DWyJS0+wtv/G6uwnuKa7sK17fpR
KjN105AVegszRAwRJ96f+L/R8zE7g9w019eLSj/Z7xNFHoGc1HpoXKDQBOcxYB6SrtCfd6AHPeKm
6P3SSCU/TVkiWwQNgfs9OhLYBZmT3xzpHbvW8o6/S1S8oyvF+j0y8GgumDEPIW/5ktRG7k3RqldW
NvQ8dF0jG3EuX9/w8hgpIxoBGo19TFyKtDzDsohiI8g1Zq7iJyKbb/egFZGAgOM6w7zbDaroOrTE
mQ6P3ySg8QFJl+bSSpQx0C6VloxuHsH2pES6Orip6TiWK+c8WYeZDuAHlzBkauadm6rSUJ7EovZy
XmZdOFDaVdSOWGu3p2E72zE3uwSHXeTq88/JJ7rckCD08nBpSkRfpVUvLt9+MaUw5N5LnlfCiLMv
IdWOnZHgeLbbIG5/6BeXr6k7E/NQ9xgKcTM7y58ERBiMrGlOwhTOiPdjQ8cbEPShEkq8nXSfgoeJ
BcUHbvr6NAX8H+QBvc1NypcHkpLVCP782Ht6tfZfdbJI6zwAQ7E+XNf/62na7Redd7sO5XSAKeX+
Wt17ZfY12dP0o9nXrn+GIdzqBOYzbKS3UcmB0kAdW6KXnKX+d9oyesl03ff9MgEGKP1Zny64Y2lG
joxhFFMMvOfT0k2qDhV67YtvUHPrSauoU15+ia4FLAFbujEFGNc3rJr/s1dC1a6Ls9dhYqrd2X/n
BeM11XVoF+BxEl6SMrLalSddqg/qTVzERUQXtwXllZT4rG/w5GfUB52exqPQdv1ESbyC8Tv+Zh8E
GELKJI2URWrECKl2SWApbIR10zoi0jxikWoQ7EdOOtiFkdpuLl9SsJrqckFpFUsxe3+BrO2NYEs6
IIkhkn0tBwNqRM3yt3TjrHuZ1ujGYYxEWJaCaZLk1D6muQy2AEI+uFFT7O1powKEHx6efqOi3GhD
w181+6y4N7DXvy7jIbMNFcB1oOMEGVvvmOkiwiumebz9hQkdwosboDQMjapycWBZ4TM9bzB6C4KU
zubbRJDcURBN1H7E8PWfVM7fOltdbDTvtGbJkvpcyfD0BeXM3IqfxHQldnxiZZh+zhZwmMmHJcYb
OIz8yN9u4PCw37cknLhpIDzrd/xKiWvrplqeDYdfwYqi1zj7Wf6fBEH9haraMGiWSb1G34NT3fu2
iXKOTAneCEVVp+p4HVfPt16M9hXOEklF+IxlFhvnTidCzJOa2oa1Ces/Gfj+7LP+W0g5wjxpOig1
jewL49LAVjjrcjHp/kTtTRkedxkzpefyrW621n11u+hLltyfin73X/nrzecrD58zoVDaTLNKFW54
R6l7qjgOuDP6DeexAwag3ZtBYjXkJDQrd2WOvmuOAwVp4MpBDSdLY20HbjJKuysSLNMyDoSaD8VH
Jh108cnWXbKl76xxgakOXPigoc1tY0lHewsg9K0al3EdRhQk/ayJQZMZBu+tlunwowjb+LPHOqvH
RhtfolW4fdxUotXDbbwFFxN/sKjKbrMhsET1A2pxqKxfRU1Q+ESxagnsSn7xrM3WdWV/P+ao7jOL
FicIuPtXasLWSV+RlvyHobVoyfKKWlrrj+euMorXkO+PKW2g7e5DYDGhan/CjybY1z8Pr5csZnYB
5A4L7wQHnHgybA6jKIOnYHURbtZtV1EiNocmsmIDcvrKVHAVtj2mJr/oMVxdXlktrgY7jMccfJ0m
CwvKATyyRYdFr6ldTo3UmzrJwC7xuSN28wGEVtPzw5GuQlalCUJoxVoxUSLaIXWuBNpwMvsJkiLM
rIosoqjN0DgMmzdEzLomLnt9w7uLHXM9gjr+WYaZj8a9Fp4HjZ7q9uMp0LUTQRcKnxFtBZa5tU7G
1Gq4B8g1Pjc1kvJ8IgR0lMyK0XD0lj2Gy5+BN7/YMrCFpeACub2aYKNxJi9qskUpufoJwotFXTxX
Yzno/jnxe4217uwchnsPdbunWGKdcfZu1sVxEtMPMbk6NZD2lPWUbDZHGUL2sg9N6bM9oVc3/uL9
Ec8UOkRj34dC2U3ytGg7rdN+GzJATKz5v3d5YJO3waLws8m2P/fV8ZlhxwkxQYGNMxJcKY/Q9765
Y4sMOtt2F1O9RT9g1cU+x0sjzIlvZwuy5kXPsUeilfRNGt5GIvXPued/Q52IalBen+ugVSUDWYFb
luCd/nBgIJuCsgy52QgZwcDiXY6X31+0vmhIrOZAGxbL6Sx/nyQaZCP+6tFF0vFNwKmiWFmcncET
0eetf5OpfnoE5pVgu3ivH0NnRiTJNO4bt8IHxQY5wIGXpHSWoSSGXpFYIyFNHGytgN+ZRFlpi1wc
tr3I/P5huARl8l7JTgS6vtjk42b8fXVqlvd7eqqQozCH8XYoC7fkz2NgTpUVjXlQg6H9c8xZAG1Z
8hllJ/Uwgy6+hcc+oqInYhQJNXRVIHY6l4kS3xn2z8bwk/syor91CobOS4w4EZLq17z2Y12jElaa
MbkhJmnxDRri2kcZFUqQ/fcYsL64H3M8aWnXCGSTRnqyQ8cLgF7IUIs1M9KiEWSG0yQJjIkIXtHN
9GFNvBzmwCI/chd8sXAz1QJjdT1BnwpCXSbfjuJaO3/FpNFBHuB4zGR72qpzlebkrgaxeShKyXX0
d3xeMh9KN27iSp9RDGXelsUISABWCI09v/oxec+NoH3YO8JvtsZobjbVwmB4HEKL0tbO/Un8u2rP
h8L4K7SSwr8kkINSYn4ldhXG5YxkgKO6vZcjXVvcs0nzn5gdUcJdtks7aogddLIatCX3Ic0O6Xbh
RoCCTGGjavIOBoSRqMbUc6YYqMWlHYYhbauXBUzBa/bBBwRTZGXN5/akNw6orpyflZ+IWS1jL110
t9S/dpN5dWZ8vw6dhDTwmd7UiYvBy610M+XrmQomIjUZQY/bXc/Nhvkc3FAnMAxbq68nBVSjNRQw
AnTiiDMjFZTFgw76X9e/xYAn1Bm8TM6PhYcaf0ph5yHL6SbQBI5VvOncvTpoOtU1d4mDH3hahA5R
O8WLqv6h/xeh2MQMR+s98pLJJDqPpna9j/ZDCoFIdt1RbksGsdsIDH2GYIVzAQslCXU5ovchFpDM
HUHlogUIJBCW70Mb7j3PFp5zywQUohczNPzveYJ7c1wVXx+5O2kW+d0NiS0HeVuH//bEKGCGxA4Y
xupc81/rZC40F7tMEAsdJQjRJjakf7yeQBv9H5orDBqjwFrtTvBUpNrGkv3PKT5rLHFEmDb+usFE
YNo7bx/Vm0kyTB9LQZ9aoz3Qm3uXYdinjK5Xyc75tNScm1BeGst2US/lV6rlof5OHDrRJgSnXqsZ
N4U4NxkKFcyXrK+flA1OuzfmsyUHq1ve5tsJeAczu6jtXfBOn2cPfX73VgRfvDsDgVPSmASMHFrO
mtRASJCzmGa7jBgT+P4lpvKToUV4wOv98hIe7l9hAQBuYi1dRQLFcKeHfGpvAxqa43xkOh2D6vv0
OI6cAC1De115+kKwkGvdXii+9UF7CFlMxG/PdXzJ7mTgpQGUXIjEdMj44ntyfeOB8PftYZ1nJvVP
lX+0T12E0WxGw7eeQqnnU4+uwipSRE9KOuF1+MyV7NdfLtxN1vtJ0z7p5FSyyh4IQL3R6MoHaers
oT87meKEZeIdxHPVfCMiRUD1Y/Vfy97htBVRtESrqxQKjyPBIZTGq2szHbu6Xp17IEcBty4959du
nuEyibLwYvWeiDOMLZ6yXamw6EEqEDt11v2yG5/EAktphMEOJTihw2Zvqi6OP3pQVNlUdGPQ0B+A
FT7fjJQuBR9M2r5qCk3K9hdBvjwH65IQmjVcwVdQeX3rRWu3RQkw5uFaOg+4eGKR6L2NTL5/UlJx
qbnZoAmbrn27Y7X69UPO7x1mCrKsg3c4zKvYEbNx+BQKTB4zxJ4VkxcNZQCfLYOJXJ7ae8IrYVVU
ZbemQuFicnqMakSnyOjOkUTpA/TbP9mHNIgYrPjmi4JMs1nADOzlhGbVMNQvhHuQlPypUUtz7fiY
64C3FT6e/JqTUc3slLiTMG8Oajc6R3fyumwY5X4l/AFUyBgrzQgJDR/R6/0oE/00fqUlcmsxt3PF
mlAQgJvOsoWv9O7oVt+x+rfgTrasuOZAziR0NBZt+jcybrdA5MkvXC0cI8FoQuXtOkyvY/8gjfZA
F2o8m6nWCr1FCfkRkdbozhiX0WSc8P/Gn6Cyb6svkDLsJymvTcdsgmZ9yII47aEEDEy197J5mEaZ
+HFS0PwN9YZmiT8yGRrBuLFjI3K1SDXbHMkcxd7f8WD3JhL9uROE165thkUvAzjq9bODPv3RGo8F
fKHgEKiD0LJV/epmSvbhmccXH5Ixm+vIbqGF81w3f3x4Tgg8CjqZe7aW5iu97nnkOF+FFjw/7HIW
COjREtge84bTLctzS5sWh9bvKXk1y96AMD+UtMMUujy2ojSVgv8Ug8xUqAbqhY9DnZQo33C1uI/h
yzpcGpAS+gfVdrVS8S9hLx0fZHMnw+BxQYNE2BIEW/s2jMrAMxvlOIcs+9zXa+No4Eu/qoHXhDK0
CV/WgPEGSt3ZSpvw3Em5danvqe/vks7hxi1JvbAgzDk70fZlhragP/3v/XI2xMxNpYOcKqIIu4x/
TeVlZhWngdOgB0zwk4A5am5JlEVeItym4FcFIQqWHcSE4Cffz5jcCyrfZCxLsV68HGd51jb7W63Y
MA5CVoBuFx3UzL57IRqn9uUCei8Y+BM0bkzuQtf+FXBLpOZr/rFEwz6jl5HvINAgPX19T+sQ9sAk
T6DOoAXDhF/W0frT4SYqj0eJpWvUL5cEDLlmBFMxhVxysDh+Ex5VxtfaJ8HFF10+4HSAUxy950OK
7Yb/7tS+tKPXpkfPWVWG77WiEko4NoqXhEXgy0SY6HSWBpHyAhbItq682B8NPs3wBwd7mLnDOUDe
95cWmD7Ri0UYmLuXJvrg9rGadEz2SeEkBH2xh1SoPwr29flW3FutOXnYsf79jwufbdHJ0LEG4qLQ
4rBxg0cor15kpi8NN1B3fjKn0mLXGxsMVfwf14EeEmRzljp72jXccm2ReAVp/iykNAA2hJbdHOB6
6f6GrZB/+wjl3/FErJQbHbia6RhPw5Us24C1nXeWLnwJS0Tszqk57MDYnqAGwWO92ZxmdqPAv2A+
RVswbRgyCEFz8CExnctz6e2yfX4oiZRuEufwANFjVIfqsqgzNCnYCbw2vjdZ4SLrPbpi4dzpYKxF
UD8VryvaIbYu1Kyjb752j281zESa0txRvPojlT+KYHwlEkpeM1Mh+slz2WDNrtfK2b6r3qqjBogi
oRDC5JvKSQT7ToKCJgvBweGh+U/LZAI34Y3JIK37xjO9dcytmkZjV4C4nWjmAsioZbUSYQck8vpn
JvuGYt7br9aG8sJtr6AYDMqLsIYKiMRrqizqLFg/Ur3PpT27qOLiIawc8N6EDtkQKcDQovV424TS
me789Ab0N5uR63ZHHr8eaaSQxHGotNIs3HG72VOQDwrCeC+BO3RuP6eCzIIva1JqBVR8Fq4ZEoib
WWRwVQELYvbNRPwXVGUIjruqOGu6tuT1Ff9krr1CZk4OZ9lP27T3rhbr3dCDQ6vjLF6HwD5MAgxJ
x8wGQwTWtvdRnGS6RiHmH9nQx8VXcJpnIYOkN5TcI0+UPIDAQzWoifjzDu7qIh8PaQ/j56hTOd6i
UL0UgAJjs0a5vDf92daY0yTNdXnxUAKkeAmkSyWuOjzkSa4WOaGzE4kEXIPkZ2D4rekrg/M/7+Mw
XeBwlbK9Me/+15UjqPSKu809VycIlE80C8ewEDJy5AZnGPDXaMNzhs9kZCGRBZZAqffHN8gQbUNP
Tvj5cZQr5zG527OGlpSL/PFIR5ZSLOtOkCYJiy7FdSGaPxgZS5dsHJArxoEJv0chzjl/G/qGvz7B
4LNwDiOQ2258mn7pDSWNdZn6wRiHaz+B3v482mWKRMD0qk9UewcnxYsCsiokdhkcrZYO4upa2M5F
vsZerhSM19IrQWPvmWgb1SPWBt4IXTGoasfaLRLRf481zGPwjnco4LMIf0pdU907UnMDnwnriPd5
3j1VLLueusKvYAbU5zTQWnSMJ0KEX8XOXvWDXZBnYCba2KbBm1QUTIxdhnK4fmAZsD6aUxmVi+SD
nNF9zneOV8aOvT9vsPkEFoEn3fK82vRArQ/EarI4EaoGT6G4uNrAfYVO4bpSN1zJzTGO8lPFswfm
L/UQDGmFeoEmaCQ68G2MOVoamDwkvCf4Q813/ELaEkofLu6g6LZ6nAS0vA+dd50r+omu5FTblCAo
q8gXtZ1xCkuVbTCtj1WKc0yHjSxMqXNStl9tmqjLzNgqxD8FqNWqcUw/FbYscd31Fb6I/sSE27Xs
DfKvxeMBht4WUfaODC7rzQNm9sEsJn9SdwYBbXCaKQnlM+b0PnxhL7T5NRpdqgacNRIOGosvXdGV
3EB9vN+vaj58m0tUmVRb1MHVtLry8gx4ODF23DgKsltUJftyskgiwJqwd2Oeh14xjVp19sPePhZk
T+/kbM6WachW3Vp/eUWkWDOWPJ7HnaGoKctAEN73bwNFkoYAu6tBXIQDw7qi85VH4TftTG1qBj3s
atUBnM8Y4m7gdtZgojq/se1mkviji5qUiUxllTlfdcn4JQz/rbfCZL9WunjkLYhjjBM8sL2a0UTO
b/6QZSdgG1GRsM0oRacIp+PBtxlZnWd+HBuq+ZMgoLKsuCOy5lsO2zctaHF8Z4YvvRa+ffbYHdau
8eqaxiIhVkUB8a6+6vuEd4pw7CfD+tbx9J/VGN+7jfvhS5AUR4hj4i86qAO0EHwaFdFtWTRAgjZT
vtzulB8qRvagoBvZihe7nA/VV38bBQHrsb/fPasPcNweUB0VuJ1NjFEwDjY07MIraOs2V8zYgeU+
nzi87GHcARZz24aXrm3ZnQu7U7AJFMmRPL5usAbIwSXpdTfE3Bw/2THtlUhi/i0txOwRdEmZigjt
bD+5xsZBPQSlqBakiDQKQRNJQ6SiSmO8GU7KxhRGCKZmhLO/vyNzygfHpK5jWO59vY8hUcQhUWnd
pkQU6q8+phaj70ganIgj2A81yoTTD6Ib7kKUdFvKRd8ol3+UpVE8B4X7+sF0FcQdcPnVrI9TKela
MHZaG/Q+Z0nuu/B4baSbkROvNfoD/fPnDSEOJCqWvzSkobDTDsxBEVtkzVolWyPcQ/50msthZYll
l2edXvXlDPM5Gp0wpvlR3dsT7M19Lf4pAj3qyVd0Z82yo6pilC+VbC8Fc3iY4iEP86GzzkY02i9Q
4OSpNrZexDn/TuJpqwvA16MsByT8v1Scm5Y1jL5FS8IcXHWrNKhEIH5FuZLbTzs9KJ04rGg7w2nk
wkAfVJCEnOnDiwWOZEFfmh5qCmtCLamf5W5Di1k9zdT2HL9U4PhYwWN86HWk+P21jQHE61NHNiWb
nM+9o5Pva23WgTXFUsOd1aRvVPhSjJHrel89D6hybHTm/Sfckap48wSX9YlzhETYzYRGDVVFN0Px
ulwgkkyftxFUBFAAqWp30m+EJeA3F4uLGCStWYSsSiaYdD8xE8h2xX53Dku49zMLyS8amypaDGUs
4UVoT2xABSTRFgu21JP7uhkEMOOLF1PrWCoTv8BIjn+zbdpz8N+/K6KZxM5N+rA56uunxquMmC/R
M5Fy7o0NKv3z8ls5+qcZy61gPOX/AJYAiRiR+ZLuUuThy77OAH2qPoDpI2JEBuIdbr1OVQzy+22N
dhgJbOqBgM7lm75IFQHKMabdsmA9fVpzPHvN+bcWl/Y6UD31aUqYKSx7K+Gk4nIeDNne+jBhl9Q8
BxMKKGknno8EkR1UwJ3a/WfIPHtx33hGeKJv2oFdHxHoMrZaCiZJtKcC8gC+ne61r5bz3xT4MNIX
ibfDRr1CyuK/jOmL1UeJPxA81ER80XFatLatD+vOv+2+d1UeuGX/hRESMBMGdAvZmtwM15rDcAi3
qjKzFt9ongrT42XHOfVwxMD12M92bCbPBshUCXvaJm3ndbYUhnkBcWSOFkcMV/D8KF0f4XNgWZGt
BKCKI/LAxRtle+Z6MuDnWvzAOC7tKn7oFjyV+FX/whwPtFvBntzehejwPI8cC0/qmKp84Ga3tdTO
Mm+ctdjUTMPffAD5ZZMYuXUfs42EFYJa+PDcT+pj/q9jhCeiLUO/BmlGgBWxM5TZQfgnNYWIZjrG
Mqu0zWM06rnU1vsJWNIRfxtLvyukM2L/DufHW0u3+YxHeuo8yo6fEQlNOmT0DxS2Rrz7uAV3E3BO
v2miN4ihhODzIJeJAaWb/5J+eqY7SOnbTCVGUYGyXTB4ECnloLROe8/aHUd4lcHnNtnhfpvSQZ7C
WFKRffQ62Au8zCwngLNh/VfD/8+NeXKFNg/fgq+eV72wu8cpo+qbdogbkfT5LEwAeP2DGl458eXO
69b03VR6ywW7nD0h3dEBS3qwOedXsl7y3MKgtmpcly9nPmlc0ujAaxBN8+bCU/IS0Vs/Yajx8E9g
gdYL7pGBPwp5GMQyWlPqDIpOw83SbE4HTBDGdy0WW5bjsvULc04dn8cTgyVMAZAt1OiYW/NrZQ5B
oiq52uCqXHMmA3DE/qsIVu8mgEJSJABREKuAzMQfCT7cv2HDkCw/Q+Cv1nOxYOcs+1oMiZ7M/+ft
hebruBiamyFnogoamk16+SS05bAYqJk+ajHAlSZZfOToAfCct94phIO6Ey9eeA6s/nV5HekaGGIt
C03k9gWCmeOlnTbl/EztFNrp2xhY+VUoNGdb7BPmXf6t3DsSahSs/ey1Nn4QIpUTdovkcDMUQ3RR
FZyzZ138q6OfubuIFcYjjhF+Q+TQYNQ5KW8Ni+qoYGw77cp49HYhuuud8FqjIHUu0Fmz2rf/by09
rKMZUsKxVsgWqBT93Un9FEUIT6p5YVh9etKxu4xfLNqjQ0FZdehKyF81GjL9c1y8Mh9u3lDgAd1j
caQpYEqK6qsuphCJbMPNkLxvGQx5fd/nBlPvjVCjwAP/un9rSH4+YP+rlVJYTACTz+2f8Jh0OWph
kgKvoiLLU8eagtRKk3OIYGsyht+liMoE36mMI2xgCE2Gj0MG4WQmiWprwB/bpdbmnDLWMInMpaLs
wIvSlPo5aMB1TpL/rID6+UvG+nQr9OI+l+JDXlBQNGEdjCCmU5io0FS7t5jTuRdmNPZPJ+LMqGPp
XhtfNrxub2+IYVYCtUpEfV8iKDxfYYEMDwXb+PVavBUDNc+t2TDMtYX8+aG8JxCn/wTlgwq81tyr
6tL1+xZJhMRJfeHZq07+CPlWaaLCnPxZg+OX5r3qHtUT+Y7/qwGzpV6hNgsNet8/E222KE48Zsop
mmrjp03k+XY2P/D5z3l22Yni6Fp06PFY1+IRLdevFqzmmBv9CMBbOlWurIgcuzCw/3F0pWZJd/HS
wc/AdNSwiDv2XH/WguVPDtcjB524iCU8QtPfWLl8x5meYVZfz0lKMRbMaK1stwcQ3mQe3Td4F1Cv
TtiVg2eDcmHLCWo6upQuXFjePPekueSNCDKFuvTETPM+i0HQQkWbKDwg3RSEVW+UjMeNHoeX6fCJ
/2YxT83jm1ClGMYvTQ+rJYkK8HSvS9vgewN6CH/Q8aNlsru8k5ezf9JJlDx8HCNecX5am9cU1KWk
Tp7YfgEBSuVbDkMOdIcIWhSyNefxOjzKisDO2C/kOZQQcO+OZdQhM8A4jOKB9u1p4tMHp3qZf1sN
7ZFzTzVzTjTIRaJcgAUavt70JPBZ5WSRX5MjgWFlj41S07YnbR8Moe3jlqcA/87mLmKV7bnZ7gd4
QEf7sZvx+8GioI93No2aN4RmTA7JbE8sApXpoWaHM4e9ef2U5Ty8XKxZ+JGtuDYzoVgFWgyri8fQ
edpcLsm5QlZSZmOfhP4aYnECxCchTwkliYSXA5HRDoJW/ZJsQ9LEZlJk52oNaBbhNNFURA0TZ5Ub
xVGaxyCPQHRmUZYi0jN3D823JdQDi8tmnsxsXdO/YdmpyaRubIAEu6M/y8xlfn4O0bl9NEVXV+U1
L283WfVs/JPB+6cIU4Jy0Yrs18q6yKtSVUHh3JDycmkEo3tdW0cLR8GbbaQTmO5jky1WX+hys4jC
cEQbypLpmP+GNTsuuFs4MpMJiY0GN+vZOWBFi/6j2lccoeArJpPrl9eeVEIMhW2jF2hT6JpXllOS
0nksAYKdiSxdWqu25G7SQuO5NU75n0jJtW+xT//bc93sPgqjrz1U7zrdmjymWJ4Fkc5+8j0eJQ+9
f/splqft/AupnVxPG96865cKj+ewHnSLCVmxTCVb4IU5cCutSBC4FykOMcaFmLCO7ijUO3uH7pDi
gByPBa5j9gSnOAjFyxJB7aN8WSorVC7f12DubQYMJNpYytorBUsF1LDdTwys4h6dcKipMGZnrNPj
LOEY593mO9nddglVc/9T7l1Z8eYV66e7iqmBN3iJQ4TLsHTrYXQvLQepIdBACjA5zB7z9V3Kkj3K
SrTGoj0ZUuPTSGSQ3s7r+fHUygKZRoLPQ5QYEz94L2Hegr3Toa2BHYJXWaYUuBLKopG3HXP5waqb
ONYXULSx4F9COMBFgHYTdURCpS7F+GKQclpvp/1njYtjdb8/Rv5Eay72xPkOawB+Fe/wb95zZ4dD
gbJJ+2KDSXvqQhyPLvoSNLqJlVr4kz8dChPZkI9sJaWlPOR+/IDGqRKPx9KqWdHYeN7bEEaQHi1C
BaGLiQ1OpWBQrfpjcWR++iPjSyx/cqVh3horYcq7dQD1flYMzbnnHbpxfHuEXh/sgyL7LjsEIH82
pQafanZTxQfX7L9YSQlDqGm3Ala5CJAnzS6MOQg/Q49zSBqNrFZT4go+nob0+1/ONS9csiXA+wce
gdSnVAcdLAVOOFqUhaLdGz6grkP9zaSW4Z5mQ18sLjpPrbDEEkQm7stuDk68XrArxBNyPcRbE3EI
DLRREpWBG8xL7dpPmhD/ZCQxNwnj5GqrZD/cpgvzq1I3lm7LNW9A+rY9c4OiwGC+xGe5B8rZJZUJ
0wKV2FQmc3GobYasGe7fyf1BU5naL8apGKHenM5QCds5ZoAg2Wji2a+TFdUk4F9o/xVJnHbGP9bu
fbLbPWcXZUjIM6ehAVA3OtihudeZgNDloH5wcbjz/00ekasj9+AEst0DA/N+uEimKf2CYKqjuDcu
wzQXDzMj8cnCo/yLPUGbSIa3Or/p8LXF9o+rSCvo8/WJgF4OhGp1yDPcxyvIdu0hOaAsEXsmeBQS
5G98gCNDDEa3/OdB11okuQb6UJ2wIw2bXEX71dPL1jZYlVK7SszGqgtTyzJ5CAu87rg/Yv9I1O/j
xCxc7APFGba00dpfM0h/pKOXdbzIjCFaPAAlEF6amP5CZdrviu/PDdOK6WGtc0zi777t64/raIhx
vGBNmoJnQcu3az96rzZKcd/hJv7qOG8zumAUJd16QFepvFEC/vC0RJNJQeA7XIarTT5tEsF5Zzg1
4rtBCsYg8ALCZR55xtp+fQnZS4CteskWYx+PHe3TA1fcsou3RfQBNa/81/V+oHM/iqFROEP+Ctk4
BQrHAeLDsPMTRtPmrV2n+SxKzQMbT8adx338fTLUEFvyzZtmx7PrOtbWf3NnqFz+lmlh9Y9XiAzC
CydXK7xhBw+FtV1LaboGAg1UJn3UoJhGQsOzTkvG9cD+9xOWFiOTwWCrOh8fTVJjiSEzBvnNU8HW
PXxGG4wMyah3CkINtfc9E5C9TIQwC2xI7WiNGgShQpJfXi7RIcas4PdD/ldurpXp7MyvYL/uTVNG
TCUmed8jJhr3NbpAwtwzUGEMDic9z3hlRY8qSmS2z9mCS+WSdf1lk/0dPKp7bFpIn9A5PyV2Xo69
LsWI+DoXqteSBnGJxQoBp0UmWnacJCtV2wAy6lMQIJpl3dJfiHsHGXZduzMPAAHu7AarAncqO665
cVqQQUr4GBd4d32nV/m/VzxR3U9lelg58w1K7K5nwSJx6EB6F2TMv8R2Ay56L5t8k59mOQAq5WHb
3aDTVpYUCvY22tvzAr0AlZHPYh65psVdQW3e/BcYeCWakbHAPq9qZmPgAZAcfejMqSgyG6eBjYlA
I2z3uQZn6xj5Di+yZAPPTfcyPOnaZsmy+KFTQ7SHy/hn0E8rBEeKefPqSUIWktV5iTNNbAzERDj+
qblefuY5+wyzCHofEHCO9M85mg8L7IO8uT3cEDgq7YD1oYir5VwJ9GuXqefbkHyUOmKQ8xo3SWkn
noozCCiAuegUdvz5jKBITqSErv1Ho1AOIKNDWxGeWJ4Dh4Y6pCic1/yoms3ogxux8mNned3euVta
DaDrFLHiEjFmwJrGhxVVrtxiRtTWGXCPk52J14teYVyc7/fgk29P+eJBD3/JYoFYlD5AOJ9MytGe
foDzzXtyeSi5PKv75PfwfJHcqkzrknCyoGVm01aLQpAkwAMuQC2oYT6Y1/YolcovuQVNNuS+6wzq
0N2X9xJaf0hFj8ZjcjnCYVtmhVNSDX6rUGycU1xMONpgejuVhPGcSs2vfxEhFylbrf5jXRXGg6O0
8+CE/0XgBbPV3Dz4IIw+YzUAL6+Bbl+bqohXa1UielV+NbHkFBlBxxH1UYdMjDc2QjkcuWd7LrPr
R1doJDZm4Id5jgP7RA4NGGG9RacS/iqkF6xd/+LFwzNUAIaFD6XFwr2fj0AD39TfcdwjdUVs2ur8
fiH9E9YegBeVOY+3ybfNC+b3U+zixTk58mguJQSdZar7t9AF0GvBlNtkD+HTcmhQpAst/QzIaneq
O1YrxcP5cuEEmvbGncnUlpIF0IyxX/TuAR/OdxdEUw0GeiycUhuagLVMxfv34aJlMguwQUfF1bc4
kmRzy2i2FQFxuLqN9QwBhE5NuFhGb9yMW5XR6YW7iSHLvqE4X5G7/NzY4FNBEC2Co9whWfs7TRLT
EmIfTrhzZ8ZV4bTNP7H8V0OoCDGxHOV/cPk2WWk32A0kqD2iv0dgNyyoq8IMWv38Gee6MMKnDpXs
VgiP39+gguPuRAzLH6iwW4Opx809+0dOMOlPHcu69NaP1prmvXGn6LN5I7+hYzLMuLQmWMqhLmZ3
hRLE8vsuIX5QPaIvcapqb0K2WXFdI9+ibvH1JfEH6NP/2k5glAEPTbDko5yeYYp2yT0qsRxVDIsT
hqlXOXg3vKNYAKa7VPK/clXNnpZbpDqP5NEW+BZ3gfG972e2t/OxdQKyqYhl2rcDs1/InTbhQsY/
ExawNYpM5ky26glEiRyh1oUGIiv3uY+KqeB32EjG2A94SgHOORf+Ytur9Z87CT6Lq91+WHlxynA/
nc/WsUpUqDZTMrWuBAHJ59roRAWilzc+njQgjat2Od3bPy6DKAOGcFRbN1JKBuwYO8wucMAmkT7O
OU/gf4l3c8RV93dPtH+KmTLX7vykhaQML+J5w5+d3C8BMHgtnI0khYk7z6fzoRMk5TooSC5/RKFT
o2uc7VZXNuZTxmoP9TEY9MA8S6N220Xx+o4OtLe2D3dNWsyBNiefXl2IQyRhSwCVpU85SyTQ9buS
3yb8nNQQPhPJd0t3z6GF109H/RvfMQrRGELJWenzA/iD3ODxRzmSE3fMpish+veemSPShWhhejJh
0cZp0IjtieMtPxjRUx9EPeHXORBRFNm6TSxixoKTSydGkFYLjxD1D+UQp6CD64cFP8QVSyB4uyab
g8F78iv5sqfZgMQfyl5+W4DkXMbP8Q4C9LUfEELDiHfzX4gXdGzMOKRiWRFwHy91vP8lRBbGG/Dt
JrDiiXSB0WqeDRobPJAqigzgYZl/07eUBtxsVudVmKZxEiA7R0oaOkjtshMqUUAJ7LsBHTYkuiEp
jmpkQx6JyqA/w5CtCpLKh3VnqEnke9cFC4UuLteClHWiUe7gIDM/0WgsmbxcfBNP/y/aCmNoNdLD
2c8lH9ixBGHGq7qcRPQEHcFT5oT7s51AKZGdlpcNJWSj6M04JSpiBV07FwYnhPvRjniSyObuAYZf
cB0JjM/bTmoA/v29wLMhFfnHLrA7NmBangOavE4bbfrS9g+9MXeRHwwLXApAD8x4SiHykq6xCqXz
1TKcUviOwydZ5ZFnc/66km8B/2t8KOUteLJnGR6ZSb+lwluLUzbrbuX+f9twtiaK/cQjoeU1YGOG
rl050TpRpculxMIU2BTxH4Q7tH8SkVPfwx/W600EepAIsqDFOfnFkiO3K9KzUhtrUH4wNmUvLygK
uN8Ypv9jR6ZHvobJJ+YU9le+vcWKD1wpE5hEJ5H+cx91qT7aOUpbcB3UmXLT4sO60Nkn6TiXlK5w
1EnOtzByhU2i0q8INravs0Eos0J4piLEno6BrIQKwzZD8sEBE6J+Ir+HYqfS/Cyjt3+2I1ce53Oc
LiTR8VYdOO1jdo5PFWjcugwKxf1oe90ff3kvrM1p4sQdhLNHGtL9mRbNscHk2lFWJZdq3EJQBRsL
OW6SsO+OYdx/RL803tZ8bK7rKIAkl8iJjpP+zv+z+/hwz+fzcFcbml+Hdxdu0sS/oEla2Ua+YreT
a56nx8jF2cTp3j053BG6O+5esUEUgfRlWPJl+ATN+qIQivaPT/uKuOIrnc1zxWK03Jf08LdiWpI4
H7kE1bYIuUBFolvlxm7on3H+hXdUvA6aQqZgpngH8Y6/dF/BPq37j+ih0IRsOkxZY3SR0iZ1vBuw
iKlZ2Sqxn4YcLeCOZP/2aNGlcpA1nPaaLFw4OtgkBosEGhy7ncEJIAyDfEhlZDhA7thXi2eDUKgh
JOMAB57ar4W2IsMpkv5EuEjbsiT9TnlPzutzbbnkSxRWS8zclDe9nf9JS1zOdHuxYvzjDRSA43wX
gHfsxxKeV5M2v8n1QgqRDKHPzX3gxEHyMhdSKxsc/HdVZz663ndTmZ1mT37xO3BLW50H/OS90On6
esl8nUpfWEtQmHB/DT0YARXOMIIocVMIVdNPP+z0tnmWLCdg6dZasl43FpVeTRh3IUvPV1Qn7w0O
7OhjuSamdOVCjErwrbvNklEGDFr/7/vlGgQlLImb3VcCumKoSMmXvGceEYKxD0CiSCuuk8rOld+g
I6VXtQaG2ZsS0EQ8C7oBmg9IuXUfTJqNewfeUaiaDjajox0iMbjr4YSLMX+VGAmqE1uEU8S6PTW/
4Cs5umktiueiNkU1vEEgq0niKlCypyrtcOTwjbW1JFKd4fCSnrG3XEVf8SXQorqg/dvQE5T9Yra0
IPqSb21fZWiKODJ71NIkMA7zj2NOfIaQH1tD4/r2tbRa//Dv0AVG0uqa6yuTyDlQEmvbTMSQwo+3
iEI9fmvMUc3Snz2GzCmM7nGAmSwcAy6rswE+RZku1C2qQ+jzX/JfmIXXCCSo+ulZ9m9sm6XTW2Py
1j+oAiLgrjBh7Wnp5lGBP/pGBLhm2YIeLz1Xukf7/u/zRx/+ytE8kMlqO5GacS2dcoxL7qfej5eX
IOt8NvpiejxIH5YkoRf6URMCHL11O0fWLEme5wmViOuB0+ZagC5jcZwW1fUK4/KAyjWfEyDJSiMM
o0IF3zAmbq6pAuYM2rNybvM/U8/8OHXEmSiCQ3gWh/h7m5kzNSxxwdI109yXTeGWkXheU06EYj2J
fBOoGaNUmvkLLJhVgSMVfcOGcKRpCOaNlzfCGEtufnKtf5gsz4TeWX04KXb/SAc9VESUyK1QyQUT
S7rUhSGw79ZC+EdF54pXvg2UAd+1OSHtGihNKDS4u4JGCzog04oCmbdJrJCM4IguW5fhkq5hWLb/
eNdlhQFNuALR0RAtH3m34O8vfIltdfIAAYBN4VgMh6lAmNpZA3Y9p0eQzQunLv/QJmPDCEt8YRR2
z9ESz/LcH8NHClhl7Wl0DXV7HPgr5qI1wPWM+kos64ZKgmuWZCd1L7CEP+rtdj0cwcD8L36wlv7x
uqXh/TRrR9Uy1kLAZJ4eVsrXXPUrO4yqj9wdMZg3fLxk6T9ekcDlnxLxRSVVrdziXJcZl5/bQAPA
ZhkQfHCNj8dW+MkjGc/33Pxk3XsK59ae5QQUWXqvtpuxUd5RXUbCNhpS2n0In3in4kPOMORfgwKc
PuVBYxDmSzZk5J8bqDdyxHiJqoduoEQ0aZ+R+o+XYsO6iRw6/mTjyA/O1d+/GyEj5ybqzXtxfEnR
WVkl0RSvQ3Yda2J0lceo21w/JXXlsyGKpu5LhDfDWODCM4jUYtgWI+a/8EQpkzf+8msgk8u3GNqp
OM7AG2/Dr61d/RsTW58PvzO4GG85cRr4cq0wVg5IhojAJltrEvCopFFGSZyhuYLTAdmkNMV911kC
q6o8PZVIvwZHTA0DEFTVBL5mzu6FdTc+DtYySqEuzW1AqDS/G3c9nxj3snjIa473KF2bui7PBDZF
mjpkcpoaIB5BJZScMDVyOpzy+OxhxuV6B+bFL0c4wGxv+PpZIr4swOJoi8hsQ7Sr4AJ4KuJlYnEP
SgNJjzMQbbGhzlPqFyIgfhmIFlsvk4H34CwkPOG3kfABjReXFQZIj4J85Fep7cyDbhyhpYAoJzCy
IA/SDjQ0wD/Ht/zVVkiBqE9mL9vJOP+8VLyLLwc1lfflo1mDd7JeDLAwXSffpn3FelO2H/8tG62x
Zso3lor2psv8nKS0W8ueO05YkRpcIO1ct6cuCcNUwLn6ohI//qpvOfrXLFDRH5EJ1rU23eik/cPj
kskWFzrbbc5Hx/HtWWmRwuvtPoDueVIvbsJL+QkBVAuGzIzT6oKWcRQQZYdpFOWS4w4w2oIbuElD
KiVwXn17IoU3pCGnygfPgHKeBBt+EuhhUrUy986bSc9lxHofnBDp3sQKvyvm2pxgpa61xY6ExYuJ
sRZ1lcrXb+NIYAVQu61v1lo0JMnd8JB3MelAqGVvEiz1i908bH+XDuJiw/2L4ohlgSGwegVxkphu
4vdtJAwFb7KRDkSO+temFv1S2vQukxf3LFwfi0N2WYgOKkovAq75dFzM/E1LKSelylFdi2xm8SXL
mFkg+IgeAuHYf+kZ7T4hnxcsb+EhTdImsusIel6L3/BWid2PtmuointWSrJcNLtS5WcFrKD/MAZb
evGy9C8ZLc3uvUia3tXbq27HXsv8wEL6MgRXixV/5iJfnvysF5UBxdVJIn903nSgOUk+mWgHEH0Z
u6jEfMfv6KOk8haWagw86BMLaRwYkkZQT8lOM8dTYV/OVUGb0XP6QWxnNk3JxnoCu7vkK0dzQtD3
L8YKN9Cs/sqlUmdkmlptqpRfuPbO68XCd467CsBFxUNjHcjsyBn2rrJHT4I/z5cq6Zi6U+DoiHDl
Foc2FI6R8bCLcIBo1A3lWSA3KAD6Vtv3Bhx+uNaGCHLnH4HGhPVbCAtM0v2NvDEeST3bEtBzrf6I
jUGFlBYEAzj5XW/ZuVN4NYJwUwEKxMQsmB1wgW6AAaQJniUJPPNX0n3fI/vACnCf1fpqQ6gzIx+z
Friv8PsauUEyOGa5+mlVZrtxkVK/tJ1+8DJwj+kTlk8FKc4254fq4mt01217ppV4Y6VvVDuhlBEA
pzFVgP9xas/UH+Zn4G8mskq0GdOU6adnUKgqXJbOU2MwKJkq/MmbvFyeTt2Uvj5RsZa4GoRnefzD
wDfejBNWqkuFi8tsCKx9XlQ38/+QBYQ5xlFmxbsaWQzEDWQccYhW4rQ13r1+YxbRaJXfodDl9kgD
USBD5HzsbIwjNiZkdgjeh/uf844jNGgmynK+8Fjb/o1uTtZWiSHQjiTjdIU/K4k1169Nmt5EtC8K
THrgeiv0YRpQyOb0E/ksElWhCI68xO/Kjb0F2bJGZ3FY7PcX3fLIbBDabA6G8/bIlUcW9q70qAnO
KCL0vWJmNWeTofbEiGjqmqrYzxD4rmvUreopM5QJ6euJrpm14JT/I6SRdCJOeyhG2gPZrGAwzth3
ekB1Z+fCc6j5/D9fqw16i9/FyNm+pp1sDJi4Npx+fwG/ibpxn0wP3QHlCCGlENiuXIaMGCMvz6WA
sSZBLK0D/O/w1l1TZ2gDUTrDQhZ2zNBAlcdNNwzgZLTlEfbakXROhGz3xdEOXjPDsFpv5XGSYu/o
HCq4deGxiEl9F+4ThS03ELSZTkGE1r1Pq749O3vBJeOHUcVC9h0O7qGVghVkjJWJ36KmZTJ2a9Uv
OZHGwj7Ok7W8JW0IQ2hik0YgfF4Q5OFeBU5tMnu/1apL2HnqatTAhbGYb7z+QbDnedMvP2/QwnKi
lhHhasbEv10QtzVIXvnRbXCNTkn4dWgfjR68NLtxcFwwXMzZ+1wHqtHsVLKI7i1xbP/W8fecovhW
OVxVNIJcqGM16nqZs3mwgBnQscq/JmLshl3MX5jK+Q5VrVeKiRLI+U4toHp79bzK7PYgNVRnvqtZ
pi/da7A0HNeCnhhHcTa7/+ZD2vRIFEes8fe2zXf6a9oHlKt9ydFmOa7iVP3oeYZpFjxskc8IyOXv
WtfeVCacSYTZ+yV6UxORMFm1ZKwV9KcgqcvlrGoQtdf/p/45orrNjbsbWQP7g0LfwnmOnGmNDdHh
moVd1EvM2iidSvTpIx+dWBKgDQljgzInm7ms3aIh5rFLlL9+tDGh1BX8cswXshvP2PFMprQ7UmZa
Fv/x1JLPJYTtNoSQUBuYK5wfa8a8XBpaaMEP4gJmvOKudFx8gO/+Sdxl571mhfq0V06/DjKJGF4f
+Q2P51DSZgoTauo0YH2Ce86UodVh1RHTl5oS7zAOXjDSQ7RxLLpYBHiwo4eTT8apLElUzKVqiRKn
96ST6Lw6L2egHiNTEQz1EWIkJSrKWtOsQkmsrQMs7pVqDAJflBiTq2S92Cwj6nTcISgo9iPYqxon
v86NcaiYiXX+tIYvDUfSHHPYzi4N9ZPZ+z5fLJEgTEx242f/gmTn4myQVebT8hBJLlDof9tQsEwl
RpsGuM+w0hD6BylofYgUpnBE2357VTMPLAqcSY+aghSJHkUXpsarcP9jqT5wwGuM4gNfAcXLQCKW
amnN3+Lrx75Aae8bTBbQH+EVOXhkcpNnc042J+9TuqLyZ/uZa8dSN3CYJfifrGvbu2D9fC231QGR
yNLY4PvA4S9y+50VxQOR2sxRB69D5cybpdHsH3doiiNGgBr6T0erNxvx1Nl0eP/roQm0R3UrkJdT
vouW7f/Z2/hqfvgL5aPDNfdJ/QMC5AkJKDq4VpAOgvouh0KmsR8JrOYSNQp269M09K/JRsk0KAWu
pNUdBLhcKN4kjnvzQVcN7nOoLBJvTf1epFO6hgsjsq2GL6Xdr7vTBONKP/NdaY5YgXIemZI2lyPW
7qSpNHSqgarbh8wCdMZcsoEvbg0epM1luRAzdEZgeEs1+WgKwZxcCSmE1IpoNfjEvjL6aq5EFygw
FhrjFLTwgn53DqhrvIpXfFej1KtMwe58uomN2z/gqA9j3ixIk/JTwh0hxk1RX+AxhBsGJVgNVtVc
JmF+TosU0ckyCScVZf9Q7ZgeSqmHnUscpyPdPDzr6ibxMuFTYldkbKX38zdkS3SmKLVp0NNwux1h
ClTOrDgkNLU+/tKUJLlkytMEHpIrXgE4WmB2d5YElUy3zKC/86dFLXyLYYLfWmHwgq4GdF/0xQUT
WmgUDFgNKks4jGpeXN+dihMsxjGyuzrDW4nJ4IJCZBpV+D3ZXwJmHW1ymrAP/GVY+Je9OymjqNYb
Q8+ad111LzOoTNzaX4W3IQh+M9VYwvas1DxHtqvoAdqHTQ3GAQ2llGM6ncxPt3oEpW5/d5Z4s2Xc
01A86I+70SBgLXUZCBUDKVV2/v5d0OOFchj9ip/QPNLva40ZnXg8FypXR8XHc9UXaqjJp90lflHK
amTAySkYN2CTQnMSeI45c3uH0si7pC1ezrldps5Tk4zFT3188lFtt38JH7OcebAOj2pUUzFgmD/8
gP07hzYBU4r4t+QHR+Ym0SfN5H30RLVfI5xjfpXOxMeCM0nVI7MaQibrRIbVxLueesuECm4z54ha
t3D77HaDdgqZgmlWPp/dbFaYN12UWtok52p2o2V1PatTqJcouy+QcJ9G04bmkDEGStfXD5rTBqsL
Z6qwakSDNxw9WXEWGPzaBQAL7fgs9/14UnZN62FpTQoS62eoOkYjpZ0/olWEsw5gYckaH0cqBWRW
PCcPeBra9u/o6I/fLdgoDqaVirL0f7VhRbjzV506WoAv+XJjqhnMKVEdavKSVU4j7t0HD/BNpGhI
4Qqqlz3iy+cplwsyB7azlF5N8LcMbwBx70r2/FSMQS/+NORxX6IC0fJU4qMnakyih5rZKIfvkl/c
sovZKW4ybu2feKzcqpoAqXIHWq/4yjl07ixJo/f/O2hDrbW5XlqA7u1bvRxAemYKjaMFhtX7KuQ6
iDjT79XrqHFKhBP+JvsGEn4v3DUPilD746Pbf7mw77D4Pl/Pg8HW/be5lDksI5GTzXi1hK5G2n/U
/1q2Cu7QUyr3f47+fN9xWfTCzUjGzOUg4/6LwoviReek+ZeOnNOKB+MFNOQJqqJgogECXQqJzjAC
vc/Ziiq7TMhAJHptAn48leuVVrKz/TWDVXkrwEgfgAIQUU0SbFtKF8m7ZvNfm1KHeFbaxfIIaw8x
PAHeKjdi6ss8A1evJhy8l7eI7slHSmOXqSWYa1cHEhnUbOvOSrlH01paiUKYlGjdcRs4KIZJ2j87
Xpn7iMZUSjP3gdhcoZ2M0AyTE5Yg+NthemmFcO9TLhGRXcdjvC7ZFkA09ae8sa7UIh8ieNksfsmX
sA+USDSW7d9j6DsnQ4K7um4Bl//F1xdiQMusqMV2YSzbH2pPfrJ8Krm4f4wyMEcskJ+2YVJLrp8Z
ZW9y4OrceCoHweyKkd8QN3NxkQmxE+cucldTtGwXsiZGGpnhxQFzApobwcwz0kq1jTSOmWDibYn5
XHmDyutU9/ZSLiWrzo7pY+w82wjY5h8wEzkH0h59fANrVePubbnhC6fuytdh5LIy+pOjsl263mmZ
E5q/j/L1Zz8xUECBY+CsG85bBMvrc8CVoMbR5YpVsTNxscA/DZy/bsCD7fuxWW1aJWk/iM2EPI6S
YvUTRUAYXJkt4rT5hPbv90GCGoUo7GsKf27li9mc00HZjtIDU4tCr+1XC284QsgT1CNZhede/2ci
BiBwCNEUr8Bx0/xxnaTs0NnU50DCEiw/9FynLsx599blYlPh8tXGUqkzIdLSl657GM+f4v2+JeZK
B4dgNbDvOxubo22ZiuK8hjKO09IGLoleAtmD4uAp8Fl0PmB7ROpDpdbDEdi61QrbApfyXtltALrL
3DnpO+3qhB2Qtvy1WC//wD0Pzt1ScX15lGU9296Tj/E6lxovlPAn2DsI6Hz02Fd0i9JRiBKpdjvE
LJ2QwiYSh/NeM1SxdCwlqu134Fw9wOwae/sLyFiDpkz904WaZBo7auXUgNF/95Ntk4P5jKZVjfsZ
TUvgE1tmhUVe5LJnmsE/JKvhw8K3WBO2qYZ19pO8+ig0u2Qw7uNgWuJfHD3Ov5UpNLZ6cMFCm0ch
j8QqHVWkVF1YWfPXVgSCyOZ1XPC03nhJn8cQtBI5TvUVdnPRE1MmmDcQvLjdZOB8tyTBIs++wWjG
UPHHDTT63Cn3chiBhO6E3YCyV8Tg4r+sJtQl7+kRE6OKZlfoLDVAlCH+Qm/C5eE8rWecj8WBI2Gq
kOUkPjgAl8vqoJyZ/Bx/F2bZTXjgwCHKi7Q3ONPOUl81a2O/7PQ3B0phPtsB1wJWL8yY0Xk1iWcu
je9fG2vym89pmBBao4Y2g7/LYucZ2fyjlSOO5S2Y9xYZJ07o7SSb24QgTTzATvDbUPauN9qFO1EG
8T/tIfPiZ2OpXI8h3emL0JqIU0r76hrQOwVIh76GVhygplz2+4vwAa5i3yRfBwqIvDyvXseKlKkG
I73SOKL7PoEoWyWqRQk3SPYzczpoirB096sBkIwXZPgGg90NQ8lqhujk+g0TIqzzG2BbKFDC3xm2
8yTDoi4RJWUX2AXLNWAm8v120Y4p6pTpqP2paFGxZAXPLnbQye0BRkdl16ZdBB+iwdCZFv/bbqhQ
3LeR1Rqt6cRFjlsMBZLqSoEJa2fbGgf1CoRHeW5J1uipVACOujCQ/m8U+HQFitxdfXWEEeJZoQmR
wekS91g35RFsL9ensUtdi57ctGn3AastYseuFSWMVlxaRxGo6aESgR4Faf9ENbl1L6AzUoz4BsFA
/E9e1PKWcAxgOGcfFb65IHA98RMHM9m+HpYPPzTOMsuZ7b1g5su3pWzz0BH9usMiTaj2npoi6bbC
IXBdz8s/fMrfEVJPjOBViUgL4Ymbc3x5BvgIH8emWk3PxDrPWEhQWAxOdf+fbVJ75Z7CGczDf6TD
UmA5gmfvg8J4vu37eYYU4HLgzyNrBvdB5SSelu25yS+fU+6XOrZxfkMHJoYJu3Nc/eqavmPWTw3f
qoR0C5qzy8h5Ue3okzHMpXxpV5Rtnt2gt1fsd/dY4k6IQJ2dtx7V1EUF2S14F1eqr2j7u4eLrO56
iX6MLumLTWeKthKEEkGx/XhFSCDbrXHti/Ped/+6WDm/7ASIF7NjIWWZJdQ4oynuzp2NvA5ya6w+
+UHnNH6TP9SfXM0xE5kGCamx/j8xm2XLoiM48zP8dconVccKkirb+0DwSkSvYZ8VQ91XcYKBIw7C
Oa4nFjZ65rP/AaIQmDET4OJn86dr0ISpDjptXON0T/NzyDNDG4vscVQClBBBrP/suRW1xaQcAcbg
51li6OqkZifCV/PSiTrJ6i+0UB1DCpS7yLM0hOut/KKLYwQ7jlaIil/ougxj0fxmJuoSTP3uNJf6
dvF1bkRl1ccoZ3WQ0sQWBTyGcW1AEbDQUKS8nCu7QV8wzTXlkz/gNxuia+oQzCHqqztdvt3zI6TW
ii3LVNvL3LczMYYPusWhbtNXV1/RUCR5mf1qLlh7EkhQdZhxPZTheHAKZoVWYAcN7JGOPjrcXmA0
Q0n+jCvXgXw/74J0ZrDAeb2f91iEMXi55UYp8xmbaflxwCiw0kVRuZ3DemkmVUd17rNLBEjbnzr1
yGpwfZBOaBIo12mWlpPLRc5c6fntneQEE2OxHal6qQKe3+3wOGPQPeVRaSA736DX8O5TNS8HwiB0
WqAS1fXTCjp/zcA2ulUhF+8HfFDxYD+r1eNOi0HbfDVSuxhidFPpbU6l5oDXD2FpPrUgRjoNWYRI
IwrrDFYwxr8JmorTdsyzsv7Qq5jhanpeHMPQmxhZMW8J0rbJxgEMMz1viqUh/+jPkDTJw6Sdbbeo
LVLAEHOVd35ApDfBC2pBLPemuCmV4CL9j5zMrYyFPenBc8DGfg11GtKZpKum2vJcArx6pevUTvx1
RqIfXhQ3/GGZBLg95CeKsufDIG89jhqrN7yB9rUIlBKDTHmUjvJNGa3I2KxMY95LvJP1UtFPizn3
I8HzM98Q3AgRoXRzIZZFYV9fq5EN0tupyz9u0Gs9Fsm1LnpCMo7KBzGhZGvEF/d7w8gSX/WUYnN9
So0q2f8IaQay3D2o9bA74N8k8ybTlRx+nUgacAT43F/mpxQDlEviQXe0luiDQ9rb36WuKoQ+GlNZ
3zYEj28k9SPH5YRvbFDf/jO/7B0UHE5sFQUReh58plsWSdoh/A1OMu8N4wM+KE8eADMmk8h43slY
aSBBK3komNPSnU9qoVggsOTUEGzC7ldz3YoTzt7yEeiTmauNflIpYQ2Ug3ZP3Mwa0WC3EBId8Okb
oMe21ZaTPbox14mnBVCPyvfA2Frg/FCY/ksyXshYtBPhK5P2k4hUKYVD+ZrqDy/ELqcbcWM5LTEW
rj/P9JWMvsseiAHezxhFBvGVA1xyGrfaPUeydvnJUChF6jPvH0oxtIOE5cAdOD8llPGG4VWIZTX4
fPKL2NcK7lDXm0eEEPKULoQ8JhC6YkZWS2JzJmysfLTW7gd3c3ZqClmForcBSEAtLfqCGVpBsB1u
rsgMfJ25SFgIEBbzxr5CxbuV1LswKTykAOYL+9AchZ1aY4DiVXaukobHBAiU9CUvwG6DudHf41Tl
mETnhfvtlh6MT7+sKpQ5tVHXnOlNGnSh6q5EMz0nuVn1mfSpuKYi0fGaEPmeCb1UABVB2WYrs8st
Sm5tD/St/IpTPvpdFoVFJw1ElyYDK8ApSrjG8rvqZhRo5hTGbtRPtes2iCbwU7iTCPx7MvpczOli
xCO75MCWcaZt6ZKQjVDyYSWbX3yapdduVyqX+7xqawgyVJfBYHr1RN7GjU2zUitIz6j24KcETcUX
2+nogBV9bopNrShAL0bEmjTzSHwJqS4Mzy4KBEfqt5SE1J3F5pqPrbtlqCRLf7+3lyeZjPYlKh82
Yrpk7mtP/k91LvNJVA6vl01zIgwPefKlDO0E/6QpsxoNRHO0OBRRcGH88CuxalZyLrnN5BT2sPHi
mJyijvkfI3cvkghgspcNf7Vby4xCTG0DvJNbO497/akcUmU2NvtApgJQUoAOrIxg+++dil2KnQ1H
fp2aN4f6tpQwUTzdvugLoNYTlKPvSTYAl5QHY7okBNk5kQFm5HeO8F5vdefGvpt5mgfg46fuCMFP
nkg5Y5DGyqXamyNBguyU0joPOiVaWrHtiYnhnZN/+XcUU6gv52GGNS6VMrD+vWrLumyMLrPIE8Xu
TPdbVsiJuvz9Fxz5ifKKOVbPn3Z0KkMpjSDUgzCttcyur7jQ8QTaq36nyJGm5bJccIokTYzo9yKb
HeX712ZfkVODSfq+96+8DhF+meUZV8TPJ8lmjXHcdUEkXFpHJtqK5ZhNXcrOCJaQk92/2D3uo6cl
d3XoE3Af04QUFbsuniW6fL6/EEIkcJgW+h9b+dl00LhfvL7SOqnLQhsPYL8GcvcvcT8xd51hDnWV
JEerXV4dN7BwfRQVOxk1RbazEuplHCFSraGMPY7zixpn5hnuZH6V7oZjbYTa/0SgYVSxvfiIir3K
k1ic8zVjez9gV4TZ5DcGvxSjd579Qpg6/cFYRs2vdN55+h5ekuFWeONmrvPnud2ncR+s8X01hrNh
KofesOc/2LkV3EYJIMxDzMzDC9fDynSK0h7CQhXu2pZpZd7Q013VjSv/DJR+1T+Dx1+uSa83e4LA
fxvsn5ZqIy1F8L6eUUUdELH0USUpGJLbuDFES1lkBuhNeINl8VunliILzc0/F5om/Wg4T4SmWtXn
ng+Rbo0857G+5Wbe0xSr/BdLoctzbpJl0HJHyM4T2asFqMjzfCszyQDK1MtGZM9B1FAllfwUIXBM
xOkMTEuPgDPqRlIfxW9QMHfCPWgpk2AFFESjmM3VPlZtLZF5vH+fgmjPfnrKDuFUbzI2lAUflKFG
u+mSTEiGjj93gTX+hxNBdebcOCJMrqbl7ULTrx/hXe9HxKbDg9CcBnQesP2dUxcRunnz1kacHdbn
wCCAtAUdpy+uoGYPLAvidLO4HEDqzW3GSSK+V4p1MTFX7YgMhLu1d8yQqspI5NWiYtlU34QWqn7U
bae/72H5WsbgvvcUasMqTKgF8lJzjpp/GbJ2hfvggRsuiZgOd5Gm9R28IDZqPrc4NG285n6Z3RSx
JPUmOTLkgmjC/M0vq80LJn5jKw7PVnxgdqq19sbJgzBaL24xGarrTUVUNqwEGg7b5AZS3K5VlL6L
VmzGl6CkReYmlKVoxaEmy0IqNoOVuuGS+UkD5pnf6wNnkH/tGhE/4ejPDkfO+kfk7RhqU62MvTQx
DJQXoI3Lj9tt7OMVt+C++dRq/vm90GZj3iqt8UCDt3cxU+yn8eKq/yA7H91d8qqZSqPzYyvTPfWb
mx15DY1GqGh99oxalRNWz1qELuLDyNupnyI5MapGTbd1DtrzcGqotcgVWGoCiMzF5wwZU3sCU+qq
iG0H5TuTkyKZToWZ4G5m5OS2RPjpjGncpLcoi51H9d4MSKmTS4XfeBkTlrjjzVSs+iT6gxGxKtWI
6P5K5ypEVQzsEdRPTUEvBgexu686sB6x1LfL09xeIetzGD+Ei63EcQczb+4jmTjlGBdIBcGsbpXQ
aM+Umafz9CvhyLTeB2O77bNLx6U/k4+vRySX2KehpWTlpm6vVO+x6niRiF8CQf40VF5MB4IZm5I0
wA4UWniOlzU2yaK9w3aPYH+eK0KiFWmUxJs6yLUIj04u5xBBl3d1p53QvWmaP6Zj7jDJkiEzLMdG
UoZENbbu3i5rSKcUDMXD64vQi0ylfr0U+WAcjXw+uLMGwPjI7VnM3suB5iA7N/LIjkQ02qgIkiQJ
jIG0nxdDVDr6I4HroZqbLUEkzHFE5Y77g77yfvqBRtl1/JV1cimxOMvUhsW9qUGC+xq0XWOAk1bp
SPGu5egTH7iuoum4meKg69exLXyPBDiEVp3/us46sK7kfYhdKdKY4DodkVRbPSarxnoL5lrFfCmm
zQWXeMHGKqKzWMVzo0cyEQ/Srvm0wp5d5PKUo4uiHJsmSe5IiEv0/UHBM4Qrom9xbnrWAYnw2Mge
NoEa2hOBatCesZV5rBnrzdXjX69PBjCTNc7KYcxq/erUToo9JW1bS1T2Ma4zE6HGDtE7pQuVIgcf
U3lt28DtKrLNRgcFfv2h02sNLF8BylOabVCkATuOkHzA0YNtilSuqHE73sW+hCf8173X58K4QMgD
X9vVrcqIuibyxaOD+HvipU+kjznICzx9xHeJ6l06QDaD9bwTcv/0X9uXRvQjjzIVWh0zSSnI5BhT
qKGAJIaPfIqYMVHckhhP1isfzPw1zhlarFMqVKQFX9unuyVotlqJ3oin2TqItb5+9f5s3rRCwBy0
2jUwQhq01hHLcFgjWCZCYWSa7KuC83KyQGEgpFBntQ0wIXUETO1mUji2lxjL5Me7ecwFMC7wBJNU
/jAKSR5d9BNCRnQMUZFvitxrBUqcR0QKPr2/JwAPtPXuGRlm36hcSRsLDbYXaMB5SQYoGL5q4Jlv
8S9getkPrY8W8y+PM73UUD+sEihfhynHhKlAJDCUsDEemjWswW+lwh/iAiL3vuqz8ghK4x2yo2VN
zqYNRCuWVW4emCStg+zX9IEG7gzZwC4WU4nFMwzlTGPnoYBQvgOpedmK8NcOwpfriX6qFXTqUqb2
Lg08LpwEI2rxR6sfxJXIkwWf5FAdgp9YJKyzZ9MRKKSIxtd2gyYycpsi+pGQ89ZSUNopERghRIwW
rGgxVZUcnZxLDu2dNzkZc2BqtxXl30n/yZlarxihMK70f6H4HZ7WwQZVLmEKcWFNZ65VaOI/O+Oe
RdjM7FvC/VyBgnPLG9UnhKdxR89hfLIlzhBD23FdwhQDXyTywiSrm3tMciSco4uquTupsIDZ82/6
fUe2tgWbh2R2mv0lK7mAP7Y1VnOEsu0O2vKwuFWCa/LtYxYp8sSR/REqG59pvuamQV/ZkLIsvCMz
StHkB8fbRN2mv6zwhXw7RUmqjP5SlMcST0z/Ba1tmDPVl82BBv0timVgDxLmd2NHgh4SioQkedfY
79SqdMNsZxiAgcKz+CBpHA/EUVt/1Z6GP1DfJPLOnA/hx3DC8o453A7YDhWINWidFc5ECaeDh0mq
mbOCKmOmWEqhdbs2Vhi83TO+CFJJ+9e26pL+G7spY9pSUmXNQbMeHJdhRZY1QoUjSZnB+PowaoEQ
+MNCZvt3wQ7pWcQgKerwuBcxaSE2KxxcQ0eGXoOEoJYl5taDRxnXK49OmF9bcof3jT6Ed+Jzna/L
PXu8T33MSZjegnkZfahsf2Nl7dTUL3qwxtLo75UxOJDlXbeCGATsvtRCJzR5dNrJ7fnh050z1Z40
c16/dIjg+Vt4KwQ5HawG2iMLQ3rrmAuQvbqWE+lE7IjO9wrv48qC6FXZpBGXzInWVK+fSkmYK0Lt
WZz2n+brsSl5qqrTvwVX3XkZ3ZBU8g/U+6op6XltrkqaKJ2api04UmeO9/kpZbYlEm7qQF7lNpRq
8V8EdnnFD2sm6I+gEQeI2FG+jjZ/Yp/OpF8JEKy7MOly38H6SHpEsGAJvchkFlnONW1ZDyDVeMPD
g0Od6oid5nB1kreoSaM8NWURoavOizupYW/Y9ExtVxFilXJBUfVcDUC4QWD/d4IcrWpOxhbZ0R/5
TkjXvRE914mf1LLx4H3esmcE6/6kJRWxteu8FtIL3PkFSZMcc2yv+QdgVYGI6Xs1K7ctbrN56Kkb
6dpoPibpg7AuMU5AxLQQChpyQWGXaFJgXGUv1C728d4wMo0iu1rAtTJGDXZWAtN9LqH5rGx22Hqo
4zPXtlxAoSEdsbyfX3qO+dkvt+MmJSrKTkTap/SxZwXophRJrAX3OwcqgZJdxjKHzktaF8qHfcTk
cVneu3hZWzYBLy3zxmMvvyKtTmRDWYSzGzbOeYZNC393mFNat68roOZSjld0g2S4EqwfJmJOYRei
+VXIDAG+hp0uy+ysEG7fYaYEla2SZzibGZM2Kg1CVK+e2jiVL5Cri7aTGKBx84iiNnqkzLD5f+kp
MoAwViOYs6OcLD89+dOWYHw0DztB/tVjdLDTczKoFscalavO44yHhS0Vtu/qwtOO3p71c6GmB1Xn
/zGIzI2mMHWkdyqNBqqxOO9Og6bfu4bYiA5HEQV7aFMY699pjL8aQTYQvOy+OfD4SLofs6GSl3Jg
RaP4eRCrbT+l945QPsRNX1A7o69aHaqZaALj8lBWC1S0L/X59Pm7bQMdSLAGaAhDdus8tznGE/sM
AA03IC369VkFpyy2/Bp1GPvXCeakVNsdu92RlC5oRhGszcnsnPyJAxZpuVjgvkh5F3e/06655+oK
EJLKZRARfrIm3I2rCKegovCD7SV4h4w+oQ5gprihjMKF7fO3CrWA52n5zt5ZBoLwgJLGwuxok9nN
F/nSYua0A73PqYGyfXhvA7x7VRe2YieugPDCaSdGfyrUGt+Pyz9DVSrLzWTUgPaG0VEY0qSokGZn
is4uuGXnp4WT6k2D+TnmbZQ43SHRqlBoyA31F9WhUhItNy9HkIeEMIvFEn6j6k9Ln9svOOSciwqs
1aWzZM5BMYJeUqwVmGCWn/XJmtId1cmNfIymKBz3nTlLB83pRnqkWco/ogyW+0zEaAnVtNfT6kvn
v1sdrwUPTQmLmt8jzR+TdbtSG8W8uJHNak67eRIGApefClV67WySv2ekjNMGS7nCIqLMHRoueEN7
IxEFpIuBCkimzxtKFte863efsgCXS18yV8kjF5ygLrnA+m134auMaspNF80183U7kZw8kPpRMXaV
L2NJQCJt31ShmxwCZRLimq8R4pGRBIb2kSM2uM3J0uvxbP1jUX9pDOcXZVKPidmjJvitiTArCy/F
xkBdkwoPZEUHL0E3vD7pFEf9liLIZx8nrvg/zAp5G8FrkBEr5jtpYJwyMIk6YOEgQ5jf1TJLL8VU
BRIpviC+qu6v6qai5ltTfm0VEIlEc/V5XiugLZVfky6y6GHKqCQPUNRWAydT1oS80YFnreaywcxb
zSuU6ZvsvVBzcZOBi18lROk+JFW27jFKFoyILJB8KOkKyDLfGSEsur7JBtGiRD0oHvx56BN1lNTD
ddp8K3Y0vzzxPfMLtO5M9DX1tF8U4gHGW4rdHkJb+sjaXeSvdJx6o+oSpHs0F4NRqWe+VEOpipzG
LrRoDBZYd0TRByoBeVjrrIbKt2tPiDn5kufFVGPW6TNLT1hwlXGErPslGxeTDm+kWEvm0TqPBckR
BqDqKb7BhZDGRiuYOp4vi6igo5KzB2rmQ1UE9Of7acWBNFxxaDrGQaPlx+icQJtYfJFGsq3FAZjg
n+uMsBfleXOVpDooygqsXfAx0RdpiP9tdbY0P4xzPLK5uYlihpTFZIjDgsfYD7T8UVzzhYj5tHZW
TXKHhUjk2Gq8qo1yuVhSan703b4pQPnQpBD7S9wdMxwQoCEeJtiYSjMFxfAI4iIIXQnnVhODEsLo
hEKOv+PBOIBEn0HB8iW1e9qiG4c4gCXQ5TH2lfpiDthq418Kpldret901HkTFUM5euvGgzxfxM9b
CtW2CEHBrmAyEfL7bOXkuCBiLTn3h0pncctfGdCyuKwl7hlZe2/H7swmTOR+FlLAETElfWiL8qKs
tG45zC/UKPOKXyJT0yfCwNHLeNfA1J2pevcba83zyXRHY3bcajw78bwNHgZDUI8dgP92Tfmdx7bk
efPb4rB9xaVoTlZL9poAXPFNz9DGJ/w/U0laiBmRFkJIUAuyooh6BB6Ar0GoeKn0HgNW41e2uZxC
QeiStfZry7sgOFAQzjRr9kLDsFRziku6bx4jdSuitfZGKHGcZO4sYNsgL4qGzcmcfc3Fj1SuoxXW
Mi5B58TvI7ehgGkeIeNZg/+tLJ/znRLAcJ+k2yrV+AdsPhqHLjdJpWW51auxup3mBNAXEQejXHNI
mhbNVu1+71j/7s/ij+HZHKkon5+5wNBjbS/YddMwafq35/R9m6Bq4RNkoApeDiPJBYM3QjfS0eYq
EZ4+717jY0ApzBQ3eQetdebpoSMKaDrmUrPe/d1z6uSDVxbIbNhrKxzcAbgvvTYFwerdg5GGFqkj
xAoTb9OyQNlt0DvdQkEUOpujUAAh8acwaPozfIvW03/8s9YWtRXIK5PJap+kINUsTadClrr31SHA
0zzCCK6lYwKFo0Lb8G1CJqqznvdusYXocLZaGQ85GyMrMv56usgANR6PUACspAGoz6l4Jvca6lWz
CkhEe/nU8rgx1GzXAyFUfJnvP0ELh5hJq04JVptbP0Msg4k0+nXj1YCJr1VrZly3vKRxIp8tMEAo
Pwmo3HdCTH6TVT1fs9pMGIBz2LgSByqICOMcFmad14/yTJYo49qKUJXWpvgE/hx00ho5Rw8yZVNS
RJrViwm5EXjPObMeWNGnRPV8HdbK0XV4i02mvQCzuJJCRvZGs5C3032k0kai8a1yctCo+ZLx5lDN
qfd0XkllQ7ouyY4yuaXP1ew2WhXOKrEJuw+vhTi4Ij4d8b8Njdx3m6AapSnBYFXseK6UOVRD4+xl
3hmNDsYZH5wymBCOX0y7ynULmvaGO5/Ij0wrFZ9UyzBNjFc+iyDa5Sz0V01UHRwgjuCIcCjjekMR
HheHHxTqH01qt+UFHnKaBW/r9pc8oRRfvv2cHMvCDbqGjkrNe00jdieIzwm7qW9iovo4tv5jn9wk
vXImT4SrAoXV2kl/pqMKLuQErYOYeAOKYe95AyLPWTq30Sso22yO1MPW1pUONfz5Nj4iSmzIZjGp
0QYTxXzxBL8DH6wGy2Q5rklj+H+7S4JLcrjofIL8k4CkZb7uTS0XjwgIKOaOW9hO7GxiSto57DvY
2hL+HdQq3890sez1RcyO7/QXDD5c8fYaqhE/eUZMNWkg+mKuKxs/sfh+ZxqDV6ld7ppJ7oNP8e93
PSMUA2L4QAzkG2Lhp370WU5rZ+cyNRu6cOe5UKFz9xTbML8CVdpOmJ4KZMcfnTgpbDPwA/UEGuds
IbiQpy6qK6AZWiZTEmYhOaVf6uWzT8GfQWWmX3lCc2KVuDRS0hsPnSl3s1hetYIBDiULtWjktbze
tBho425enIK2hIlrWTtaNCb7v6EFCr7OHENgz8spzuw0IU3DwGvFMdREjTpzf5vuDEgsktJM5DgP
pLuGjEd6q1yL2QO0ktWgaF514e38VDhPwWyrJ8Lcvp3UyDDKQrYeh3TpdQLGb/d0jdV+tKnD1Vxl
pQvjm+HOh9qj9oWriiUXuMT/OsWVkWKfVPmm1DogLjBqRXGhlgYo/DuEqAIGmezrHqcASOd5IDev
dbhfPBt//v4zkA8DIPRT23TY3gdGir9eOQvwHUTEUVZR7sTeDeWEdgGifFQnLAgCD+B1p50Ekbim
yMSyjTCTAL0TGwi32XmIu3UwuykpdjCD0beiFuG3z2dTX8SU1lhWMG6mxwFWPLPdRbCSWANHPAKR
EvTgXBG40B7INAWZwUrZhcvpb1fhqk7KqjDVSXF75Wfp4Zd2PBCPBG2cGGko1TQQ1eHyIpnTUBlG
yT/kXR5WQNmtYDTbiMThV6jyq+65s5w6K6OWxHceDsvELdK/FGgruxdNHF8+E6gVCqlSorPge9qh
zr4/o2b5dpXfTaJLiXFC/4ZbwzqOZIc/daArszjylpUDxxoVnxKciB02FWZ6q/CZTlYpIKa7IW6J
Y5bKrOhvQ2GanW5rpScxEMhmlF3snA+8NMWOpeRv3/IrJF0iHglkmyL0QI832ddHReVf7sDxuxoh
9cgBQha+ErbPP/8RFpbCXGDfhyRZ5PAfnslzOELpHJrHDaiptHpU6YwZWNaxclFWsgRSOeeYrbfk
LeCJzxBcnznRClX4057AUQF073NOR9jH4xwnHb3ctFygmggNCP5akVI6J55LwOKxvQnVChHdlNsd
HfRbzyW+kpoVme6LkwvBZ9cz8fKvkV8r3mm2Mx4rO2NNea9tES4dy/frw80USGzTXqe4DsTcKTK5
4Dby8I4ILbWdTZai29zn6YdUAxSLiFBD62whr1SxQ3qiZxX00mKaxY4vwj2gih0M16blyfr3sRcg
uJ5AplVJrvU9zHTiQ+oo71uwKAJqWFpQA9t2CDgFGqsAGjWz8tjAVcvKY/C+23dXGmMV51t3QKkj
9rHLQumvLgKMHsv5jqMKr5kNVR5lJawAaj4kABVpKQ336T9WJ0kyO5fXq6nBw+os2bYI6GV6qC4J
21fA//bFlym8cJ2WXA+z1XDfOWaQYl4TVbl4mravc2hG80HzhXyh1JFgijcwOXOoU1FkMH/Ce675
hA08z0CQ8MFISNgsUkNIVB83gKzb3qZM9dUFUOiWp9GgbHI9C6dhE422hWmm8BPUkNVl2UULKX7v
FHvVL3oZ6fbBg9taav3TK3SzTTjOVskfFw3rdr+v4g/TSmvNWmXWJR7Am+l2PxI2NCI5kcn8LBr1
MoQ1gtie/VoRIbBYrrDo4Z8NdwKAV6csd37Avd6NuWT5hVicqmn3YQnr47NSANIGXkuHkkGV+a2f
vvdPKvIXCfSZGTHTvK4fRIYS715W0f4hTmg05MT4bphRppYuirniAPSG87pM0ngfflM0tgIo09m9
YjdjzMIyNKxM69jSn2bewyekRm6mK+yGTWQYCdWbHbSjCGr3FKqhAy6HdM8B+flZtukj0RJJ/t6+
hDCgYeO+h7+GjRtvithF6GTNaPuUHdiGenOeAHbbLUp+Oq4QlYyQ3wGS6XcQMf/dChrKhvGAfzxB
KhYvp8/fzyeOc1jVnuaBDU7QRRGL8Cf+UPxIBucanY0engPAfYwplZZofj7UWgqbSlvvrBPa2P3Q
cE9IJn+sex6l/0uFTV/dYBADStWCkRFYAoc8vml+lsqwmTtpp37rNzHR2QV0UqBddweWK3ztEuZh
3ktxoD41ZocdS5F97q382W2SmQvmlKsD/yUD5i/9EkirQODNcFeL3j/k8rxXlHAU+15/SFo7zJpq
ZeOiUL9+mY+brSM8F04LY0jNnTI7ZGA+K/ESfJ0svYTzutIo+Cu04xErU+p7T/2bOmPBTHv3xUMZ
PFQNybnW72OfDoJkmq01iw7TqQXHT7j/1Ov4dteiHA+mHlbUHyeIS2rKCvAQBRk1UjXmJjGyTM+W
X8YhAb4lqsaSpErn3sahM++vQC8+c5a1JpbNIRsd/u6jV1U18/1idyRizJ5sn9hZzm+Gu6bfBlEO
kOpNj5jipOUNvn50ytnXuG3+4DznzUvcb8xuK+hYyM+XKOc9NYBkoog6vcCq4tqFvRe0MMUjSb9Z
cQKA7w3iAR83BWO9k2XiwgnobUycms59J7e4xxTeRk+Vbv4FT1ICrFAVjyHjwpCEVgTk9qE7GSaR
IqxEBYEXCoDUYHtkMM7dWdu0lhyD5u8hMdkcPar8LDQbp+PIbpjXJ7EKtTNwgG4bYmPxbYVza9gK
2EstNZWXt+zTUxhod9+j13bPuhV0+ziESBqcYRtG+TZJxKLBTKB+xqaTmlTcBeursjQqTmD68pYn
PoKvmLYI8zGQMTSDH0XGa/Py+c+dyWo8j4GGE6sgeHMbE1qS5Aqq8bZzXO5NnexGybnDLNmZTiqG
Q6G9kOQxyFFBpoNOFl+ixloB6Wbzi6JkCAs3RZD37hJbMXNAUcKxftFafgJBv2o/5oYlcHIWf2O0
Amq5tnmADm0vvsv1u6GE/p/jD4vIXfNrQm8h1q7lmfFqmWDz41TV0HT7Gbsu6AGFMMnKnUrK4f45
cHZNjTI5+e0CgVgJdrZBZlxiU61eyncWeo3dwjsH2pOeVyUk/1V8yCpN2WMd1+jKrpdXGXtTAP2o
o9c4GYY6KEuENMGzmYh+eRTJnP/WDcx8AHA3NXZfZCsznnzqqT0379xSho5Ierm8Coy/EVIcYRXC
M1vp+Odu9BqTbdKaxb5RnadPWYghtec0EWzkD7tHTrzVGL4q57N3OjDhp5RC47FdcXwLLU2UjeGu
SGNv7rqUiyARWLzZRRc/+KohFsiacE2S8dImlnwAk8dkz5rXk3Xt934PTXecc/p2WbdalpWZ2ACJ
AtbsTYQYwi+wEBofpXgYOCzjgIt0ZgGseCc5qaxdOAtQ7g3EsU/WOuGe8mpVRFjTP9/9+FMEnkOY
xIBBLNFcRvOFz3tZGMOPhRs2sPx40LlU00Qt/NdghTrOw7RvzeMlAjjoCYsQ8vRafwO6I4sCAXMb
XjZ2Sg/Uf4TzxhiXkp3NRvtAtNSvz9BxdeqcWjYZk5rKlUYEkH3TMkQiX7DLZyKismIjNSUQInkc
lWp9TqJZN2XrOkyp7W0lMATm3mqvq2lLEXHfzEyO5IJrOWbDg0sinUD75wdzyEOjcTyx2pb6KmKi
mN7xpbAJlTLdqMmmnSjjDXQJTxYb3Sv38TSmDbiev/gIo2WeqVCxVNTwaavml14g82DwAPr9vecv
EHsdQ1Wl9bPUPpZCYiai4AUdoG80Z5Mhy4yTpL4AAhaLn/vkrHl7znCmi0sLXlm7lG6Ck/63Pln/
a2xvLjaD7AaIi0Q9jFSdVjS7MVBddaqpuxlmrucgnCBTPZsSDoDLMinsCpuNc7dkAFjsry0u0w+m
xyvBMW4KMwPgh4aNX8o/QePX3mziij40KVhrcXDtv63y8CIrtFdeb8nyeBNewaf5xZylN7yfcDGO
P09lMId7QvlTlNayzn+VK8hh0qMRFKtogbcIMk4PxgXcgwscI8/IO//Qr7F4AKYAmGSJza2ivMAX
TcaoQbIzHr63p+420ZygyJgSWLUu2ivrjEoxwM422++dm2lvmKI4ilh8rJPV72xEtnqNBf0r5seN
2sKfsvwuMONC55XsN3oDdogRziUdyW3a7jk5O1y+t711ZZDZ4TKgo2/PYJ1U3IMv5JOxuv3zZ8WL
8Ij1FCO9/vpV8xZaqb6klm+7KpaZnLpwiW7FgGPouFr3nWr8EKHikLdrpBgKuLaxV0YO2nwzaoAM
Lhdu6xnwhAVgnc3dBMiXidrqmMnn1j9icPwnJx3XEGNX+2ljFCLDpUs5wwTq03Q2yXqJj8HRfiFT
l7KrTmxRg8ieqtcbQl2+kyQP6r1X4y6SJG0+ikDF9qrBvrTWfNC8tPTyAQTbedEvnxyNGq5MukG3
+D+yBen91m4pQRGm0E7ub1FniguPKwb+jQfYzK5YxCgsDScVlktSX1c/cgjEF0KA0JsW31HxSo5n
DkwIhdA1P+fONPWekKKrq5iGUEanBTswCBycUOj1IWkFdl2cLnFEVwnz7Z8BWsVTN6XHlSiyqHNm
WeDtfc9FHmSBM6ObqK7USJgGqF5kwpl8eWNkrrvfLtCWR7hL9eOzBWpygh3Epy2JE2xfLxjzb2+5
3aEIPE7xxlQZ9mKkygmUTFWuBSjsHnU6mIh56ipSp1C0uHXJhb5z2pPgx/Dm4eA07/4hUaoMLy5V
qBgSAGDuOn4CyTJHhkL8vhwe9yrpjTBlyYNFD6uFAYG5sm42AW68mnzz4m81Vnt3GhLDaqCSRppY
0Xe/Avu2nPGuGfkWeGgKZwqLSPacUflmDHVHaDC8d1rZ3FhBYmCJlQc2pdJCjvjcTJ5pAUhGNyfi
Gna/HJM6e7ZdVb3Cfpj8+sD4MEtTqo4Fstbynu/5P4uiQ/LnJa7Qb7ao7ZXmltuwXxc7MYIFuk5r
ZFXalLyQ9/bpmEu0jhLVYb4NDItLW7R3mErDxhUZy5rSZwf4/aSCLQ4Fnb59gzDnjSuFdFSSEY0N
UCYKetIwwCkkj3H5mfN35lDWmuZ10XFV/n4zaNiHLjaInLkfaNkXd+UV/+Kzb1BF22v5HGSD3zlb
wjdaII3wMgn23VQIRR683Mnau1V4ph+F8fy/gs3jVLIWDznMU1wLqXd0aNq7/9cIdxQbuO8Sh2zZ
dBgi1K0cY69A0Q8ZN8oWxkqD8wp7ANkfIIySaXY4KA9urpuhbD5icpbJe4Z6L4KbvSJwm7SvYmAF
adJqjqcHXSSlk0W+x+x16qx6WnX5EiQ3/KNgs0/JNK1RW93UpNWfudi7aMy4uxGS+3HnXTwUjUqG
sLnzYdzhpVlKNRpBltQV/5OJYT2P7jGz+Su2tKhAnyxsB7oWLZwIfmGCPBKQcJUE6s5eHA0IHZ9m
j5mfWaOeHS4ybjGS26YuVBV1gl5xHqIG8g8WZ4juOM9mYFrVSSNosIAZ1Zbkq4iAgh+uOdYUAucA
UUE7TVSWfEhpLKT9lffbI7EV2I16lSvwFq/RZD43FnvR6c4HgSv+oFQmJoJZkfaAYm650SzS87Fj
ot/6fKp/xhxafcahefySi57kwZj3D6uy44nwn91R0LqqZQioLLi52HZxkyY/NbSEu7rA271k57dB
GVCoKPAEwGunn4rEiCzv9TAyNeZHzGNBciTqQRyyJzCf6f79ig38ZDmq/4gtp5yO7/IKoTICAoCl
c6YRYrMAI71z3axrefZJ6lPdgT2NHZiKwVIJ4jGx214xUz4wpFASw+B4nZ865TTHCg/fJjYfWRgy
fw+UVLv+xvfbQBG61RUUgk5Pj3kgeqT5CKOx3M+oFZf9AZdOk+6co5uwZ6P4e272dfrRxA6pW7B3
A6O96qb57xOVxSiz+g/CLS322s2XUvt9FC7QVjqjQxL6O09PgS4IZ2odSsQDf+hgjkgRERs60nVY
JLi+eWPgeVS0kj86aNCNtNlzXYX0qPjomJ0Rs0MuzExoHmuAHyUF2+qfuc3ZFewBIdChsHzih7Xc
tsU1z+7VN5wbRTj7WEiUuMXwakMHpe+DuefNhztOVPnXF/eeHIBSvxcwGwu+DXYFJwk+T+XMZXjj
p2uY/Sd+wMEPkIRrMaVZdNvDUwzPHl3KNzpo0tPf7aAmC88/+Mmoq6mNAecS59leYIKBS4VN3c+0
T32YDqOcX8jGanafQLQClfiR6Elq/01s68VEUbuhfIxCFVtDXbHte4fqwBSPOWVnwvyLUhUCLBDe
xxq8J0eBzo4Augp972nIftj/hnLaWkBtynyflG/QtsdbSFYdRcrlRcUnLouVXKbCJ5gWaREeaxZr
pi/p80UrrzFt023mu1O+SGwG1ZnX2h8HBfZ8CRipap95p8CtQ3uyKtaaERM0TRBCvVHHvvoiVEM/
DthgddXPRRIe9VSwu6juBMgSjWj1vj0ylHgveBDG1p28GeCxck9aMw+KseedmWtd7EnzL783ij47
mNRX+vG4l4wuYdZbQMWxy4zqW/+wqosLPlC9dfgyNbQeKdi+0P5TP6bpjuAUmoizQC/czsYIHBRV
gCL2lld0yn1r18of1hVO1JfMdGODVm8rYXA9CT465GsiRooL1iU3YmBVt5juSjEpVrNivBDJzNbR
+bXAJks00UYK/PLLJF+Hc4nSSnTp9zKJJrl1PF0Zg24dSgnUgs7Q1dG6tDP/yUF5CyOi2NraqNdV
rc2xMFev11j03cxRBnbpHujQGxEWsFWWELcFepc5JDj3WJY8W89Efb2hgB0n16VjL7DTEOROXICO
fOpO7iNrC55sdhQxMiOMnCcA6bkKJPBzNIzFSTF6EbwZQISlZJOtF2xEsImc43dge2TK4zNo8pwM
hfFQoSmF1CN8FKW4lmE1mPzA2TrYTJrJn4ZcwkeLAnozjjg47sSGS81VDYOVfgEcuYuiAxgvin/3
2YJS9Ksg2L0WCKyZdBrFwf3VhPYQO85rrjq53TRFfWGskt7xKNEYxt+ibS3OSowYCqedTVDSY1+x
yHuJHiNjdGpoUJSttX7HqoVzRCRZjmiBvylz2KQb2C5y4nfwaeWMXzKzlbINd9yumTt9up1IGa34
4XgAi0bw7e2WP1f6L/w674JvgBywo4EYARr30wVRVfdTQ0npjeGGfLCaAvf0Q3l6Zw7CkZA59i8P
qsPgqrKUet4eGUxWlk/4pbFBvYVvEvl2X4kV4qnTmA+cM8uj2hbJT+Fjzbdd0UClRB4pMAun4Jz8
/RmxXT6f7qgwaWkGsv631RGaS0lqxdGzyMoYvk+oAabswWc5cQTfuRhPpqYQtZ38t/SA7F+bMJpS
rmJaoxq0GO4H7+2HwbN5icOkdrZru0xkslPSwePpoqpMagtAbV6/pJo/ZCaK3LJlEof/kBHhz8Kp
dKZUzX3R+uEt9Us2ilc66NaEDd9Ezyb/VAhFsnLPDG6FlozWcnbl7HWFpeOs1RljZpW19g1Ww2Fa
0ypewTXvxuEImVcqPC0lQzZv6/fhdtsbR8RhsiBKYTTA6kZSWZRqu+y+qhMkhnk2J9rH1YAPSjKn
+jBS8PokaYyZ5ZOxBLrOokOPXhHsPACOVKcib3ZlGV+Rb36nGFc+HLiNF04OJ6qvjuUtv0MtQwDT
DllUuC0y4swLUgz52+xPhN6X2E/H+oiA6sRab33RQJ28qVvDLPy3KbtRpVwoNkZQMolr4XQi/AUs
csGcI1I3797azgHwa5eMOgt/VsUAoSL1gzYoS4BrRM2mYl4/YnvfycM725fe2NQlaGJiKfz4dHe2
VK5hPOY0eCIix04UXOXQ9quB0pPvBY3iKQFzbzBnovE1HB1SpREBHvbrlXVS+OMnKurOkPPmWDv1
9vzxgl4VUMgr5ycB0OALTV3/ZXTnG1Nml1tMHs849/RJM1eZzwlJJXSNWJBmR3Lc2rLhuPmQPqXA
PprN65L+8KpJBXT8SEc3ramNZmxhd7VcYInyk3qORXKV2qkER3I04zXCgZZJ7y7ilsChW/AART3i
Fxm9AdcV1COhfuJpVFgGrqx2wkwDClbUw8sSUY55zidlfumvR9LneI1hpU8zKSWCu60GSAZOBF5x
FVwNU8x0rgsp3bqrfnA5aHgSYV5n01BY/jKszVMzX2D4EY/dXjOYBwuZ6pa16iXElhzu3DU9tKdU
/soRvQc/YbNTkGLK8iEFCFKff/cq9WFM3ArCq205HDcHbhcd8wUTzxgSon+1uWQa2WDfjsa8lbLS
T5yt10xZPZr6HhIKLn/IOwjeDCLADNC36t5QxLel8eyLwrUyJ2RdMETC+IiVInf/bTUEr+dPRJXH
oTHbyATpOIUpYxtGU79c5mhmbD1KR4bn/CHhq7VJA5M8pIjxR3GleOX9hXBqLqeiGgXUE5j65bah
D41dyOOZnTjQOtuO/nC60Fu1MYMSKU2fgEu4Tovt+wVctxXJ2dBtb5XahkiR2pEPoie0EaOLeeVB
wSVw2BkCuY/TTUEg38lMvTqdh0bLZd7s4eBxuIQqdqUEf1sFXKVRErQodueeg0uJzYNQ3/SEfoQx
JrN6J67ngE+YXFPCHSuEEuCny5Cxt8Q2Q7o+1LoDuWgBpjoE7kEIBn5y56iU4l+t/1xIDlLMcYuA
B3z0gXGc0W5OLHgBB0GQAI+T8CxuYPQHUUKvqLfes6jcOQEDsOyaEhpTLJyfQhDMcYEeCjn4/KiV
Z7y8ZVmjxdJ/a3Ky++c8TH6ZinV9NzJb7gdk45cWeos65XEDThK1ReTKL7H+CPJaWN6mXMMVgf+K
fIhVsCXWxEaKPOn7R9w0xHTKm6UF6ALgVqGAJz8umlMuyU962Lw1SvOVXo2DEKce+SOncEiZtuZH
dL4rMNtSkNUB6no/j1WGHp3NOtbXBHVmAcjJ6PVz8QVDZINJsUzy8jyvtf3nKRaWmwKVsj2wxwob
hPOJarMEcrNSmuiWmh+OiOAyTSkArWFTGJQ3qfFj8yqL/P1C6iNKyTPiQQBlstEIUwRYDeZdz9tw
26bYIvlMWid+8j64ZLpI5+9R2acNJ4N4K/qEA92fsyeJDve2BtkxfcEalM0q9KzYmWHPrR+pIv1E
9aXCaYtDaK6Tg3wOrgJNOx1TpW+2KaVQ23vvdpLB+nMP9IwJJEDqK8ZbS9MCehtVUhI18+IZLcxj
f9xZlf8ZwJMpVCUGVh9d1neGAnWCY8dxM9Jjwt2k0dJ3gFAurGva/yfdHOHbzM3m5rbjOATBvddM
Wh/RIPYRx/FpkVBPKMRUh7QxXOyenKBZTjU96rHg9DmH87R8eoNqU/Klpo/K2XOKXXEb5TT1zZOr
QvPRAfqIRvngBBuTQTJKzz8ifnmJBwRsK7PrVZc2RAqoUu7Wu8R31ebsCQ0OqU9eJ9THDPkXMFmc
kuZscozVWnBrBu6fNkZD/qrlBsWACVdaTMqFBOzScmzD675eBzvfEQNh8m/Ihie5UCMKVnSPzAIR
jdu/rSQrZ1N55hjmq4VUUY5h/5rR+fk5ida9gWMoxF7YNvB4IgRaPYY0J21E17KWcgHIswgj2OXz
30mekNPY59E2c2rKMckDzEhPaz1IG+J68yO0pzGpA5/nkY9w+FIoW0Gd+73GLg/l4zCVf8pVSxQk
qxD0Am9awgU3A5VExZCwFRln4uwDXaYMwM0pJvku80K7PzX5yyKWoCU3cwtmjGLyMrFhxZu6BCHy
v3YZt0S9XGRMnKzfnlQLFeE/lJEV6zvcPgtA06EH2vUpCpqMQvlM20yGZxFBXQt+b/wQydCM51iF
HBHvblGVdAiQxCkhNrdfQNZP0LrkIMLsk636IMH/eU+OgAD5+9Bgdl3FDAtijbYs0t5t7uvulTV/
P2n/20qv8odb6ndmnBxiI8OKms1rc+WvplbERGzEF9R0NT2RYmrxncVeSY8V6QV0Sgcv5LQycU9y
kZt+XOJOac8oYLKfphf/M+8fu7KFJpY80HCelP0XzFk8gR5GyAMBetfVNQsgp5NVoTTC3ELL5AQY
6U6WUmnUyqqJvR4I2U2F5aQl+aNkVC34FgbnuBSQnhtbYAq/XrR5vbxawx5aRCdRlTG/16NcIw39
cLKeJ/bFhU1xe01Hymtez2gRkUSv2RX82bOVta4St7IY38m7+lRTKm+H7e4PHfv3Ej1PKYkT2NLA
hOe1sOg/gHCrypHJWe9KNA1hDiUh9gCKv0jrJQ6ARulZBpqj/Rxp7rLpw/Fxq3aTjYyXcq59oaj8
OOI4XfhEol0dx+NFnObSY6fQjPmJuQNDQq/d+LPLH5jM8SH0t8VuYWlzuaAToz68t4VCN6eofz0q
mmE6OSekF9YNSParGr/TsoFFNGsh3VuktQxBHJYA+bSmREn/ZRoWxTRhZvYDphNXAvSuqbdoFTKI
rqAN7vHnMp7a1ScNc47FcSLwTKDhTLPoc48NDj/uGSb1XaC9fgUWfaWu89FO+JXtOmBwERb9DCyu
3vFK1wS2PWhruGPC5soOIWIGQ0V7t9t+TZkIr6eXrH3mZWjOuskFvNFA2GWv2BKbP3ez3L4YXNE/
t1d+8JesWaNxV4sWE5Cb78+f/3nIq/7kXAh02nE9aQ08T6r7eYH9V9qB6l1e8vMVsUf9GaXxY3Mh
f8Sl7jibG0vh0yH0AfjEPPeSrCpIHW6b6GG5L4uKUqpAo8nnpjTNNUdG74i6T+aYeWKVN06gZ9x3
P3P9he+RjgUcBLf8+6XgJ+34US/A3xS+pcnpfCFgfhws/jqdA9Lm6p0kwZSXgCLvjAHuwZWZ4yVO
oOgGIBX10MH+u3r4sNrqRrvzxjxzOsGlVyVe08RCqwhRyhpgzM+w2o2wrawdKVSTTNooYMOQ0jnb
ktn+T+Lb3iqp0npSi7nAmybMuNAFZ9lxON2NREtT46sLoyAHjEkzllfkAsfynDSANUWkuJyfMvtU
1OWN99Ds6CAlTesZOe3uXUh3M2tVLW/lDIKOSlwk6pLO55uZEb626vp5Nisw7A0N1K7CtoX7Tibe
oip6egaiAybLbgPD8zMNbeL9Z0ob6ZVdXQYC0KVuuRQd8hyHjy12Y3JSgE/QChf31ESM0dBg5zVL
935O17GhM4jqNDdVFjhXD5ppJxS6RdxYHbW0tckGNNYJ3hgsmMOk9p8m62nEBTAh2A8k1kO/WtaK
VgSiPm/mjFX0AJ4YxpPEwhyVFl1MbqLhebg7M3ZxcLbZXun5NtNXzdN4/YUclOTGMNXXWSFfh9Pm
+gKuwl/uG3WDbyqMzCS+Mr2S4XWz+s0TH3z/mV4Nc3O45Khg6Fgm51sAU7srHOD1B4motgFzv6DG
vVHovhqXDbXHfKnWNzTaiRTJ5M1tRZSVrKe77uQjl7W8kf1NaqzeOv/P+cEkjtBVvnKGHwAPtE1B
SZEqUH80CSHUIEntyl/1jeKiSRXLK18QABEXl0nTIbHEGLqcyYLLSxT6fnaqMUqq4uHYl37KUeqV
wHEzRcuGpOklTJdHpcTENW/fW+5mPqe/jn94W/FzB5hGOXmHFpW02r92/KnNbrqHOQOh4EpHlye5
iP22suLQdOzN2No/aEH5O6+WYV6FeTIHcmgtqDSDkIDZ7PAEw+a60P7FhmL7ozn/xPv9ByvDUCXU
SicLW4kg9j+gooyTi72xTjCmUk0HEESJz/XzoCMNL3PbixLHFHsfrCqOtmthhTQ6EGASqQ54Aeu4
CF1uR3fUGLRD8h/4nmC40L5xryFClY6GdjeGNV8oaHLoTPNuelssA4lj0VS8k6dUV8vIR2igJ8+C
27lJvfCQtAw0uhpMGKDNll3Gg7mx+8S7l/7J2FMkaFEg28qy6AP2Rtg4u1e21e1+sdzqACjKWnK6
QcDlC75l7eMoOLn7GSMtRahvxFNvTzFlMB/II82ZjQkDbzrFnbUk2LtOL0PI9prQSEV9QOZQHdel
WNs1N7OQ53nHnAU3LQBDJz6RDeILyA/kehRL872hIxm7saSV/eWxNn3ROCo9spGeNGWDw5smu8n0
EL0/otTNs+1YcN2nwAg1jx/Wtvai/wPWEzKfZdqOlenfx4DqTmPx0jdMbugfBQ2LY+FOS9LisAzt
PFvUaVWl4lgiKPnuHg0K3ougSj0awTUJ8x4+IRNahxIEb+OtOXIueKLFCEq3m7XcWgk/UbxzsnZw
fFekDBqXgGDOFWMp06lFFmoZV4AGdVlMDxM+LD0GMasCfVgqBelxBDgDYV0s+8T0wvqooA3IIARy
eXHj2tOZp2Ev6KRZFu9YJn93BV4kKtj0Jr+dwW2aF8B4iQte0iP9DeaUeDldUq8147O5l7nRGaXo
J2DzvwMjbNIZlG5QcDvBfkrBPTf81Sk4HOQhPc3/uUh44MWw8VRLK6ek3/zY8isQDnr7CvQeOYH5
DXx3heS/Y0YNmPzY+Xt+R7L69NEi8YpZglxPk0z0uJBJDw9O+txqwJZQ3g8xqOgwv1syKaCzBbgb
P514lw2LcUpWUQjnrNc/uLqvQl4AA5jWEh1DNwBwcJhGRP+lO4F6tLuJH7dzTnoNg+2HC4rJy40x
QJym1gw5hlb4GD8eXkGvPXRxmyzdQ4trpS7Dp8Iu4KdZtQg4QxJevB5BuBGzCFtnzie0Fd2OuF1J
93BSVj1CovxQbV/FcBwF3lQUq78ggq2+cKxFeW+yYpJW/4HgC7MB/dC1Uw6jP3zMVkI/WDET7gfB
b0IMcKNDJ4V6UwciRwkrmaOF7Ud3iGiEdXQ/0Z7yctMy40uL12n97ccLsBUOMWOYobYM7tQV+Bfu
yTOiMvr+5VKLdwGYmiBDF+e4Sa6lfNn1s4E9bD0OZkx+VDrVw79QMojfO+ngV7H/GKj1XCjmlHHV
YeqR5PDpsmH36Vri3IZ2nsZ/hXdOawVhPXJaQTsl5PAoV0xGGm4aiBlA6Gi8dUorY7E6q/PLan9N
vAMalox8RompXNIPgvdoEwQE4bdtbpgFdHFv13hHR0XsA72BtPLk4ZSz2RisLbkCZjZKQHJWTTVQ
pLlZxqXbzH66lI+36quyHx5oHnDcJUow4IMg+zCqvrT1IerH1Bds3kCANwB0KpBxQp+gIZTjhkkp
8v48hhIAIBjlaKXlE6FPHIgCPsgwg/fJ7lRyHvzg4qDF4SqBqTcRSr3eoeMU1WrRG3xLSn2gAscx
B7U2bUojaG7rRNoS1k1oSLNnBLGVwap2ry2AbbKFYFULSOXXVoumO9g85UzhtGWef06iTJkj2thR
Q+7o1vnIe2Fi/I1K+eXXwRFiP82dUkBenQm8c9iPVEjU5W5yN1ZIjmbUHyW7wQfdlDU4jnDFllvK
tCtnWyrpMqAXLPjib3qw/V8uCLK1h/jb2DDj1AXMz5E7f9AXuDBQavk5rnVABONtoV/+gvfIreuZ
QkXqSlgzcDWrcZ1hKCdJGpbPeMFMOWVVFAfQI2gw4+DuwIFq9/UiFKnQprRTTyd6WbEzgxLo9udi
1Po96lNYl45cyDJ7H+ign671R8SNMLTOxttF5PVo7KptEMoKd8lEKWz2ViDyt8jzTopuWRZZaPBj
M0LvAzoxxBlJAZYP9phtzY0q/zPzHLXroaDwdAJYDHjFfn34FBHYFJIXxS2MAVe3L7AfKcEktDIV
z2BLOBrW+SyXQyyWUZ5S3BtkeA48h7CSrKrEFBWP6vuBU5s3AdtaEkhNu3DElM8c00FkySsAqbun
Xi6ry5eJLEltTxE+lk4UOsLTUY6CD2ITaSwM/uBbWVvHkVtsbPZU4x2VC+p86kbHgJVeVTBboRdc
AlzYfj+hkUl/ebMJ1h6smHOkTvFuK7MQVWNgVi0zGCMUNJ78v55PaW1hIIeRpNhKNysmiPrW1IJT
SqiKt6p96feiZwbmmjT6iPUtALX+vGUX3sk/cjjifdFztKxzrmp/t1Fvip44RtH7ApXFWiLxbOns
NlivoqiD55wv0XYz7+tdn+M71fvMAeQrD7TWpu0U7xRhp+1o6HlOfEk0MAMu1CNZVSdF8wvKquYI
gpp9NtpDdhMHdzrP2Uox863RQNS8Twd1vxb4pOCaDEgSIdeADDimIxXqhPRDwV9pwFNfyp3yd9I6
j9XjqmXGsDBi8k26/e+NwBhig2d/PH7T/Z46qXyEBCosqB+m/DnkBnT9ZyPpnlmg7M4pSEUJZSyK
iqTg/cydEDvFBbzVHMoAN6oFnRVoOk+hJqXHoyGSLuiGeLc+/cvwgPOvCrFOCpptxLd4BCZogPSV
nGORLHs03ClyO2iywaHC8ITEqx6hqn0mtPq8TsXL6oic4gEgSBdUH7F0XhWYIqU/e5KTFt9KJtF+
JM9Xs/i0a2MKAMVQTBW4TmDjNxlQQaXv1wVvKZVIDImUJXYrFy1vlKiZtSRXJHKcun4IfV49thsh
r+00aY3atvCgWJhgfHENMk8EgO4Gxdko73y7FnP2zM7Jx9pNXYWBJOSR2JywlY3Nm3cl5LqqtihT
GnZUpX1LWZaP44XP6JlISHxZKho1w7IWCHMOzdMiIzNkQPXirxjJN3eCLLdNBxf+WCoxCEHwCiXp
WFrcloQoG1Wg+YlhoojagAqE2mEUTavmyNJnNTbnP7Ek1i+Qe9N+E1vIvnASzl7NysCd94LPvRuc
jcF1a57Lzzf/Cv/vFK5LCaWBWhKMHciOyUeBWqV/EYUBCj41gsddYumsG1F/Vbw+JA9DRgwcd0Ez
NkGS6H2OOuInN3i2jrjrXiygpZiJ7x0syZDS5HrJhSv6J6J+HgoC1c78e9OW/rbzO4gRlEBXBYLE
VAqfES3Kin04wLin2rjGR4EpLA4kjo60YWvFJ6qRTHfDgSBrq2yhKt3KIgVwswGtqgVmutGgOFFZ
GjzgGQJ6bvg8EIw1shxeCiSKdQoPvqJHK22t9WhnI9zEcAVvdHiyl/Z3/UQ03wIqdvaeH1uzo02y
s130bgJQuTDyNe0kDrj8soTsOA6icv1Mkr6iXVHiiDDKqRP/vPSR/+f7j7kWpRQZRJflximipdmf
xTu+7vHj7hABANyVOgvtRSCd2jGeYGGKqNIbTIq2wcMp+LdnG+Ri+g1Pkx8CRQ00jXdWuION0kty
/Mw+wkGrxp2qi3a+ww5Mc7ZM47muVhyU5XnqXJ6BZR1a6iDajfURRu4EsDs7+rYA4qRuHTdeUN/C
0C7LL5gvA0SoqFgTYK0gpDhIj8p1A6uwW9mIh3ph6bMaut7zXEIc9vubFXDtbJr4xxnw8teSTc9i
iZBni4wDoazLe8FLroBmjrBivVoRbrE1tN2Sfv8jCUgY15rOcP1PS5rGV0MGSfxjA57ete12bAqq
NHuPHQK0TAyItqVSqFRri5hvdP/SjMGiqWy1zx9ItAq3GyksxWyQkIllGNfuxxn0hsEbfuq1IvzZ
gpsV/wYDxjnW1FcOw6bVNR0662PnrrKnik+DM9Vu3x1/6h6CBvNkKY1rMgkQh6qdKPI7B+zww+Ry
ZefS174Z4tF9H2G0FCHumdOkMzKMHffvdliRWOIVNqOZ5wC6H2MPslXfXV7RAlWmhIifzMqumwmt
zc5XDW7vrAnRJhtkZwcJ7Q2gITNsUw9k7ukor6Z3iQz2xdpwoVdF2RhPhP/1Ub3BfH8MKxfnUIqO
77VUYjWBGlboZFOSJvVHljgjn/msIxYHA8Mp1iFpwqTRhAZytgWFfb06uibzIY5K/iXuhFds4kno
B/psgE+llAkOW3aqIQByO6oi9NwV5l+D/WKsl7xdU09K3hq3sjmsc9kS1Sq3kXmi9Btc8Oohio97
WCOLje9evR3ZrjQtxNZ81SAPE/HedH1YZUR9c130Fa+jdSepKfAsrp/Liu5ZH2x21QHcxtrSAwLy
dtJHJo+5tTGT4VnUtLbMys2vNSL4dqT5mK38UHHY9Jg+Dc3me0vLdKbC7o1Jpas5r2c8ONy0rpsT
DIIJmEDf88ncamD3kjhKuRhSOORm5GfmiRUEeHd4ZzyKYPAjtTBa/UOAPsM86lw6xmXVuex4bKEg
8LZ6Shdv6/nA+2CRQl+jc716N6VuHa0wN7g/3mZGUtY2hEV7eXwhCLe0PTTrxusYwEIaQ96IvjTV
ObVSAkYKMftKQf3P9lzLiNf0rstgCqU3lEpRP6TaTNCue6eOoWO7h/JIoEoaVm/zPHL6hN7SeUC/
Mwdui9/cqE+bhJ+Dr+3JuZ/U/tzkqz79tB20FyiYYMDOH9BvDwOrlMWsnYfyaEQNIGxB40llT3qA
e3MnT4c9KHzctbO/YmBblUs0tmbwRUmKDdpHnQ+uD8st2X/0ZE4PBj+i4Z3itfgIzrmInWMsINtz
lpjTZV1uzsoG2K3DX9JcmlF70A9H9BnckPrkS/qWdjoK8JhQeYlY2sXpn+Zrd+mFDNGi4/a1m1mK
eEAJw3ET/fLuyatWnLiWvl2fU1LPkM4TQL1NmDK5yE1CFvf1MUrqfy04sTgQBR8qawUz186oiHI0
WuUlCscoGY61/C+OQBrw3TisfyaipXLOh3fXwgFbr3mYe1u+Idh5rzF2LAPhOs9h327YGuGDGixR
aFb/37+NnmykLUGis6B1OxNdQ97FREpdEQRAsbADPMIVAKvHC+sACnnSE/areiVumRot9lizE2P5
M+6RuPMbGgenDaYIEZQ29NTUPwNiJqMRKHfFzILhh+5IkHOD5Pi/4ccSXciIjgtKfgrJiUL2nXfJ
x7zgRn7VgedLIZS2HutAZqLn9F7MY2tV+zJ+Es5ufa8G3T9LT9npjV7F/RRz2n3xUiEczM3wPUPa
hGg0xJbXEki5mrOLYd6q8yjxZOYYiPpUoowuJIOHR6RrN7klYJ7n+/QQ5MeYzi49QfkqabkKkb8t
c1tgK8N78y6rPgt5JaJ7L/+Y8YZoPAUJuaOSimEZhhmeJypD4jLy/7ZrwJlo++ar6lv8+OsVnQbD
U9donyb0A3MniRYxNH+yCK4bTd63awxube13MeRE3MsrAL+17kvsDPX1Sj8aO6uVJ+THUbNFHNjr
acypi1ENYM71bDoxh4WPaHJ2lJdEDedVvfZ9n/ZYGVC2zv3IOSS+OZE6SVllaZEZGDZg8lNLH3iR
Pqfav8ADCVCBGLtNuZUBP8WHg/T90PD0fY+E3KLrsi1xIAd+C5gMJmsqOl1GUC/Gp1jHSzKT/pmt
Knr6vpOYNBe0VmvRpZUfCmhzMZhzcHOJQB2HCdWmWFkCn/dvK5BJGWFx0Ica6iJIY4CNdmvEq8tz
3NtbGTVGoa1dZ7lHuPRimz5OtSTSuNQlbDaHSDQxl2T1OFV+jC4bzsfDs0eJovU1PUWCHr5wbG7f
4URiLo814ARc4qVny40GKeLC3d/+huZ2pzxaTI7zBPlh8Dw50uJwzlA9QFicbmQhdgE8I2kmaExo
c56jFr0yQJPFdgSCASagxQGTxfnBwzyzpd6LO3iX4qZwAQ5q2UuN+32He+clKLb7IHV+ukt996O0
EtEaDKqVROTVWgXhYDu3eCHTVJiGWpSUHNNRezJebmBmPb2+bJu2jl7ihmzj+6hrzUHySRV/Stmj
jbZJMRdgz5FCy+AM4+3GQf/gyq6k0/hI48s5FrVwcx5oebH8/jBCELYtkQ56qx6eAsEZrzM+eq0K
8Tas5pkFoJ6BL05dScJsEVvosQ5slcl10atpFbaS+9ORCtSn2divQAEbK8QdzPsdLLNKu6KaNVtu
m9S0qQ4SarkF+RE6scc5r+t9Vs5N6aituxlIAHzffdkRGYPgxcjFNBCFIOPO+kUVgB/13VgCWShP
Qw7Lrp2DAt4JUOenu1Cj4AzgYDSNr4hPBtpwWmunN9m2nYVBaU+uN47eEl5zdc6gjnKwEusNNs/a
zX6273i573JnxBqMENERpNLV5o8leGpHumOy5W2s04qNTamlxBrb5bZqPn5TynAj3Xozck4WCUHu
SERdRfYxwElIuf2M4h/xNHXRpCHi93VVJE/XzPZOfH3KA10R8FNScJBuRCJN+qBTys/QhKLHXo0A
2egdu41+PEAKgnRygWCHmBxepmtD4u+xibl/QvguIXqFbYwNHyAyoZ+0qHJ/YecWarDJA85UbcRU
yIPTQ3qOg7Zl6wAV1VsY2KbWfvqP8T9FsYfHwfi6IcRo1ZI7eEL3LCuqsGEcdBAezgQy8atBY2D2
SjL4FjnLgR/kQeaUmf55xWQNicNgJO1dPnb431GYvGCBu38nVjqEV6YB4So8kaHemrkb1hazR7GC
ivaKBGNt0vo+EEj0OEOMW7j3Q90mtAaBQsbTHYeuAPNOO9zoleEUbygLH4gZ0CMMVB/wyqA3VF0V
14uU3uTVcWHLY2pdvHMZ5VFtuYZhPGEsm2XiSkNV4nW6uD3dB6w339XUbIwFq7fW0GwFzNeVbRK1
HdrOaE7aQ6mA4JeM/+x54Ucp99DtjIsmNN6hHa3kq10Mpv2gZIg1Qm654yyT7oaRRcgVvIqU2UBp
MxpPURXpthMaSMAObdJdbVojYxBGXTBEHPcaLtJTTzhic5/46j9OujwUhZa9peZ2PdW9WaKBNO0T
P1fRid54dYH7KS9rcwQo9Eyf7JpVg9Rvyyr1nRrtsnFtWfbUjDrvyvDpKV9IizqNB9pSQqiZLBbL
qf7rCNVz7LJILFJqf8X8rsBflXZAIHar9Lvgb1qi5sKVKoK/4PYLU+owFuwQ4w0AiBqsidoNVzA3
araQqtMmYH9UU53/K0MMifp155/yy0R6jhBLkLfFeXDDLQJEfVmc3NxyGdauxrN+dern3zKBsR+u
9C7Xaytqpud/xougi3OFW/GmvUt4E+QGa93LHtfxkLQaXxAF0QgHpXCEmbJdW79VmU8BusdNuUo/
k1yB0djhVZ5/c4BYIdA7+OG7Q6uNtolSbbv4Xd2BYXLJHVycwNjw9qvzDAAQiWJn/sqiZWAKJd3K
2ePYgEJ6i8gnFbod8aD1FuqPafmXmcBWAfqyH2c0Eg+zoReyAOYcI2uQQFEy3u7DvdPLrKiwf4PZ
p4rpRNfKUE3jFU39QuKqcpmot1zcFQYY4Wd3izLOZQcDN+cx6mBes8Yamos4Jd6bsZYJsdbY2JYj
ZDAt60ssXbwF6vniM/jltCitGoA+hPdqEfoLfxqA/PyvOlPcfWYM2dLTvKJS1eSaXqAPKXFRLMLI
JItvQI7Q68HdkMvY/9ATbEHXXO5FsGcd9YXZQ5o1zQXUNq6MeJriduUrHi2H+wZCPtSFmjj/WE19
ls+E2R+8ngeMNAbv9SH6A1ZHrOFKnrX/odNOO6YclCNqmJT5Vp6E18pKW8OF/Svdsekzgcdk2sW7
Q4Di8x5R7LfKk6e9WbQq49yZwNXDUjY1DjxWF8mOIJKckQybZH/x75LS+HAbxIdAwW+eQPyfLEUn
3f6iCauz4gMgL/Hqd1jQNzukvaLKocSUIEMNoDr2QuupPrNMGRummASxv0OGL0UWt1NlX+Dq3c1w
IlK3skz00xAAzL2c69ULF6LbN8tv/lPUsfkMVZ1WApUO/J8TSz/9FVHO7WweqTtHyRyMs/DWrfE9
6f0Lxl2oMqnzlO18TjRzxahp2Xsb1XO1Cf5Z5xusFYBOPYX/VhaYC2mjmFiEWZJFi5SNFTNU6+Ek
SqAdG5EYqA8+tyLEaaTBMsRPJbYUGvQT1///JvmOWdZneBWdvQ+UdLn5CdyPL3MEByu+hNFeBnvM
elLHBKVzvee8Egb2k6Hgfo36VmzYKtspDjAfb9yR9CcGuMvgItbf1r8HoEnxX2QLjNwj9Gn+7DOJ
SOWizb/9cY4g8VQssCgt0OvOS8Tl/xykIycMi/aGHiMbJyr/xXZ1IwRbpVmBX7fXMujIBkRCpfwx
yfah3ycnORTWbWJbnyRyE5IqGXz/0DvEVlya5y+gbEFObVdXPGWDQupiii9P4s++cuqaQkfKE1Ed
f5kAPKT+xIhruRHh7ZgrfbdnIq6IGIVfQpCclgs2iePjbwot0JG8u4toFY9WLGuQ5Zzg7oTjDqMS
AoL8LX0T8M5kRYYhEJQS3eGqh/KJGoPSbVy6mi+fL+B8aShf/dNBQKQ93DcG+DdjZD9dnQD+39aZ
oHM/UC5mqNFkt/U5fI5fY67M3Xoa+igV6aa7PcuxbDVHOBmYqCoSRMC+olxpRKLA0aX9HTtF2LK2
gHyOqgLRr1fVM02hE4UI3Bk7KyOHJJz02TEtCj7fpCsBaEhaAz+MHhg0pyPaSXzfVxDRW79vwCu0
2ufRZWVzB5K45pePuZE2+bvUuMM9A23OwkG8MwsZJ08ZIIKKSNpha7V1OhI259He5u6RX2tzSdp2
iY85OaWpreqz9oiIVuXD4RYrFHJf1Q0+UFj1wbaum5D97QqgT0rcD+9/M/KzHULGX4TLy35EMPMC
B2Ra3N1grcAb6EAJJ098doyE9oeUG9pmqOH3TGiwysYHX23+/1OwiNP1BXfBIFKIwOuCum/c/iZp
w7SozTLHt3dNdWwGfH6bIbmRZucwbX4uH/2i0czFClRapMss0Ye1YfyJ7EgnzQfYJ8miBB18xpbS
oxd4QJpJAreY8Se+dH51pgtJ6m8J3CD3Q4uGVbq/HY0pH0xkwn9e7PINLD/iWAaVI6O1HGYTnJoj
48ZRT114hEzZ/1UYgvb4q4gMQSnP+UkjOkkRDC1hDHrYQKzmazaeIbJvmhuY2qkROv7qwdeE1rkA
uZezRHhkfClIp3rTss4tHt5J6fWB7LVW4LctbYj4VE4zNAH7cquWbBsfrLeWujH5v/sNU4oQ+R/a
wlth3arogmZNcNgCv2lWGc3poKwyhbbTXFOs16lCo+X3yzAkO8oW2c23ZNheULu+EwAmEZxm+Ge5
lXmVdB6zHsT3de61EYivSzOMLih5PcaWUze/R1G0VJo1DGIY/02tyzKCS8XhrWbPB+NhzAI/38Kh
L6lTPFx3tZOmlQVorKVdsJyNxvu/urY0hJUCzgr66mllGqBGLXCZLMVVjWI7CDviORvFUR9KHKBd
TcIFIQVEZl+d7hztUj4vfV/19PbPy/5aKmSXlh3ftMP0LRCZf/uo7zrkTyGHciUsVd9EcN7n4fjp
lmd91MDOPKsUhOtjWc73LkE9uvj11Qex7PwLWy/nKbAFhn1htQNzYTf4kJJXGktnSirRgN+i0vSF
uxMfgVY+5gYbx1tWgVUQe1V5SqgdgbthdOaU0B+ajDJy7lQ0Xj6NhaMaGVAqDWmACs78Ur9qm6bf
U8Mk2Ndawl7tho53BH2yJkdlCx4yJH61G+0IuOL0KtkWmDA6ti9u0WVnr92WN5mgxOX2ASypKOSE
1+NtlDcx1Y+mXX6Y+xcmBMMaUSoR3K+fwKG9VuLvYpBJA7ccDqvFufUluUiDNruBDzQy6Uivw9Sw
g3QomlEc77CHFehbFpWKqxIbfpgi6T2211j+hgCfWoDPHPfseiimqMTDpKd/pGz1PxNnKnapK6zx
jCVMlnYNEQTmjhJkT+q0cerWyy59zijL/zbjMXH+HxhV/BiGx9oCrjpI73lKK5G7me+e975bRYjx
SZZR668YlDiGzsAHReLle6GjCYzlSY2FEPpTFjlBu5PSKXdI+RSoLHSWuqztHsEFGqMNaYmjzQmH
iMG30fQDHm0EqpJmbArMBOk31hR8nVOxuUsPHwgGkL2w6MIdZN0XlNH4kWWHGm0NxgVZ2VNnnjXr
FY0D6/7EhG69hvDhc4t6m0iyCg3qbFks3suGrRL2t9H233KghO/iXG4ACUm7SvLSLUAHkgory/nU
dmDuZvtfV/1ctZw8Cnl3hmAQSUrMYjstOKy3nX2TlMiB1zLTanfd5PNt1lIf57dkdeXewblBsgXv
Dz3njn+QxJv7Xxi/+sdjKMvYbr16BfXDU/Iv3cMJEMSoOw9GhfOfVNmpIE783Ik/lvP2idl1LXSP
XGX5oEyOnSAkX++Q1SYEbulyrWL58cgCkLlmFf7cbyN05gO3MWG19lk7CQnuAU5vADaDw/ZJgu74
uSCbFOk9V1OpA0eLBdcKB9jtbHw4e4eB5CNQjmw0hwsiceiZwOgpEVBcpXM3Jiu27zHmHPK/CcGV
qaq2X+QiQ8f6Rsfrme8b03WQl9nM1V3NNUpqe2GIZRQC2e0CPUyA2KivelzsnBxqK6e79rWiL5bm
rDKoqwxP0MUwE9TUwYokigTmFJkGISbv9s1NVJ8M7sKFy27rKEqInSlAbwzY1qLaZqhqE9w8L6cr
aS/IIFKdjyDsrt4+C9BzKOnlwSp9ttY7H/DCMFSlv2cepIwhFeVjwgmYIw4x848o9mBngBLTsZQ1
tIJXs2T98xtLZo4lyQtphaSwaPo+9vlNLK0l2KsjHkWKQmJRxWHmoWs4I2XqM+P37cDYrNc6wEX8
awgg/kt3QHskdwZ3isQu/vMG0BXbkEu+udkt6cib2xn2v5dURdpPxcsUy5lrP96Q7cu1UPDBTZut
ArGd6xxM1RFPwUSn2aWxXz3d/lJxug/R/Vl1Dgz7zPVFepJ2Ymp4V8s5LLYhubdOiv7oHcC2qzV9
erP2d9jTFPM5XiHMF8gti2iGtmExZLaPU1875YJH7pu20BpTlNppKDf41DM/YaCBM2RijnmLVrmU
4HrXXoM0hgwFM40d0U3qxer+/5O28Ok8CJK2ygfySQEv/wxws5L/T6vu9NtPam26MHhlHtFmv8Xi
awONpQRKYj8iHUBhk0H7xU+8HMxPmciD3KUqOhf4yFgQLbiIge2+Dqk0NG0IXyaRsYjW3jThywND
LJqk71ts6tiBpeg4Zd7rtHM3B5sdYZLAOXbMHKhoNtaarRoC0WhvnqYGRevxIrNbkXFVh7Di92qP
Zf3ecysqS3rLGIu1dz73soxrAXIhQErR42yOY+SLVAUcdPvRaHhSVgFJO817YURyGGLpH9OKXMez
Yfprxqp9ldkJQxX7waBez1b7DUzE+Z6mGHYAL4fAAMj5QtqOCjbwLCbF3/Ry8k0VHX9B/GSOreNB
D78zSRHbCAcTRD77KFKKsCg6DoqEJomnKLl9UR/BzecRiOY4TbFTpnuFcgW8s8xdBrjOIyPcHzvx
gVqAedMrNqmVTwq1Oe75LaAxVl1tOVzH5xp6IqBoYLdmyytvZ6NGpci3mPhA96G3wAze85T+2cuy
yPsZN3PQpTTJAiSNvjWzV77xdRHaoMm8YIqoRhvvxi7KT2VAHN2NjrBlUQKEFgvCPEfBG/0lsLiE
/bibF1G8yxvLePQbb0Uzl7XMFvk+lGYY8LL8+Z6YSwW0+/UK5Sgk7+jQA0ajrhU8JjgVw/Yo5yGq
GRUSzqNJOEGBK/VKE23et2bm84e5JJE1ZcZrdlO4Ln4cAsbnh5qYYestcDZNy9Dn0qu/DzYpLztE
3Wbm3RwdCGeAawPXoxSnjxw+xB/uuaaF7xfEQBtxYZK3PYtq9zP3WN0hY+WP07u0WPliFD5xJMsH
utkXQ77yzUrkrnNkCAWm/1JcowiwSB4v5PMyvqBN/2Pdhw9HqfpvPeWscODvE8T/X6k8zIkz68NR
TkeL7o7j/NX3xJPUPO/07vQJjEhEo1+Nfcq9vErrALWKEq83CshTGplPbBs7nDPYYg/83altr7K9
npXBHEoDskuxauy7MFRizBoHfxwV6eH+1FMt+WCHNP7LbXipYtE4PEqV7guYszH4nQpFHHvX8aeU
rR7XonPuXy96MfSP+PdDkIjiZsTL63pQ/NC1bvJP/qzfArPIkplsXFOSIIvhPUBFvitVDnPvOdU5
JZvLEIcFmO9uTHVyxH9fF0a16/+8T/4re2bMO1GFmdryQY2HKAZWk2RWvTC5p0XVGJFqM47nALc1
cYZQWM7KSahjy3y36bFUf5M42RJyYI+DgU0XQ0aG6qC1fSRtIONAYFUNeinSI3SpnU/iGTEYa+pQ
McBxvlwzQ/xRIY9IHvXBpOwjHPSS986MtJXqZCBAEvTwHOUCXAzeGsMOfvYoLwEccrwWv+Agv8SC
pFs43ngHJvlTQs6zlTpNGx/h4zdcpn3fko9mfsRRbtL0xtdKlUkhYEOasXdwJxP240Jn8ZNvEGVK
u9cpN0r2HqDYzS1QP879YGQWVP3K+lHGuQ/pQ39k3AYz4GcRaF6NrNd/JrkhiABTgNYNjAFAX+S1
tKe0sKxJf1nBc8cvQgslAFffIq43zP22tht2RJYCLTQqJfTF+7Vk7orq9oFA0iTvL0NwcttKyT9h
M23CBeVMGWlFAB1bHwz72qpFljW6ja6jR3dnisUUTaPWHWm2r5PDl9MwSVZFWWab0BqXAANjP4hq
UqTY2jOYrHxY2ZVpX7ZBn6Ect9sSHAUTPAQkJMwg0Mwc8EhBeM5VJUTgHbAaPuuhWJLAEN3W4TN1
GcmKHmfyKg/P2sErlw/TUNnC+tc1NP8q1iXJb6mkXAU5TbRZPXV893dpDrrHrkPOOxIM3zpz9mfQ
/R4y+7Kr8okZ0qecLc3Vd57Zwq/nVwoVxIcX1qKNxsmouosXQNdXFDe29wem+EP6malTFtDqIYtG
zsryJwXV8IHaSlAQX5BOZa25t/8pGiN6QWGmMpsAaTfHeC362SbMq684dQJZVcJ5cDQWPVYhSCAg
76pvxAQveKZTkNmOq7/bweGkm323J2btv0fpL7Utl0Ak83fXy8ibpNULGVLNcM7trvilq5hGRaeL
rJMsYgUXGNdFk41lyCZesYPeOMNPQjT/zRTLRQG+75G9dC9EFTGcWofcqZ+0Z/m/LjtIjdzWmGS6
QkZKsZnSt6XguaVOfkDCFZPwNu8IS5aOrwzR71CHgNSIxC7AVdnQ9rl5v9PIIY1BBvviQBintD+S
5NJg+rmBnbQdPLgicNY+TrvYflqppaEuNpFR76nrBjkZje+/1c7FH4rjO3LiZ41SFViV57xB7Dbs
dSfqLPdv82bLJ7PzbbSDEjPL5wZ8sPVUu20lZqkisMxFa9/MF1YvwYAMxdxtEigAhKVqbURVyBoV
O5tey4Z4VWPrvnXDyr09j9Nt9GPwF8BszQh1KPNMoV/mZ5x9d5t/mO+wLIGoxKJvyZ3IVi+Mxb0w
MO92FhcxdoSIq9itemhpY+Z7ytKcL/wu26ZafexxPGCzak5x5DqIDdcEShqMGh1uUEfYewPBhx0g
cwFVCFy++4BP4erqVT6OkM80OiMqhfu1rUfUA2vUHgRySa+9H09en7byqbZTJEIdwj0LFX+pAZgZ
iKV7jvSIQhPqM+08myhZWuJLDvReRmWrYCRz58AmZ6XLpYK0EwZSQhc1VL09dHEw0xXjzMd4t9Cd
EUECbcxWQBoogB+1wGjKA+kW2OGs9nOz6j5l/UZuhNXJ4LJMbQz08ake98Sw4MPLoVLq4eu63C2x
9qNXqVpjhBUbWnbxt5OTWCj9ogvGC3GZttV6JcxuUQiLWeJrXrqWK+j4XbbYZ3b+U9xN+SZK3HqG
MnDOl5mQoVf90StWcdfGSjMNhUAhF4Zc+milGzYX6Nwqpi0EwaEuOIYtbKRKCc207ID1g8fGXW8A
awk7T5I4HK0Cc9Vb2sTogGXpWMjzo/x4JjJPV8EuvGsaC509amzAH5KnW2WOgEu7x+LUcW9ZVKa1
dqsoTmJPi2p4c8FBy/xjI+A6bLjHhGEB3jEWWC0CvcEbzC5d1DCcwt7PCxW3fIdF07bBHnAmb4L5
3ybe8ILqTJSOG5yUun0DFFkZy0J2xP9YSZis1qUGkFXwRhzevh+HuZDlwU8xAhkspo10pjTQprJI
0T5vPzXNZaOEA8ANwQwMHOroBbo8rAuisRm5EhnbY/y6UUV7lYs8Upd2zd91B0fkAPkQ4xLSjkm5
cQdTqOLKNBAFjZqKwjnzSfzDfgsd70TkEMtjcujFmyhGIgUxJr08gSBDdu0nsI3KZWIczfF6Ham2
aW27Npup2mPGeQSL+sEmXiLxJ4bpFj0GK7EhQGhn8hYyKmRne6pBlgR+Iq/lVIOJzyV3Ese6Rv9x
k2Cw4bHoMVETOPklbbCHMuGghK5xKu0UEt00t80hdmu38sdNxhrypO5tDuXsvowezmA9XpisJVTR
lq24R8bx171kbcBKlw7daDZou3rdJEmVnqGwvGApv/BX/p7TUMGMb9ToD87CYoJ6yoO9oQHND0gn
2w48jl1vtpm2YqL3Y5mjjZpZ4QG9CQivzDdILkNR7oieYwG1tjAY6AS0rddJ+x4IxAdvE8xSOzN1
G2dwQBcGVlmPGmtSr32eJPHCEKLTTQWizBVdTjbbc5y1Kr6ECc+2BbvQeMeEMNgPleUbfU+zjzLY
0JSwagzdBYbpLV+SnN9rW+1hLS5fWLJNLx9y/e+VQ0VTUGMq8VA4I4QUhN8BuU44dCPuFwPOvGfY
sq4EZEcgTjCzegx+9e256n7Qt3FPeJN/25Hs3FuJmDetujVCQCI6jqkBy8KLeFPwVwuR/ht9mONZ
ztP7pu8W22gaBBDpZhW06p8GHYVyAhESGksnqeHQ9B8V6OIstFW03V4HM9RpNw//zhgE4fLIFZuD
3RPrCa3+CccFC/PRQiqQuW96F7TL2lh5MHYfc5TS+GCLhkUIY9Zf8kxKUvVPRgHh8G8nmxD0yURc
4Jr2HZKd8aPrV41YNUmFR+y8pN5ohsZ4j4SpoWgbDtooEbZe4qucun+wBMa/FsGv+ptx3mPIq0sP
evN2NiCbFBiBh5cteaE1YWpKK+k88+k3PY9ahyB+/gCJdynoxU3oK2lcZChcDhskk/YTIFowejSP
ovgEv0iTTK6442HcA1a2KOPmGRk9JBeqIjATyo482g5IkCTDAbcjxqDPLPe8kwYjCBc8qwt6V45B
MuRb9Q1Tpovdt0QeG7+1qhjqgaCgwKm/Fo+s5YaaHCqrOkQKH1rJ/BATL9UHamKLPkCdwgteFrkM
o0umoPv6LmiDR3KAWv4LcX755oIMVPqcCZVlUkvfHW3B+w4UDUEG2+WyXiMjpsYv+6b3p+oxrIjq
tQMxwQJA0Fv9+peYUptnVqTiw7HDMi6ZVk/9OhSPzpAMkhSCskbhwUylg2zAS4wlJJZ+g4yfk1W0
BkaSDP+mH+QGoLmzIfQAfFDlBhEjBZ8Lv5bkBl2PSWqo/lSHYh2sxf7JdG3+9Mfooe1cpc/X/77H
YynxRkYflIbZzjjR5U8bYwCuijUJ2rlELDoz4p8u9D5AW1KX+W+/So97jLATZmFaxhuyPVhr3YP/
BGvRPvT7jg29gz7W7RGCkSW22AS51dF79CiqnTkm2Mi/k9S+UhJdQXzL7RbuEr/1g5RszhV0iroR
XEZPMp0YqeRfuVYaWcoKTeqoEKdrOggNIyxZcRU+MHX01LM/U7Rt5c4s7tVQIr+9Of11AxyhKydX
0N/KRwP47yuq/TeeuEou/Fa27k7G0qCEDc7xnNyV5HcKinPO0BrzR+DRc3UBDc39ch/+y4T2DtKv
Ael3b5U3mYVxAWqXDYVi5QG0rNaegi4zQVR71E+wIkbcZLFUPpICjmVKMnQ++7bpwirzrJuqGDBm
x1UpdBxjkOVZglGce6vGH/ESAS706q856fFp3leY5ZyIDQCOSCixtcLfmHhalSYLkVc2qidoZSi9
DwIkDhnMc9+ikqiB3WqpaMaPVhvKGOudRXdDPDA+RMe/Hyjaq0cwebRdYw66hcXO0kLbiVoKnjOm
tKu2LSMqLtD8AMHY/9K2lFcfHJWWQWhXdYN+9X0lVjuQy0JyVJlNr4tD7fohTN2yg23WtDNG5XYw
HfMhU2nUrALIsRfxSQ2NddK4TENt8pNY4xVSslWGJQ2PEr/E+Z6RblLvsc+qDX6cXG+kFOd/hqqv
6A0WY5l8UnMibMKsdOVVjgPOLSmqePkhH5nHi0yEhpNlN7CKLBiPMY4WizRp/lGRXuYcWe466z0r
s5q1008pJ90Cywq78DWUoXzwH4cYztGb4KQ50v2M+z8mGPE46E12QxIariWov903t8nyk3b8xdWd
xmXXUi2jhx6nAihnyZycNNCmx0ViXMI4WbDj+8mTyOgTgC1cQMesC33Aw2+wTv+gMwtyyztFkXIL
nXKt2fX2V4QsqTh0ZsWBeQ94AF7ltz0Qf2PQSfHUa12z7VMorfP0h8MrJfx/cHTtOVtClqUfIkCO
tBYiM6b6B6NYYfvaZcKSPrxogXD8Y9ky+3kmUZcsIn7DJJk4VTH/qW10jVeiCNwG990gjmfGP+20
Ybs8ElSafrG8BFSlgbRw8bKotLX9mssB3AfFgj/MJ51UaTMHG5FCWbeMaPSrOdUYD9WQfDgF8YwY
dd36bNmd4860dHJvBnVheyqEoVwEdLOyw4JAiFXI0azHvxtIOutQnarazqDe+EeGYLQv81GA+rp5
BhJH40whVp8o3UF0SCVGi71DliavRBmUC6UeLbF6Qzx0/ltCVDkAvRkBdz87LORgzAOer5cq61xa
H8LHNjdi+UQGfqsua4jVIJZiHxVpjXLX4pLJ2I0f5j5/QyX1Z3Mk6xBfOVJVd1KCYIPY4R/FUyWj
q3F+BIYoWjTvlqZRqM9SYLR+QGPK6efWmDVKv5fmoj3gu0Y4UPEnxlUnDO9JwomTnJVuWGTKVkdy
HdRVTPlNhSoCkYI8KG8VA+cjQdQrz6kifAyGNY992fbp3qnKZMlcvB9bi5E4R1pe+j8ehGwXwXM+
lw/VZQ/ogYQghwCHDWcTPGPWGZ1tLoBH0g51n/wSWY5wtyS7EJee5zDjZV/uWOGsFcY1fD7L4+iy
wVUcAM86NBT5EJh+oIltoQVM8nnTVWmyReD6iH3L9wYLYhFByzKe7K7Fm93cInInfjUkLmFtm0n6
DwBdfwidijZtzXuxJLretrSpBdpihV/RpofZZ/j5r3eDsSkToM3euvc+igP7fU7qlbx86sOh1cXF
CmrDC8ITaNGPYPPb860rSeUmuo5clGP+pXg23a+Hm8ihuU/+u6UhlhyfvCepiimknTHynMUlDBAB
/u56KMzqjSTAUWWhcZGDPxWMTW6CG504cL+u68Q+ESU7Wr9WAOyz3GdWqchMXpcDQeTfTjHwmaNq
NgacQgtQXe7EWeWtfkkNoHmmPUtw/RZDYjdQoXU8utohISIQuwHWwFCxBHOiBOZYkBe4qVdMhZiC
Drz1MPWr1avmlMc0LAQohBEO0pgOcPzRajnQTppmecsFzb85lxSx4IhZCsqKXFVCpFBMV2XcCKbT
VovNkFOuxrsMj5+N91PMIh8oX53PISZwgyj6lWE+xdSwRMCt8pyTyXVvwN+uu+xP31ULvGkOUNXn
UfWN+0VI5Fpp71wuEeKm99n33xhCKlDaTbJF78BDXJz6W+4wXszsftvF7n8OWFVk1pbkeU1dUh0D
XskEwSi4UxVP3HzWOgsvoXwOs2ya/Uz4oib4uCbdqbRFuHy06dL849D8VdHnq8GnqPL0om+kxlHy
EQ2VxvuCJxzHLKItYYCM5kyZoF3jnIv7ZGMf0fzDjY0ZfF7KccX6+C5KQ7H71Yuzh0g6iqnozB51
OC3WIIVsOiwQk/bXdRAaUq20QEVCThiKyfmIMFebb2nN7gmcHeE4B8yftsZDw8u7I4YMHKu50+ti
d37RM+Xc/LzrV3CA6x3T3ajUbvZqiRBPvro/rsFNTcXNxdL5lNLagOESHnfSwIOG37qr7iHRY8La
FZQZjZPKfySHgQ2zeurWHg3+eaoWb8J7ue99kWAx8BwCIGgb/d0q2BcraGg0/BiS3Ktgg0lgJe3A
VZabW1ce+1G4EixmRyMprNMTrKX9S1+OoBw+BgcnjJbrtQNV0V3EVopIBkCZAVn7LWO3d8LIt8/M
a9CZKnZr88bAU7BMrkQK7ENkzuorOnE2oHOSNkKwXGqJ7wJE1rN2MyrIbZlPF49/AuBLdsic5Y4y
cJsINp/TY1Dlqp6hOBrGWcR272ur3KcaXLOxA+IdEcsKDBJdRkgfnCyfAjywhW2+EwEs5RG63Bhi
z73hGJObvzOt+hgEUrRT0vcCOmYDfT9Q0x3D3lRWCwgn0RnGcR+Pt6TgVRUC88PvUrTuMCa1WdRj
glHqKL4nJW0qW0fw9vkjjtRJBF2XaYg0I5V0QIuz0loIENolPouo+vuUxFhqzNANAwySwb6PMnq3
WdHjP15yMBrftolCuuprR/5tLwzfLT/h+UX2J1OGzufNPj7ARovzyiZsthjRznJeuMBJpXTQFKn8
omg4YLkquVFomkzT8JQXgy9Q9GP6rsQVOMZtCCu5EwQM6Q4CRSrMslxpb4T2TFkGH85z+UAKSjq+
ook3YxAJhxHQpa4RMeP3MsUzZ95sDlNsAOixC5MyGliXym8qh33Q1Uz9MEtijyDCh/trXT2RCiJf
oT5DJlSDNFLkxgjbrLURfcul3nRnPX0zeEaVQ5jhGQNwHqcfW4BHh5uNq3/TOmKnoiMD9z/Jqq65
DneAuO7doyA4d2X8Wd4+fHrzFeUPhscaEzcl3LTBpZoLA5FNxr9g8jZUdgvKL6T8FdjScHQ27TH9
6ADBSQAZkzOVX1v3M623rsACUzPPEGe+UzcPCxmPueDP9tFlcpgnY+MuGJJrCqb2yw3cX1LlKpKT
84zNLAEBy+ELz5vLuTZdZtKfnWCCO4kfKppr1QI/BVtgp4u8Y0sqv8uN/CGvSTeHxNrxV+0NmD7B
wmsyN715GH2TgGsRaiSeys8S5XG9SkqX1SU0EBT6i+DNyYwkGvmECXx+8QTY8BiNOyXd5Y7jz3Qp
0nao9hiL3UgzLtj0CCUmmWIvNo4i++AZ232Nx2IUAp/GWwBpm4GWzPK+Isbz9BN7Wdoiuk/y0QzJ
QHgnBv0WJpJuTD9mHhZIyCMb5CaLXhUPl5l9tzcPz6t/lkqzvavHXQcZ7s3aI1HosZa1z0fqxLSv
skHkAsi3RgsqHiBMcPPaVS/hSh5MjsUAnU8b7jgn16ACH3U3aHMsHPrg7ikvhkts2M6hYqkqT7eJ
zCAxlV6XFi+vecRYS5lLZvBPCznHHRwFynA2P7U0DcLPArWxJeeutHMLyU3MYeMS8J7BA8Jjj1xS
r16bN8vonodoMkppWUWyhmEhvK0g7gIQjgNR4Pou2ZOlWVDjh2nq+F849TQ3q4N9l63hsKH9xK4r
OcxjHuBsfBDCW89C1lhtJa8TLwQFWnQKxvI0lLnSwtkmAqVQghEvEjJxWYQZvPcT5nmQfQQ3VO1q
/MOjEM4VS5FsEVgR6ZMjfUnwmccxSsGlEoHq0hOOu/ht3+AnhjcIL2DLLRATCY3m8vswijW653tT
+sVlSa/hPWl1cOCjvZ9WTG6WVqVTxagQnbMsBR3NJQe/FQF0ZXfUYfuv9QiwIBLangR1J+Iy8GC0
VTin49c4Osb5rcra8gwchzAKuRNQRqJE13aen9qpcOFjAAjC4+97llYmR2hEPKTzuYoyz+qybjTq
HMq9nRDTyCjGPj9xEksGvM4urHLOJiVHBfBiUkLSqa+dyxJEmlcdyIJtMcH7IdQXwJPbYhu6UhEm
fVHustrLL7W7UnSGRMqLHNkhirBfQ04PgETXb8DPYdUSVRSvnJnfL9xDaRP/tIkcgAaq2/dXrB2T
gFed+YrlPX9CLXI4XcIjgDg0QCd4+M9rNWxVEIBrXAI6+otP5cxwajDxSL823gUtrSGIOkgBb/5C
XZrz9GFJG18JUgX86VEUrUddWwxqxlCqjwzO28lpuUkKf5vQUv4bik8lRi3AlJTBG23CEl7UzmLK
wMaZQK39V5BgG/ilcvSq0YWU2Eq6FLfDguNFFufSUgmFz8/jJ2NhMnXzHNMyM/xo1rteNkdXk+nf
NiiL5zWW7kAptqeOEO72OqWJh8OO4Lw21jB3sbtoIdMRx7oDuuzuoy8QtjMF+kqujZJGcuMByWl2
t4zyY1an51Yx9fuq4a+jt6jUrUSfqKD0E3FqcLfmoEnzXNcdMHMf7WBvq+Emt07Y1hzhQXz+2ZRz
oL7WVMS2BeVa3dby5EO0zRh5myRKRt6mD2axhUwpBly2ZIHh8UUTUfEE4bbpAC/e1VNmzETJEEzr
PjMLK6ht034L/34luZXv8b34aXnGbXFU2tNb0m3nYY/BxHBFoNL99MH/sV1WiTo8lRwWhjR3Mppx
fFqITB2KurQeqr+G1pbvzS7rcEF2f2TauZjLbKjQKjWHaViX+RHxsXUzXfe3Z4KeHAYOO192NL7a
dI8uBx4Lrnz2SOStZZ5WFpfiyQYc2+wAQojxC9IP2dLmvv9ZtsYOb+TOtqEHAjyhqnh//a/rFCc5
5OD++QdHUGPKjPRyBieVB+m5dajhFTRAcdoUPtbp1TMn9FlPqdARRcIKVam/Q+o/UjBBLoGrIKfU
GPWFsgyM1PttMyK9cfS5SRe40wwoXwcBT0K9ScVbU1V2ccO15Y9DAX4pSECgTOs+mq2HgfI56/il
fZlX4iIMDN9e2U6nGTdxz1ehQvYjR73A4uMENPcUAqrXycH0kzMyFcDYopeGQoYW3DWH36xNrWpW
n7We8fPHGZy3NzOreRoxDm1HnWblO2HMuGRvoN1EpbgVmbiumqBpReDnY2ouLE4lsvvbojvcdX9M
qzFfaMbsjufkoBrtjqmmNcvpiRk1+zXD5eTN7AoU+zBXEdkgJqQA5nqLJj9Mcq8OMbAvFoBDxxEN
UDcmnEGBbtXCWq9a6qegq704kdixIbgxxdXViE85AqT4jqiaznk4FO9wEwIWio4Kzmq98jB1Setb
3sStTOSFq7+FxNrbp+batAGbiJ2E0B4pIR3HvWU5a4vSoxZtgOF0Gorr2fEeMIiFYtGAt72aXTEr
/f8oVY7xVEK4uDGg498CHkAShjmlRhUGU7eAaErMky36NimC5OyBMRogCYjDYhh3tszXsTFdcpi0
QNYFkhwxvxXAAEiSnFZhHfFileekV02FnF6uim+/0NtZTx3aGP09B2vgU7RpC9bK/NY9AqXoXyWa
SeM2i4rM9NR4rBNsIOUaiSmIMDxUZHQfk5I/i3zFogGXiIIpNDdb5SbOhjDKv7FGefpDLn9dVEV8
Lxkdzo60thULKrParNZYZmBcVkxnT94aURHBD9vr65gv2a5ddsySO1ZddvwC40c25/97XXrfjtnB
WdZfxfW1nnaiFleip1XKtDZWQ3ZNqG+0yWBt5vpQnvnc1tRA3BBD6Yi8sg0vPvqqRyx5W0ihK11v
HL6Lq3yyiH673/+F0ks6+tXTahHAozbRyfCpKLqB4/pWNS0lRWxYRoUv71bQfef7d0FmYmXaqdli
trPKSln1zfXD0sPmT6BpStyx7x+u0Z0YpwNSHfb9L/x8OngVmtw9+2yLOqs6rocOKqLObeGLrKHk
PHe3V25TJuXS+VCXFBcdGXLXPPwFdi/fTkJ7XaXHcZzMQd9/hgEXXSui3ymLdV3HZO17QPPZpd7C
8yZtU0ww454OdE7qiWRMKLSNbjeuwF5+6WopFVh4wpMyoeHFS2pmDMZRWOyD6vvkW57ba/OulbaC
flqGY2ma2buy67tYjTQenOE161VkHdSLnSFkGEkX/zHr4VZiEsmQXuELDsO8EdY3dyy4BIik+xPn
YrJusc3JkTAiSaYx0QszNB1zXdL6k1SJj1RL2v46froYQjTl7pwIW54Wd2c6w+D6GeOcLG+ERQSL
noYWZRJfnfOrUOgvgYpkMkEXnIQ3gnXswVAsQn7EgQRRKOOYLsTSHWVPy8ey46TTyqbJUoEjofho
qS0wUUYXR1izYscpuRqr1F+027OaXKQzM1jH6Q1BzBF3jzmlQoKLz2YlID4DhbQEcxigaLKQwObR
XpcjAQq7m3ClHvEWUyupGKTHp9CJSwE6vQebt1O8RL1Ki24vEzbPmz/CljUUY97jPLghj3R6nXrf
tzuJFWmh0GIBf8GAXiQ+K0C4wcHqz+WVvMo6ZQV2a0OJitI+dOR13Sr0Fju2dtcNaZbfVTeAC2On
HLF1HHY716YBB/+1yhXVNWFE9av+n4I9tmX8/IZNTxU9k4roxwaapf1R9h2P5UqVU5Cst2OPNn4U
JfBIdrTGEFoD6ogARmAXmyGpeo0aKmlZ66+EjYaoSEao7tCs/gMslCD8jVjCF1ugXnLs8AZBgOdv
SfCFKScYF6c+1pvLrXPaUJN9FzYOEKmrCLizdW78SJPAgKuI7N+MGBzIW+NzqESEUBGZZ1mJwi26
/hpC8Vghb7e1z7yH2houm33Cso16tlB7EKbHs/Md7G4h84LQ0kSm7g3+R+EhdC3il7JpHKzczu0T
Fd/AbJ9b50ZfhYbEOnnbQYK5asM5nVcmSwL9iFvOwqq6FSOTtNeVtZ9QS+dm9568abJ1ymE6G6UI
NbMCzosUS5fEPw34XOnkA69X06cpeb1IvHgTEOfBJnhcq6DT1gKNvBzZnCzzAa9k/qmT8ZfPZILx
/PAwlo9XZV1uwI9OreSEtX8pVy4ZY23oCI3GRLaeUhWPppeSCU5H4GDkoJxe84fdEFwOBkLXN+cQ
vjgWuVVmFYC6FdwIz77gK6mhqypnMrcTb3W61y6OpO79GEi60scAJPwq8tspZ7LadYb2xZfNo2o5
R9IZEyI1kEpPeAZiX3Zgc3s/uxQtWew+P+aBLCrHGHGpl/ocvrPXjnHBX7lFswXDX50V5v9M1Czd
M21raS/lnE5R+Z0A4mLMa4w8lP2xpD59Lhfk90ULZCdzL3EkeJj4gUXYAtVbgXGG9Hf0jAeJZGjQ
FWhVIVwVoiTmw/fKZmAGdCcoIvzJwae+EkdW84TCHYSnuqGTOjv48Mf1uzdyu9aVWsyz2rI2/6Vf
VYT7zudoMu3ZcSGtBjIh7CVCFB/udP0m2jbhlwhCuqBivIsu5EHYjHeFNv2ICfEqj3pTleLP/0AU
wro6pG9z+ueJRAr5iMR4CDBw5sbX/nvjE7BF025igK7WoMcWUDqUqcZDQypl6X5NszpxkMrTBwx3
vyqJdw0ziF7GTfIMrR2XcgWIOb1zTHa5hwjMmDpXsqgLfd/TNHUx+jRXKfijVzqvkbmJVqLk75oD
YAiXD8T/k1RGw79r4Gktg36KYlGoi10bLPunK2CFG9lsXPscrZzfOBocZJ9y6Ht9zdrK4q8w74GB
smd36WOjrrM7PQ7xrfZfHRogbxrWscn54YuvISWGMT34XD/jZ+sYp8BfyJQNyrRIP2pVyurPCINo
cJaXcHCSn6Cdy1NApeHvNlQX0v3qwGCVqf06hQ85o+kuwlOVawlP7Qu0hKR32pWQBMmsAhWmX023
0n6UpQvqQ1V0ZEAPfsZdNOEdQylrtQu8xCA4eq61BZn2J3vYoiGgNScTvn2X76G1lJ2LVzRNOcJn
AjVFO/dALViB7fQDucIEyqrtbXVKOGFxESieHgASptBXZe2r7Lmibhxj9UUN9WMBlPx2fOqB2Q+W
0HNeHSdKvH4pbX3AdXyscG1wznOMwI9fnWzMPZKPnC1L5DAcyECFbyncLdquTVqbJdhF5gN62PYR
9pPlsXbEKHofHmcT9YQmO5bOt5STHGd/+4sl+61+dPfYm8ikBBy1Pp6XbG/Qao2NSObYLzxWFW6F
xO7HvHqA3zzp9aBQH28rWvUQoKnhHbI2VL/2OLB0aQbs48nSvOJUpmrmLt6JeqqbVT/2CfZvt+VY
XNAvThE2mjt0T7TjMbEBYrR71dLw7pg6AxbeDwETQcLviYZ1rzmfG5eev5h8dF2uA4PXO3GWxPMU
Hp5odTLHddNNZ1W+dKOWpaGtWwqrgaDD27P3x00Mq2fEWdKj6DtvR+gz6S68WRyHvRysvszJghlS
Xv50l/NcqP5jqxbzILIyXyLtNYloNivAk6In9bWV3eXljLKuUjTsjY/s02LxFCWSEIxo0d7pF7z6
5+Ixb6sE9TMIxVZP0sGTSkG3frQDFiwwwVxvrkSi+rgGQdIK1rY3RN9G3xM5GYA/vROHjincGN99
7rpo9ecIBFnO6VxsUg4XZAvdH+ZzcEDuhh1JvG0C691gVM8JkfHFucdFPHxxioA05dcYUxtBEJBT
TgNjOwswV3Dfhws+TVDhfGaHmngCdWqO6Jz2ZoqWZTDQCCxEibGHE2EhS9jfHr8omWtcbieqW9zy
QOG+StuVsjw8cm7wnkPS2b2AOXwMW8kpIsKJSRVGAg9qaMTndV8KEdDJ1r/e7zXY5XGa79tPhe/J
sPnRfU57ixwRHVy40jH80lP03iSgngFsKqsQ2WN8WkELV/D032sGR+WLK/ROHFlJHQZZZWl1zTGT
tlRJXumukPNHETIkqL+X6c2LZ6SEh0NEaleF0X+Ldfo/N1gm3vVIS0ltRyS8e8C9EXhNlVCTMvfC
wqtNHCooSI9JF7C7FFLQnSGiy4ocb/ejAwWypbKbxoDKgN7Op85XjQJ45StyTnf/XRnW9nlGaaN4
odUn1cYDE7BC7REng2a0BlN7a39pSRollkhlCvuO4U8FNnrgqxbd4pP0T7Iz82aprcbi31cxJVR+
hk07Fh5RvQ4xGtsk5vTSTlXgpjxaeVl4LNAw9CUG8oREmMta96duj6JhiNAJ3Yyk0srxRU2SE1By
rTrNU65f4emPsmHtlhx1nJkRoL3CIdWVhAgYyaBzwC8rkl+QRPj94tSG+6oQMCcZaFyfpClfyiCE
d9U89Nx2PsJozT3gRPsfih4K0NooUsTJGmIHbKCs62HZcgSp/IgeVisuqYvouLK3LElwPGx7wERJ
hRl2ilhRitSy6PAyJbLAzJEIoex4+LF+YA3ujUTK/qHmqtSAnfE9GakKdq6fO7aqg88cULbue8JQ
+mcHmKv3FzoPO5is6ycs1f3iegO3Inz7ZE/tS2BhgiRP2KrvnLoPR5+qnkzwCIVjm+QLepwXleYC
81x6zouOfA0MUNFXZ3wzWb5i4tEKZaFm4fWNolF+/CdK5NKPBnId8Gg5LIRHYAWoOqS/a7Qriz1x
pWBYRDDNWAHGqxCTw5H+9YqbNVNm2KANui7/DQyH/K6HpPIAuHg10yY7dUzD4Eqi8y6VpDxvrBYz
gKxrnmQQG7DpjDspKVx82D9YbOwq/IGFv16ceONIeaQ6q9oPHcGRL5NBWJGGHMqh///4HigMEJCo
PyJiVNEdl6uh2DBwYv7OPa11PCRCRsQE/bJ6FiIbtkM2mGSjf/vWtAyumd83NaKd3vpXtavGs1sp
HpVyrwhI7AaMwX7lQgx+5PT0sxuY/irUBFpaH1m3mD2w8nJEFVkyCAMFn96XQouRDQZ6qTj2utLJ
PYJMjhwNgUPft04zSt7Yd3Qh8lroePU/iUexg7Tzj8QgzIILwl0tGaMxetA8bYr4kLqti7lgxsc3
0M1DxT6RZKfKgjhhgktI0CEJU2MRA6ZfxZ2iz8irkpf69HfSTkb9wlrK/shMeFzisFol5dtbVJpa
PSQq4SaMtP1JSuGinJDqk4+mDTbRY/q3kQJ7Fhae0VLiA7NV7QLe/wVnufnbt4ZsJPFAnxeHYjoh
Yx59fwqFqATcXhyMUH7R5DAlqc/YZrBK3w9mybQo3pJZUB1bv3isKRp8ccZ7ZxaAOcipuk6irk26
58Ks5/0KNWfvPsSnrghQIMvftCh1q994XmTZxgW+b1paoB85Old3zKeGnGpSN3q9Yt+lHu9X0TcO
FNp1rlRUHI2EjnjUg3ZAE27ijgXlvBNMXoSFUzLEbQdN4Ssx7KLtbfpsfkGIlRXFLcnSw45QttIt
ofnY0PVmo6PJG/clFCb2pWV+0qDwGQ6mcwo1XouOyCt22QYrCagDnLjpVBeelhP+a6eUZxAe8JDA
qfLtDFaVLW0sVX5eWHWKTnO9qYAt2ukUPULsL+eTILHlqf+3Fv+U24a1xHD6HVSfxzhQivXm8Jij
bndY+LalBMr2tnKCie/aaE5AbzePaWg4xPgXmo/Y7NSbmySt/sCmEkencS+4HzZ+59Ia8OdREpd3
ZZ6R4AboOdGHFIsUEfErRgR0+FbezstF/8cn3MaiZ793GJtwWoxKnU1GuZdg/2xvtiBAUTKPNaqx
36Bbd402R6Slm0lJPjFCDjRLp5EMs60Rxu9Rl/R+O60FdRmILGBGFZDwJoUG0WR/1B21ShdXuTNK
DdjlNitXhaCNUmg2Yq8sH0ZtZpdc8Jr2lfs6jutmFOERwERJPSm9rUZBo+9kCd0/NveZe17D37HM
sVfRMXB4LSfXlehTCD04dn1wc+ZI45fFaneS+ZeAj2X2pnwWvOXZqdjRBtKv1UJSyxeTvjxqQkDZ
y8zjYPKdsau7fbfrJlPwAWy9q+ueqstDJu3tFvx+jmXlKzA+287nWTuHyi4Du925ZpFB6o/X7C+m
aMecUbOPc5PN3Gj5GwoSKVDZIgvMkchvyb4xyRmJiNJITNBN48PeSUwRSjrI62rR3nSGKzEF+kso
ZB5FztAvDc/lRhNhJWcMY+uekhe2r/fFwJqKWk7tN4sVQgZYjdgptzObzPTIiD8Fp8Ox34ubAKKp
86lenQ+1P0z/NiiOiC9UvoYlA60AOIWqsIzLCayvuNOVa//wDo2Mz7xW7jjC3EDj+sDGH97m3F96
gTnsfZMuAr8wwSdgIFjwZXc7LzSUysqxotRuRlxn8LwdlZXBTEkCd0+u/u5YZiWDI4sZZshkCkRO
5qE7dEuHGJUugLmaIEqx3VTmnHb6DmU3tBFXBU61P497pQ0aFj64G0T02/C8jLbr6Xu/jT46FlD4
b6/j6xHdIaiU2l8haWQx0u0KrHGFdLklPGigGQuK4Y6MdgOS0+v0HVa5ji8o8vpyDetNZV47Dkyu
fBenx3dTuyK8fnX3r2ym+ETDhyFPjgI8dTDfs7O+N6SbK8LWOkpM4zMQFAM55Y+yn2g/1jL9ZXPD
9xFOsLPKFs80TLTGKsT293Vv2Jf+ov0P2xbuqfWZk3aIheLVjmaqCQEf1GK3I1uqs/dO8Y21/j2l
qDWtP0M/xhkE+YC7JnEut11/8WHRxGK2e4oKep4QNoe1bR608Wm89fcAUbM7tyiPuwx4ihfIOhVU
WCDZG04eHo2aAa5XhgyfQnj7qF/tyN9GR/bGgDMOnOemEsYu6yyslLLH+czxILzTUT4kZ70c9HXw
n6EzRMUgFbFKYWuwdD/rfSUfT27FNOSwEg71f7QQR7ypuxfq0g1aYpQJAsbgsdP27DmpSlNgGRv/
njRmSe1G1oDOo/iisZ1nEU1BAQOnUC7GdJRaEYa99TVQiOUqi51MdkNLi3Edawy5Wk9doCAgT+9P
Vva8mXyWML1vTym8RJA0cvFecy47NywnaPCg/JFc1jm3E8gak47Mhfu0V6cn1i7QfMN+P5ggxyNK
gUYbSDRM1SQahXVVQzUPtHWGBxTiZDWD3jyTzfaoPcMHGdR0Bl0/E0CD/W811P0Gi7uIKpxVnNtH
UwIktDiclN4tJMHJRe66XJrxjx2uu6+0tlJupIuHicoJUa6pdM08yre1XuWnDZj6PjNPTDcUbV7y
EfiO7u8xmQhku5vNZ0DdGq3XAsrC1080wHFrGlnArSi3U2q1ocIMUJThkvXt4YWIQTzlmyNC9afN
4waHYUi0zW7ZirI8haSae8j7MrsxjSaCe8HYuxJ0GquWyzMSIPIHiyVmqUzbn2zsS4JFHKMkMcWu
Wxg4QYaYND+WcqJQ2GHOGaE84XUkOVx3uGK+4ZzW56gWoPQdkG5qGfZmU0rqBZlsPALYaaO/HDBD
78eCZ/IWZLWGOw5O8/q5GmU3BrjRxpeT1YX33sbPWBjZkWyoDcgrwVKlQB+T6Tgj4ika0vVC5GgA
flyptG0eQh6RUdYoWtqegduErzCHA4wvgnOt9VFafiSezjih4/xkPg36j9bNSSvqjZKlWyczdZUX
f4OUvjKpWLOP24/A+mt2bhz23phUHq8yb+C3E1WuazRXxT76XZA9jcXDnxqQGt4s8CcZUV5g7EAg
mRH9fZrrPKX4Em01IfvEJeAooAWzIS6SS/D6zwwWd8cwGYpsgnsULuv912V/T9Izhgm3RU+JqTEM
O/LOqi7NO07mQgsdxXQbTtbMrE2mBYm7K5oBLmMkZuUSKnymnJiOK0duMUEwy1w7GWVbULfo08Dy
oQ9Gfn9IYfCFrPLK4gOBmmc34/9X5rBTV+84MIIM1MBlb3yOJpvfFYGD0730T3suYDip2ZSpESwZ
+cGOQomJLeBqtNQRFWgY0l4CExz33DXWeTW+dySRSBHlr61Dgns8jzFFkVcFfrOBlyMzR7j8LJeW
3OygQPfGQ1ARqiO3hw0KeWexm7JP+tdNDGh7CezMprhcujCCvxtEwi4QxzAVTgGXKtaSZMmltbFt
oGzWlsGIhPM09Tuf51enO2g8DIdFeHeN88gqESm5TQyDyPFIbqQroW6Q5krHQ7hVKWVxAmUMySFx
dXwup4sLUkkTAxad5IqQncAapVCB60mf2MT5xPdRmQfWQGE2kGrIZu8TtIhZIN8YuHRJjPxQ/q8a
1rjmJuzbtPbwDqApFKaeVHuT7pELWdDxo6xkIy0/1FFWLJuG+7oxRLbEFY+1xXuom7Dyg6cRB1Zr
CUwUNAfmOQItBDSFkwowytcF92BEFTiod4dDWEVU1gbPryRUUxYk/72RO3EpORG4nwLEzzZfiQoA
sTJYCLQ3IGPqGRdgTAYegodl097RMOKsCF5vXaSxPUH1UX9JGKk+qzE7RHDXZgHPCUmCT12NnCfW
DH+/PHRr5SDX1pRjNyJeN5aYUpzHdJU0972/2l3H1S4E6/lHlHUggZOV78fe5KijWkx4g2xTsPRv
O1hx5U/wwhwpQLl3ecBRCrDVmxa1MQiuFiTrXgEt5LY5fUp0KIAfLKZb1BN97n0RciFGQ2kf3cRQ
8TVCREbi8+D7ilSHgRVl/WKgswl5RMVA29aVHu05omwJ8Fx1bbWWhjA/jj70XFbHm8tK9UD+bXYi
IxnJrl8ILjnQNWdDDmwr0FJbsEb1Uv7mPRvEeR1UsR8+e4WINqUVTCHGvd8GxV3iuY5l3WPLmuyy
MjwcUXX+jKb9aqxB/OapbCIkgXuY38l17K8lIlegUThUm4rI6xBy6NlvYnti0cgZiwYS8Bru7ZAC
vmSCMsV4NheF2MrFp1fratYk2EVRfAHE0dvAjs1tOsHzNUdQ99ruy7+WtFBtYsHeq9dv1zkGBjap
4Alk7jWNGW3mrbB649D1jLR8rvUb9fyzw3+rzHdqORIUzH+Kb16czoOR1oCRtZ3S+G5JeHbo6w8d
CWSqo+/vL4CfRdVLvy6/3q3FvnPn5r3Q+QCW28s8E2BVbnOyPJWFGjdx6OKwaNgYXiWn/Ddt45Sc
Zc0u7bEQ4ops5SXIrTtGE+OTANw6SXjrIHE/ciPNBAyVauCqUmEih/r3+YknniHY5Vh/shpoIIBh
aAuPWVYwn6TwoPXudFpeAnd3ErOYqeywg9uO+WKbj0Q6KooofUSMDZNEe+FaRcMSGiEv3Udp2k91
HV0nVJi58ic8XCeLc3Mu+P8S7a8ZK6sbHVed9W+EOkJE0SWM8yOagYZIlb0j3zFeGPL40/7Rr5b3
clHJgZTOzfmOmbxHcrBu3COemfKn4g7OxK9Z2XfVTAITpV3b6vkHGMD0hBla1aJLgUrTNYNBpekD
1mpkIdkH2MdM4iIbiVE9ISI60YdtLXD5eBh4GbHdCqEKi+QMZP/IebHzBlzGvNie/NqNdJlp5fhb
jOgP1mxtdb9Cj9LPS9i/bXegE5gYxMqMvMF/adMOYtdm+tPqf4QN+D3DKUfQEUsvtmEP+c+EjJAI
HkzvqAsP5te0R3MW6MISg84BPvW9327EksbT/f+Mg30Uqar9MMgytqlopq6r+ssofGnN1YU56Ftd
7qT/+Mpv9uZCnzRRS9S6PJ4jN6sRTD3jM5FAOvC7aVVDwA1sUw7dfmYQVUmk16PK4C/VVYf5GwxC
kq/VAKdzTAERHnplWs3B/xKyXd5v4Sr4A60dTC3X3xMoQF34Yb6yOCTBD7apOrUhS7623/aj2Ydb
3z57KzOqXUb2F0KNpJIm9M57TZz9IbTcle0XtwoGCAM5Q+OcxvJn0zh3v2JTFRG6s2PJPERI46jU
iLv9G8jYjM39642Uu7GBAyl4+YGeG3vGRHsK0FMCJouMHpkjtikD1he6SzkBvGnEP9Xk4slTqJAS
lK2R2RRQi1EItViXs50uheeZ3ckHgS+R4ciLw5i4zpzLSjK+kx9mMOy3uOOCkBV4JivJaiTTpOi7
fXE1QcuLnb+YzsvwhCb8ktKM8g2bpJIHixZwzlhpQZjfdCdZpV3DHlwV3tHUZP+GpG151AZ28266
jtcdoP5dIaiEr4LCArPeYN2fIWeHVzYiU8GRHAbo4BlU49CSxjSxzMEq90Q3GzQ8WHIqey9QP85g
mG98tiDd8unO9jlpFDVHkMZOd7vyXwboNrgMkGmUlYzA9sndpSfd9vGsHl6jF8iEknetgP/qAUty
yLBSsQqAsD2ek+9H5AL470juKFPaSOONVYvZiSuM8WdIjoQdjjL/bxLsa9lQaIkyTnjwx9hSqAeO
3HXw2WXR+a7+KkDqn/SjwKy5XRnSKJLTkLaCvgbIHD3hiHIHZyum3HNRf/61KeaXKzI9gbVQjA90
vk+hWJcp7qL3tRv8BXm6VB/A5AEFeB9axDIFSBVIi9/s/aaup1BRUgo44xQMVYci6QCh0BO6d2If
OUTO1bMfvhljSVFx7F9iJ5CP1HAT2LAyTwUJFZv3yfnpXNaOYGwD4soT+eM9GuI/sXBsSnLo5k7g
t933jiDrAUZlS1hmskk3PmbFjgk3YvsIWUlk7uM07mNFtYLzISsoxshKHAR7H1eWXUgOURTQHj9e
VzrDdW+dwMMUDtwTsbKfSaFzzzTDEX9Na7XsbeF3Dv2tTW8emfl0/E6ulUC6kc2ZVgljN6JZKXfL
fArLfv9EVb4+PwOaG866un49sUCgMvRzQLhCBr0Imay7+DGU9vs+w/o/eJd8aVCTf6WqGEFeYcz6
/8ezoDcfiLPs4vVGugxFIY1eOIUaCBcjuZZ6kkxspt61GbczBr3ZlkeQw+FOeGwF0mvsCtxGtHSM
akDWXZ2fot+6JwbYVdLDzC6ZcJJwRZ7VQZsxmhAZ0tjbHgUklGEc6qYtnwm0kARQFxb77jzUIh2z
0ubrx2mA2OhIxQxlyGlcYDNGmdIH/p0WbVfQiMHntuHqnEEM7QSzf2tA0dInswGdCs+jVrn1aaUE
1cZCaOIuR60GzM/d6M0E///JqjKNs62Jx4Vq9QBabaSjSHL0Ru5usUbjf2kNLqQsNTNn46fBoNkK
OFaQoziMyoCvCSQaOj/THmyKJaD8C1N/VlAWQHEyBVWtrcz+48sGwFJ5CuMHYVpFJizC6SQObJWV
nZQ12gjz7cOhbp9fO+LQwZUdcsVuZQ70cEfrQvyACQhh/PdAvKQ2V6/L+NdUi4Wafvg41eAfnIlJ
Cng3032FcFxdpK2zpMpyi1oLyoIHl3fU0iSBLnNkY9BDWKUX8uzGimNYmd+t2WeAGD52evV2kmkV
1rVQyMb6Tm7VlILDi2UPZTkA0Uupe6M4SpKrKVNHJuLd5hIE+98xCkL9B2oBAW2n1izXGiNSRXCg
gyXYMYuwQrKyS1O99YEERVCqLu134aDQZ7tz9WracaCIwpa6WhmrpmVZ/hViKXQq9hznHk2cuVK1
t0her/Y+C8BC+qvBMV/JUz7ngGGkKsxe0VmliAsGJCRk2DYHZbyTGbvhAQyf9cLrfhMz67AdcRC9
osCWNhAiZL/tgeZkoPCPxw4QOl7PN9wD5C+iGVDKzrM0cSdyn4AA1JBeCLCALHfm2smIetDz0D+B
Rnn9XRpED7BvuaMlrk+eBvHUr+779uXEBYEx7VXO99CmVkKcr/X0OPBGCqhQXXqfxfbu2ahfQ0TS
tpwbF7owzRolPNmZzb++L2WFq5T6l95uq0BE1NTCzdTF7K/vQ8aXc/cG/ubRmtbl2ZMohltodXUs
10DZZJzAKC2Mwd39fe71SDFOk5KwZ7GzkfS25IM9cXCLZ9m/00iBiYdkCBVhkl5wCQXVi2+xveVQ
Fz+vjIAp9M5XdedNbHRiWNOYnOYEzTmAnchte3m0Vbv+CPq7EFIGUrOjUpJSleFx+BivoAdz0d+/
7o1xprGyO8a7wnRkP+FyXwnNl66dx9OV0ZdP9lTEOkAFasqarP8uqgSOY8O3sDwn6x8fofy1RWKI
X8u79rSitBxacdNXVDpU5vrcRl9A/C1u9nB7de/0FTbBt0c5UvBGqgyH1a1byLiuQ0MqrHs2m9xZ
o+xOqZI9tFBziCAQCN2v9+ZxOACJTAtU3BtN50X3GHI1GygW2Kluy5iLuXzwzghz3kJaOG5n4aMW
xcVLb4BaLHoQaXRN0Z+9cFn7qpffKgp7Kus6HFmYmfZgzEjMgoWB6ZzVtJD4j97GzjoaOgidgmKf
/0JGOVeRlVP/pyEAfsNOoBMiEJtWlV0aD6qiT9TG+WnqCfdQD9C3OUF6wiaibn9Afza8UNnAgOTi
W0ycsdRK7Qp/5QxTRk1ZQpf7+xrs46Iz4CK5kX+qANY2LJbnXfVdflX0VfOCl/VD7Az5eF4OmFTo
D5KY4lvuzlfzuz57RZmscS5Su1VYIf37fHAfI3b5gW54AP1fVNpE9zQO7azlKJTzAJN8J736GCCy
fASKnb/M3r3DsHLs2W4c9nlXqU2MQvw/8gTZ66FT6S0SyvmPpsZ6IfqaTyz0sG69nhAptIoiefCs
SDLMs4fc0qozSezQCKEMs6xjt/GNaiKjJWUsQIYR6I63BkXsI0Hb+D4qoso0Nd6CY4M22y2vlK7S
M9BAPxRfsuowI4yHXfQgpTwTYEreExTPUZ7pZvAxqBiXT5kq/iJORSPJfHpSFDz/40U/9iXwy/qd
/QCXzLf1Mw5fHE0HYrlIyQz9RlAd+od2VwZej1J3dcWz6x3POP5fR/MLEZfyOah2hdyq0rI+wHKB
0qzTYHPmvGc2GbsuzbxEG+QIw5X2h7A9Q3a6PaL7+GAW256lRPCWul9CJ6Wnh6g2y7CMjY05UKcY
I118U9t6vKd/idNK3n4adtERm+XyTVu+C7Kbazmtwez+nO3BTd1N748bPabhCdty+RGh6gauSUiS
kd0o4rdWyQszzPMIOwHhQjL2D1W8pQn5HZ6WfdshMra1UImLvyxoQi5oInw37cTwksojzwo8wDYn
3wKIsBMC/5Go9d3huB4YKuS5R7JG2a+JERRdjzAITDJF6vF5hV74h9Zc/tXpo7zLSTlnpNUDh47z
ZNZN1RU2AVdY7C8yxb1LyR0Dty4iFTNvdNXVbewAD++PNQpV3SnGONj2IoSxQ/u0auOuMPwBHmu8
0JewIromvx7hRUaodBe4cfnvT1uvKWDiG+FMMkklxLE4lxg1S6U3rz4ja8MSv7a4J6eCz7nC4kmQ
HzCyc3+lcrfHkE+i21EhHBp43WNZ+aXIOpCko1xecS8IY2mx9s/gVzytY+R9etskoZmw7sPcB1rD
ylbDAfuBB57TMifC/6z0/1wWjWcDAJkJDAb020iKQY1hwB3RyHP3C+uAMQyuzSFsI+ONCEzRvBwy
mlwtd/Tb6yG8/vtsr/juOg2w3nuK2fS8cgcmXutnMcYsvxUl8vv2KlUYfty/9+RaR2CMQAFZdOVa
QWF25udVdu0otQ7U1C8AApez9y2rR+aFKAUnXoiNB3ChYgbBjhA6FheqxNd/StBOzAVfsHrq0dQi
4HwZFkP7tQjl4rO0GFdQ8VJQ3MPyut1ZS706nRrdR/dse/4G8gf62DxH3mME/mMyuEqfF/6GfrcQ
gwsWTbygL1Qv2GOcwJtmVfDyONiWhvsOOn1VBGwNXRBFoBWyJRfDrjVhyCu/M+zSkSLSmJvokI4O
2l/81c1jRIH+GPwDGbZOReG26pZd7Ee30TSPlc0FSgYVQ+wJT5mRB+aeYsJncor+64rb9CeBTPyw
ARdfS0o2rQSXN8Rhsjxg8L5DZ6a/0TZuJSMuWIjo6kF51IU3bvEb51YwkTYQBSYJ1GTBH5/RWrDU
yfILnUCn4d2uc6Jybw/+8AozAMashR5eQNtRDbTTnbezjLHpMhupn3NxJ3W5Ce8ODDkXMI/K7Kuu
6mKVq6D2ve0WWFZn3PaHb0LA79h8dyPfu+rpgMsqMCdXEwgfGsbn7pjusomch630rm6seO76/Ji1
U2dkQ1dV7n9mVRm3KfDXrCPAPVrcj0UBcVbNdXgAAdK3qugrMAYTkiIeyfaJ4TGNH7uA/ZkRcXAb
uciDt0khGNOwwFPHQlWAbm/f48+9LrmSXQt1bBboD1nHIMsuB2ymaHp/TEkMHPndNGOlamooHbr8
Z1cmbuZkHxWTHE6rLQF2u12yncOpP+V/Hc+blgC+70mFSBSV6Na4JlTdszPpSc2dCTOOgg6qpAgK
Pws3SBdND6fZBrRHJgze6D4oVavkjtryiNz4X04aN3Mlm9zgizs0YUq5zUqlntD+KZuPSwOfKyFx
d5NUMvJsZTBurMcl6lCu2msw3FFpAVWIugLLALcyHfww6qPuZ8jAF6Rh4LS9se7YwE55T0LjgAw7
uocCEMcB0SiGQnCvaqjEkAFfUAZ9XOJpyzrCqXmJtj4ifaHssA4TFpGhctOOOP9W7UMmKCaycOv2
kODHQfNXJK9Ys8hWqymX9inV5cEz7m6slolaLOHPE9U0axanIU60QnRvmu6uXm/dZ9r8GKEt9Zje
ZZ5sbvvV55hVYpnCl8fRJLgO8jgi01X/d5085twaYtzU+3/3ch5bJaGB5GggAE3a4gOobD5jXcdx
3zeS2JcQ7FmR17AUDcjvPkiRyYnAiSmI8OuOEmNJQKAp1e2uBdCgbVPh3jgPPsZk390hCudSm9zs
96WZailOfbr3ouwwobNVhw3QBCs0ni6GK37wj6MInM3XSvKNFVQbAO7NGT0gc927gEEUgVZIiuY4
K2gOTdNICaltYd+m2jO0z6gexFCnXPxaj+1DOKOdtBJNFTKs8+oPZxo/FDwaL5UwCFlq1jECDP2k
walJLICAeDF+iJ4bomeWJH7QAnhYM9723iVI0wxbEOwWAJwXXGswQrdJ0lMgkgi7G6vUEKTWypcN
bHh28cnwLA/DfkLpQ95lv86kMLkU3c7032vb3SBjpYkfgYOCgqoh2FEmdGS8PBXh5LqOIdMW5kDD
f/+qxILrE4FtPRrfqEjW5uKSeaApuxZyNXeULmPkV9+NpqI07ZxmK435ehAKcVsHzuZF0dCaGeQw
D5V99UyYTAMGP9akXqSTreUMe9T9Q5ljiFEqbGHX1EiOvZ2E2g1HWkszRYGPfU1CNvrFkptqJjjt
9kIBc4e60cMxkkbv0Z9yHvdQBZZ2aARQhWq8ODuAslia5lhxuoDfDM8rmeUuDfguvtosWMhe+kTf
XXi7WXxFf9WjJZncvqnZRCa5QvuJP87Tji/kJWciZWazT5mzhMWcGEVKBoE5SA1EZEzuTjalGtUq
/S2a+JRpg5mTezaiwqNamx2ZFhrt6XVS0JTDXpgVnyRZcP2Md+kKVdOUPW44JWd94G8ij8/3zLXV
KBeX4eFxXRY24fow7gMn1JV9KMw27R6pz/B4aNNl0TtukbYSFh0AwpQuMWBMHcH/hCRzXSjm2FXB
aGFjPzPfpxw0cMhh38kFpdKb3Lm1SZmnrzf530obgFzCJinDzdipLQ6MJDwpUy3VQGqkhKpfdVA6
sJFJBkHmhNRnOcVwNmyuAwDzixf/S95SK8CdU9hRBqJeZc7YfeqfxJZqkkA4sF1ywgWyCXbiL/2t
VlyatdMSkk7P+wi0TKZOzOuZXIzNJo72+11oGU0pGdWpSI5g1kpGs9ZjffTr4C22vF2Jscci85OE
MXNKZGlwRFCELkhFOdjPH4ndV/M3mmAqS0hTHsNrY1tA4QvxqJs7B+nXKGRH1db4RDas9WuYLBGA
1JGjXQpSvFRXjkyFEUNJY1n2JUKinqJErmPVeqjIa8bvNWJu/VvU3vWUePuC3g8DDOwEfQeyt3Z3
GWTafDmd9EpGwuM5u6haffyovxDA1Iz698rKCmezDE3EivD9XjMCxyXrXNfXnGEpTRzws09aaVKE
MUhMmkGQGxm4oQkAzLEnwuo33JibnMgOAOhdTGXqdoX3HXrYSiCQyds5hzwa+AvLMZRuY2IkdWff
POG0leh1aRfOvkTHWSM3hC62enerxyeSg6iRFJ2KFVeUgZUIOboWQCHVM3BznRBWoNL97XM8glo7
yVW6hdJZfJIF8Ve31BGkDZi2PUNuzfyykPpceYQXgvtGJKSp7RDXM2e7niI8DKZPE3qWpRuvcb15
9Ulpux7K88EciLWvazCsfTIh6F47KFF+v599e4MIl+NwolcqtBDjN/knr5HxP7reJOXch66tnJ+x
/JmpB6I+a3Eo6pL7UwmQ7s0PwZMqTtKAbjPytGW0tsY6ZMq/aIDyGkag00iDRPPunuQ1t9OtI+T+
JeidY9k2tCBADWHO5r53GIbfG/cS7LKKk3dc1gAw3HP/Wq8lsJhkLQHkIIml2WieQkm2+Dm9kGal
qZvZJTZtom6Jz7hPi4Y0vOC4LJ6aMuVnm59T1A/Fu4eBLQKDrJ2oOC+Nexu4mPIdAT5OLhVj+qOq
qQwuNnSbwfRfBUtvz4ZtNM6JdnCEoKabRdXgglYdmZvS/ZutfRo4xzBKa5Uq0t01G2gexzYeDQFF
sCEyLjGqvOKcgVPTCVWuLId1JNhuGU08e0VWG0fM1oxVEcBT7abbjVJqk5e+enOKsqvyfuf+iZ3h
aXv+5uaQ/fPBX79W5AfMjA5jGqT79UUQBBvUnOJzvk2HF/fZOvjGdTm4iRxN+/KcSF1asffKMoCY
P2f0oEb1bt6KeXBo7WMTyX8ngYL07Cl4DA+GDRCMG684UsjVoZkQfFDwC2L1nreG98Gm75R6jj4B
u2p68VeJS1tj0kVC5nnthoLD3VAZpM5b48sRfWPNLrgrgYAFtnijCZ0awi8KNZKoWHLwelSgw06F
NbKok8BOYrS5pv1WxJjnC80r5CfEMpX4Ho3hjeKWZYCzeWlcuUQ/XnjKABRKNUHmr/hYmKl2nTvt
9vybom6N+YE/BJ4VCqjAH2J8rPJ137uvqNkOCQvQgXlwVOhutSf5fNrQnsYfqYSpTIVZD0bCxwdP
liGS2fu7fWgtolibLnkFAv9QMgcjADLh1Tj9d6LakSkFNMYu9997ox5it+WG81YgtSua9O9A0gvG
M/YnEBu2X7sE1y6kR6VHiL8+ioFd1ckP4eHAGhSJ2pYENsQSRjqn0l9xn99Q8MNx/IAQGGTM0YDl
MWe9tGTWf8qyN1GBKRlqRkM57r/YbWaPeWcmT1bVekTybjFqxL/E8il6EEICX0jBRFEmcacu+FtH
SFVC/0Wu2ub9IC2WO3fWErP/Rs2AIhu9veVWaPLryoLZNtmnvDKZIV8Yyx16iiaiDlmIdaK8cb4H
rG31V061A6HqgK4kNV60BBzqmDo3bqxWsHkJMVmoDvnK2nX6pLw+TPChor85lmrU29wrj43OcEU+
77hNPz5otcwmbMAo2Wp2MidsveNtawlvIrteMbJsOOPfNPkq3DhH/wvwejwrSYzxIsHqId6N6Kdf
dxw0jvDP9fd1E/MrTyOASMS+UmQg/asphO50CYHY4NtE14jW3VbN/PT/xmE+QgAE5Gj28fwU/8hH
irrSPxS5WNKjry8J15BYz5JGc2tFGFM//CGz4dX1qqW2A90uN7e7hn2KMaGRsSd0RBkV3kIAsMnn
Al4mLNcUvmN9450M4DTtrswgVH9G6tY+QCduK4gpproBYnvm94Yte3F7AlgmY62HjAjuTCAb8Q5u
vYPoJdizIL4P1D8q1wEGhB/eoKI6Z8hF837gpB3e43jcpAMoAEFXi5x1rP7wcBLZ1batBHk1hJKd
a+PXxZ+5lb+51CbTKcRM2Iplagsdj5xKd81pE157yxCPZmtR08B2TFiT402zT7n6Iz7W9oavgdls
jBtS6h+JMXtRBQn8BsrvHjEKIaE/+6gL2tZcGd3LmP+9z0a+W0x4v58MKMYKcmpcIINxuHci2TeW
JiiF3OeQZJQhPsPBGztP/UDT4dwcHKcbjX+kl7oygPxVvOqEuvuMI//UQ1Z2/el/0w2SU3E/AQRZ
DRIx7AdTri8GMP9uTkcvVzKXwgnuu0R4TyHGoq21lDD8RI/LH21j3IfWPO0IYlbJ2T+C7Xzk5RRL
GlllZ0pi2WpPZxPX20bxUONiFA49JmToC7qruCTa57Vubh7Ch1osU0CH47IOOnw/fXKuJQh7yNC+
PcN2kpwoI+/iJ0NCZCJmU9fvMBjYHtQrGRgVLZdGUw6LUCxOVbc82JfoVseNfXexkXdeu5BDXIAK
CBtxTOF/O18JtYe2QSBS/88PUTOIHpfJ3pKC4t9NM028lmiGf9POSxtPlbiNoRrl2Th5YWvEm2gl
CmY4OMvtg29VB84K9NnQ6yxWnsVVKPmEcpluR1SimoAzkdDVWFQogthrZfHlao0DzxjsnsPYPxJx
ohxapNNs1OQ30yfuvN7HLJpRrnoeA4h4rjjlyIaPedrRgtxeO1BkK7lInZ0hHmUv3S/fCUvrYNwh
3PZJboCXptAdBtctU0tXBgKjgwbu0dHvZm3w6j3lOAZ66kkt/OkgZEp2G0WKxgH7uvRVx8Wp/Vhz
Tl9B0AzeeiXnW3VVGIzKaaRJO8ScoOKRD5PSHA2xC9XlcxJb7mJ1gv/Z5qmJYfbgG2FN80hIwhw+
86LovZT0zFU5Gr3/W0Vb4p/DCrsEMvi6Kv731nG8YUKByWfEtmG51TBOZheeWvp/8OznLndwH/UJ
wyFF+C8M2PNMiLLDh3yB3IFcQrp5CBZv5DpezeTEi6XV7bexSr4plnk970kJU4cyKQk8UHLBnvEN
TNRMlg7B9O+ykrU95cV4DMzRvE/v2GKNI86epV2mXKgOIXOMonHsYifh/NgaXc3Dl5mMmuDX6Ruo
nVARqASJDSK3LE18sk0cQKkmxlM4NIlnn2sV0wiZuKmmhtotbfYLglZ4JkEkswNKdZYfyHuWCyUN
s/R3Ddb9gHDld6uO6nfCBVYCGDtGBu06I9qTsIO+lj1y9kDUJc7jzUzYs5i4WFwMi5G8QBQsyf9h
TPF4HREnrh2GW+bhd/4HLnYbf0c+XMMt2Exh529+bhyx6DT0hxVQpXwLb57UKWnEG6wU4NXid3DM
HDLFVyEagog6Ew/CM1jNWgPBEdHNlXVUMbSmhFLapIDhu1MAXWaH0SM/KA8/kEOwthI/izG/XNnl
wb04cVhbw7FgsKcnEiSJeZOPFeXuMY4Tt3zLHBCiy6tigpEPvZM+9svbrRt5UiquPCrB1oN74Z+K
IqYv8LRJXQFu1y6E94TCJAYwcuob+p6djnDcdaWlDVEw0nmZl0U4930YG5cBJyF/5o6RS7mNNAFR
bJrtVY99acXh1Abk4VwcGBgF4Kp1WY0t/0Rof5uSUqRQuGZWL9DHAuhQV8NVRvWqHC8eXEr223Ng
vB+HBOYPqfeFrr1uUEAe8TKzq7/zf2oeJyJ9a/KgnN1GCkQHpINHbjzqMF6QZWTwOdY2pVbPOcZJ
ee0NPjfVAv7stgZ459ylOUuXcw87zZRXZB6OLd39ukUYekdEHRPTwxPQfVHFFWto58QAvo/wmRer
SL/XH5DVBnHMkLIHi1KMQog/p1bHTEM4XrOl8kQ+qV9ebgxtK71fzHvtCeYASZ2xQs6Qujda5SeL
gBputZTswOeeU9KDJfMBsQCYdzM2OepWiwo26AOsjUzIgnCSRe9HVL9OXLf8kQ2Zcz73XOBPOILU
ybMjdA4pHXEgUlk+ALjS/R4kLQu/w52qYdoI1gazrOcyibaBSWONRdwMm4azLzPIYgjctmoXM5gC
UWF4gMMTHAtO3weyBWXlHDeH80aAIa8ZI2FSwJ1fCXypXr9f/NtKzD/1cy30zuGHWIWM33KPmyR3
CS1UIDZo5BmEB1eAxFVS/ULWmOq8JaMRma0A/IbM0KhnYL2MKLmEAEKwXZSUEVYFJmZy/B78HD1H
QlWR9INjpBN2/CMtsVJ6Ui8bOt6sAw80sfg16X3eHwTMUnUxU3fhIuCKzUt/xip03Hb62LUGZnL7
0tw0IAU+fK/WMMeOi6KLURONl0086e77m4mcTmZrggV/a7sgZKuj8/dk2R+KnLxjAg/KRvN8kZRl
xB0tkY2hbhNM2/A7ApSaE/5V/U5OXXloX2tkg2q8A5uy9x4LxRNiTUl4uOh536gl/fuAJwTIy9rg
AWXlLhk16ymxe/CTwDE+wTjPICMRxFMAm8o1MqAObIUxvIZlIa2GWlWIMGWKuxJtFmfBSisGYbpP
IxsJN5+EbtDp1FpSfF7tTNC3jFLMKXTjBgWffPV/3V1mRefqt33vyLR563gv0cLtrqBoo6ZPxAzI
Vk+daPSqNJwIzKWj2wPJZ4XwDoJ5pz9UuV19OsKBtIYnnbkLlVEntwUw3bQnl5uR2l1G4n5tfuii
KPs8jfU5ALG13m1IObmh8xFeErjEsgh8N7W1QAJxyBNAYkonICTVS56FxCu0LNSkf0QXhYdgzBB2
OsZei/qtWgr0WnMfGiTlEZxmt+EBr+kV+R7kNw8EiJ/fsYU/oIMAY4PwVlx6nwNEoeooXDg/bTqs
+XOY9tr5Sarc6PI6gFUepmQs4ilVHLgwAHoGnVKWJ0A+k5lR0ikigqPPoQO1SkmqN+XIL2NVWZR0
OwzFE+k1/3AHdVqy7U+cPKlvKQu8WX470vNAM2n/+8zTdVVjMFf4ZiWYaj5+NDR8gha4PnHelmPp
fYVlTqFvYdbdJy22XgMx3ew2Oa3nb5vyP8+Bu+IcyzSkSY7aW3NpbEqW/1RcbP1Zsm0JMa44tWiU
Qa5TbWnd/ZarTVJZwdUuuQr94DxZ6IU9T3c342Llb7uTVOtOMSJuM7EvMtmNAdLGe+rTrptl/18i
RzQL01wKbOIdePBV0tinQfsExJJvffegUassf//NMLq66BfuL0dW9jXh1UiGfOh8C5APsMhiXA38
OA9l90c+2qNUayqK+SATHGy2opnw83CIKhfVx2aS266eFfeiOSI8mUhxDmr1luuEOYSVJmZIchW+
7LKIzJxElukA+EOdSHhQ2iklX00hMBwm8JNRuZdSyL0aJpzZtF7D7eiHXTWQn3sUCZIiFBBqLnnx
i0MGATL75TN06eFgl+HK0J/0/mHs/1DStvQdBYgp+9h10/Brlq8gNRQ1CcYWOeT8fLaUvcZGJFOC
4ljWYmhx2glgZ2yXAfoPH4UK5QBpqBJT9e98w2MLlx8yEt5jE4ZNDvMoJYsAYbv3ZvAKlTn/iVmu
8cnwoZ1p3N++5izHUCbNafcqiJQIHuRxrhWhGDM8vrIt+q/5aMs1HqcVlCdcWrn5z1eYFctkJlXb
MMkwc/v4RFwFntFsCflD2WesvzZcqko1HLEJ+msydsLjirk/OzcZqoNNY+VzlAlbktZWI+Hg+1Lf
GoH9pkihuMiaRp+6AI42l6h17hbEza7qLvVU0vbusk8m7kPw3xr6GOTv5k+k6Kom2gcv/WcpFn3J
ggSK/EzoOJQC4XIE4jSa1rH/TWcA/dOzE0gnHryT2MuRje8jTqUJNJ2B8pHHCAbUD1vvxWMn5LtZ
0tkL3sXtzEsLxVkQ2kz+bsmoFHIYMHaUKEiT3QnD2hoZdlLwL1FlMDH8mkjkvCr8CczbKwhWAify
Xctid7C6zx84VfRmnr3VAIF+GKakU2WhaDQOPh7gWOtDjsg5T3qNxQx6xm/fGcuH205IIyhz9SkA
WWYMWvZY9+kcmu7aQjcEOLDXGrvpqjRD31tK1XWk3F/IracpWFe+T6p+quWDD+mhQREH3a+UWggB
ulJmY2c7UCySY3f07a7NErTtOudeJHnJcA1QKFygT/CLnlimKMuZvt3+R5yDmE5G/MwzAgBwQjlb
jsbkcV+ZMFhcVOoyIrbs7+eTlggJa3RLUtCNg2ktleF5dtVTvE0Or8kl4qV26QrrPJ08/HxeolQH
7pDW1bKFl0UlC5dqaUoEMxIneP4du/+OdJ94CVWNqtyTNhhjKAE+YukrUMh30rtxZLbyotb6Ni2r
BCyr0R6T/Ay+7SXuViIuuLgu2m8ct6rUE6Pp6b3NqDOwmPShuHIaMk1y57YfCVgHExCUTZ8vPlXL
hFntXqW+lIEP4t+BaDEg7L7N6rMHLQFQtkmeA53VPJ40cq0JkqGLPAsMZzbmv+lNfA6n9SFBGmD6
bv5PyEBpIQmRal3X2I3KhmO7Ta/E/ifmZ6Px8OfRChmrSOII9F/V8VKYKP3v08d10rRWT/9mxmEp
oukZqMp0vLv/jZdVOKLBklYnVl4bniAncD6os3XV2NWgsuceM4970cJ2upB3Mm6/OAEy1ax9OmMF
VNuAFtk+Eb25y6qMivqCQvGHJvVvULwyQLZAT7WlAllNVdJnDJbYzoXv6R5JLpO9XYbl2gOpB7Ri
ap5ub78uQJmcWI5V7Idw8wRkwYN9ZR1MMfNqE24MxAt0/1tF7mzSk4sp7kHVeKmuR8uRWbnZMF/+
93Vg2EEzvHTs2Uxtlxt+zSX9qlIL9EqrjNwAgXxUpGTTyT99mQQRiZuIUsUDfMvjaZ+pfUzGfehZ
lWcpIwdslBw2B6xhol7EgCE5M3NEAthvVrfYAalSZSOi8ZrnYkQTYkTQqb4AKfoCcu9V/wjuEiyt
YK0KuUn6pKhLo4ctvqoyiqQR5xmde7l82wY1HumVTZsC8/6ftgBh2cWAwYdh+KyO1XQqb/ur/1gy
KitMJxxm0FncsReQYrQeSXiMXkK/39xbyzZHSq50Zmtp8Q4WCNFBjF5P20U/pW5Z/rx067304jKg
EMMLs9sPMuK+Etk8jGf37sA3b5MEwejdDfhvxDwbHjricoDtUlyp9ZVWozVIjRzPro7dtBPTDVg4
OB8/2jgC2HIgf6sZP+us2uFlGoMgtJr1lvUahPK4c+xDSHyCU9fDUIrSiafXPJ10/x8agwik6Mji
Z41oBqSd2vcHQXb7iePobFknDAArPTNCzlwcwIVbIX/1f4Y/7T0WDbV0f3tpZnys+ze22FJnXE7M
sBdfyKpKPZsF7BbeF94XsTQuMAiLvTb8ZWQboFpq3VP5hB6ljACWAg+JPd72TiPcLh/x6YIZpJ2P
eSzi2zxmLle4HFZfRPQMPTvA2g7nHdF7IE6u2cQ3fQJ/UaVF/KlKMqU80VzcTFfwq6/6RNgcKaW8
bndU8rD6h3PEeRtGPW3HTpxeLJ3dhI+FIw6wy91SYU1CY6UDA6AOfEKrqyXmxfJUy4v00GCfJe04
6tVQrIGZPSaHUTz/743QP9vTzJ9KqDC026a/neXJGTx3DmhSFCO8pxDhTXfwHP0KgO0GBjJJ3kJ5
JGTlhe9XEF1ynH/Stf8OBcaIAZnSvTSYFQ0p7KlqhuRK+esdwexj/QQwxvHYlzYdTvUMUgN3WF1a
J38QQXYMCfwp007xfeIIFgl//xHpXc/pg+1mNNV+dNkqPrYdHSMpMWFNtz6xJpMGHvc09m1cRKVO
8NbrfWqo24gctPq05gb3kwbauTPvHapA5+pzx301WJ0GcVONDG2xTZeVKaKK+ZZ5cvtKSBtkp9WH
nizyI5bjv4UQBy6HGes5RkoNJ419ew5WSEwHsY2KvZYrqSf0x/cVz0HKp9hG/GBaF500nTuD21WR
HXa1KhiuUoad159gw/R+gW3E2rA0s9w3mr6BttRehIAaRvjLlBaVfnuIJKezQeorDq+fzwspi/DQ
adwGCsVCdWaQit4bvYDCIZ97M1AY0HqSIIITUjBNPRG/rxWHLgmZDjVM9zZ7v4IC1cfdqL5Bmn4x
BJ3GGWBZf8ywlAVyByZ2bAw51EiictHYsTEW9cqo9XZAkzI7BVf9S89f9irLHLZksJRSAaIZJ7NH
zGQiG8F0N+vY95hyTQtLccc1q+AGAyjIkIeOKAzbFInr6SNZNUkOahW56bDiKz/3/wtYWQWa3R2Q
bbyCDHEJJClO+QsZ0reZmUPWjMYYDLzER53lBFdlVVDUKtt1E9+cVaLh7hn7B6NlmwtGt9GvymhQ
PxXGnLIcoj858T3Gc8K1FJc7fw8TM9IdhOZS2oFJQuGBsjzYxV1CHT7J9n7Apj6szGQr4o2KTN0j
gVV5Fwr/moQ1pIzQO+3rSSjKp+mRUkWAfKHOEyKllUx6SSa6in3VYzVOgidOXdzJlvofVJ3Xyeqv
w81QiP5k9/nKyw48zA/VYKkPH5ybONlvyPJHaWK4Bk+QqcuqOlGA/GzJiqssHTSGlzdBhjPHNvCK
ivXrVmFcr+SRwQhDkhrCFEzu2IrBPqym7kztAIcDdxLGBd5/mpqR8SoqKYFcAuHJPl4YaoZTKLm/
atTlVHZiEXTC1J9btAANNw0pOjtTcl0bQxk7/ztuXaqv8gKbrDxWOENdt1vXWE6tdW8x6RaKX/Xx
z3OZ/GGwqEzItd1cD9d1A8cB1fNUvaQ4aqDSlAWB6dnjxMoRSguK6P2Ezz4DbQJfTs5tQVHpg+ta
/Pymnr/APGQnlcIBL1e3ZnWArWzCtaTbBUNC8YBDdCcsygUK6WxzglIKgIucjyaIbd6Ejtw92jSu
BA1bLtDyEGahuqHYdPMDcD6dvFkPLdlriCOhodM59QnJoe19GozJAIYwZanSl/D3HpNd50NRYgb7
7n/SthJx+2ryfJySCd7VKB3aegg0WCp0ArzmYDj+6Q6TlCfRvA1YZOxihiNAORu8Csh6ExB/76Lq
PyTolY6C3Jpj4xak7BFqrqCemJ8zUubjwtgisYWosOYTwHqSIQ3yVlX+fG/dxfJZK4c4211SYzEH
328g+aP5/iFxyUJMSP4o4XKqe3/7uzrnhz5+/oAft1h8VkXXUxB+2HcGmurur6/A+lqIkAYGA/3k
CHWvcEAh/L4aBdWHTAhRZeZJ4gYXJuRgKYzsHON+Yic9qV6EF9/WQqFdQX5xhmK4UmsSYUK9b6IG
Og3raFpjdWxTLtROn9Tq8O47NUTeglGL3wHnmNVurCc3cDCqvp0W+80e3Pnauji7eeXfuJe5UZrW
uwdlKsUN2EQsIL6/iXWQuOkuezCVe1zsCvScrsax/kMzTGaP6SHe8+mQet4igMk3He0bScfpOhPm
D9W/lN/q5X3OjaYyJhgktZVIahQV4iMLpj6CE2XYxCAzhjg+sB7Val0nTm/ovNj2cYz3we0OU71E
g33br9IjQu9bDP05WDqv4p3CLeIuL9QIKkKhfWt0ur3w0ZQ1iCrGeSy2tTuFIy5G8ZQVwF72qkZ3
CL1ME9Q8yinqXYWLgRDwsxvOxQYuiii4yzFC9fiwopFNdV4B5nNlYPsb/koT83lB8CIlOexqYvcV
3WmwLfZ3oSfOpHGYh5zxD6ujwUs3BRqSCnaEmP27eHv0b8BDtc0U1HXtWCBAkHMf9dW1TbKJRIZG
iuQml7EsLn47X6LGNC1Lg3Z46mseyHGh5XGkMLPfZX5oYyKA2Gm1EFUMgJcsCDsMqm+TCukdMXwi
9anF1T1bgQak7XREBQgKS3Q2ISapHPZa96PAH8DtEGA/Nrozrfx9ZNIOUlHug6YhZQGIpd39j+D1
JG6S1vaKzFEh4l/LQXARyq5Z+C+uSb17OxAtwpuOlp6lLiQQMrJ6ftxaafEw7YhzWy5Y+MCkRSnH
9EqE8uTbj+Q7YKZw7G6v8qePcknbp2c5EA6LQxXAVWBd5KJ40+PNEXbmyxpSNpmH+qGr5c3RqzQy
J/URML2PW9ho6Vpa0ZaoMhpcFw8RVGAuYwMnoeu0MyAzeCmNJC2qKTlV/yKdJOkSZnhjJmruNc7j
43yMt86O53UQzbyHzR2StK0zzToSDAUNMiMbQ3rpACerJ/IdrFVfH22queVd769V5R+XtMCGxMDr
tzZW/Vd5zzd3UzmYkyTtCSwsjsQR6/aMNx91L7ChcR8HKWXdeKAWolqdL1q6uARtNyy2CXb2ujWQ
7x4Zk+M0J0kUycVnYffOGzLQrNg7gdYGGErrXtFcrSP2EzH8mwGTuFBWKSpip7lXJmyw7Mx4ouMI
TbIEJABsoehyFLZemA8mWtkxlQ021QgpTmn6cdE3jBL2Q92QyoRbvTWsRcCKmWc7p0305c1SQ7BD
9x+ahUwo4TgNhJjJMvovj6D9PrDh5YudijmVcnu5d/vD6jfay51yJwD0rqyrzI9+dOBiBJTpTxJy
c6onn7YVnfdUj3DgiGIuKdeTTbEWnqMPRQyce16BztBsCQYDQrRyg9fJy88nIum5c0p7iMBXwMQm
Lcaa4OlaCOHdViNPZ3ddv6oUNROCHJ7WBLYcIPmKd+Qw+8pa3BYtd56SAzihtN+hTJEwrjbCTTXZ
jIOaAcVRBpSz8kd97be56kauBCzgZ8VEXf1igKrIveQBQxP+x+CVjJSEWw1hxXgSjI+61qL5emCT
JccOYrhJLVtCL/mWYXjyQTCx7FxPm7VetDUZFhrytGpbmc5qC65kws7zfuj9RhmKE0JA0tqr3/XS
niUdxMPFndH4dqjm9cAqUh83mqGMFWn2jRl1KyE5ux5jFLEb/+ANrZotrNAagciHTlM6TCykE2+U
bcBoC9h06DSymLbqJL9KjUeUwKeoWJEMs+XBjH72sKGGgb0Z4t2Xjy0KwMDZD8ZdBNC7sC9RVyI4
2ONFPGVLthyWRngLupQ/RBZUqUcP0G5+pqZ/67mToyA8HK7TqW0zhOCdwoTpuV8w6iSQ1x21IhKI
mk76G/H+qS82YhGy5a0IjvSQZQGE/BCdB4C0FOeFS6iak4KuK9+5QP6fm995uAHqubf2Gl18Qma5
3I8uPFBSLP8ErtXfdlr8kU0IzLj6KABx/whEW99M1vdeDde1B9j1A0ppY+1pYlAugHsgf/tCEbif
I2am9A6g62WrUbFyBXZ63xOJLRsNf+a2KgfXFV+oyw3eUDT6OWJYRmoG/uYzFU2g0klS8uNlxq3S
FewCypKUN936St0ZqOQxqHMjfjFv+xI87HrCnXcwOw1zsMb4PrV+bNGNJIaCAIoZsrOgEBewBreO
uv0e7Jy3F71minNVuulZ0OBp8EuFYf2v2DrGMxvByzg3pYmz1yDWy6Nxg/MWlyWCWPYp1YjcMCWN
aBz8wtOscIzB4OjfClONF4L1xGxOBM4adONY3/iyenAZxSjzvYg1UON3XP+s6oTaAl2K7tNwmK1P
otwPFoQDXNsZ8BVnx7dyfTSWrMppKlwkHJ2gPFUTssptFSFgE8CPH4R+9NvWPu145kd/lDT9XG+I
GXkL07hdaZhhT7jai17FMZN5ygNnLO3TwIGJc/KfDIdl6uIuvKtgNmae1SaPN4L0P4x5LqZVxhfc
eyZavNL7pPODs2pKAV6wgTdpgy+rsHIByy8QWEY2XnQr67MTAI07BtsPQ1XSkpfT8iOe5+xzL/Zm
eqRzhoH1uPAUQlXIcxDmkhWP1vLfgJ4gJr1cgRPowCgIQVhgkGqSUq6UZATg11CCPsXTyXVW2Zcf
mjZK/JKBVz54sTzKsQPOCIzzOlNavRY+xfLuf7hVhW9lD4krrsdE4Svhj48SGIzSAExydvmN9irW
rogr90GwCFKSMnXNbcqvJ7IdkEPy5Z23jaidyA70nUWQeOUU3P7wVlUJXegGFYrw4j6fQn4CEC+8
zDFTzUWSaT+jEDcZpHnVbRyoAgQ0WswXXY+dV+7DgyPax4EkT+JHaDDS9gZFNSBFTGsDc/KQ9KsD
XZ40JQ8pUOGjgQbk7ly0yVxXCoBnE8vI0z3CbhyZajX5MIPlOJnr9Uigtt/cgNMW0pYJnVDMioEq
NRnPgk4b6gKq20n4cQNXt4g9RomG/hnKUnsSwWCzOf7KZBmr7EoedPmTLDJlcG5fuG26YSW1OJlp
PgKtBK4tWNVeNoxQuQrN0Jt0P23MELducZ6zPMAHY+kxkRTWwccFW8mdKiIF0lOPSoxLyk8Id3fV
Q+O2k1U4P15XsPUe8JWmIlWmjdrZj/1XkRlhmlri6Um7tiknOKvWfe7zgo1k4KAVzlNMvPjWhySK
ZsjXTdjXEBCeSMu7NHk2e+rh9o27GgZNpJynaMZ+U5UJfuEctaK9FBjpwDL8G1EWVXdW4IcoA2pW
cCiFHWuL86Fdxw1qVfotBIwd4IhAh31w915SjSnEFkrNltrtxVD7w4sxpIQxu4lMVt2xKF5ArRbQ
7R0+orYTkB/a+HIZ/q2SkHDQcF14x+oQUlbKWr4hOJxGlkP17TM0Ns1djW1imUgwJDxv4+705NxA
9lZBGDYCByiScFp83XVn+TnI3Sx9wTZtwcBu+u8hZX8haf51XfdIB/PVTb9i0EDgyuUVwv86QzY0
gY7XeskVuPiS4OY/fZLBOXMkMIejB18Mr8iEeMWNQc0akLfzQItQN8N7HS79mLlw4jdHXrC255hV
ACTV5MLxFbKARgGtN+1thFVTQUHpcO37lh1TzLdqsifyCmEXj8STbvxOxsQ6mmjICfMwJkbG4ufc
PtysCA/QdpPM+JXw63X2ulbiuvReVsKJrz2MSLtcrIe7d0+5tms4SoGjCSs2ihzLiScVD/nWjU6U
6ZWUhnkAsRjk63+1Zsyl0p5BqLg/qYxPoSeu/iG4o/6tUtTVF/mZgkjE1UBbD/+5jJTvsNQKLOib
Cu0Mwzakbm/Vo0k3RV6/QfUKoTtDQZl74jGgBsu8bPkqqakCAfxJ5t0/iTq+Hl5q+XdUeRmqYTBj
nXMXetowYcZsmsasfWfPXAnjS7hnsfuxftywi+3RbayBrIdRh8plbEfVZoMCNWFNJ2zSYOJ+K4nv
cOyN3p8vBBniKAg98xLaiSa2cUuJo9G7+3HkzRSbgvUm9SN7lZUXgQPBeonl7YeGCsYRHrz3kvAO
JbFMLrkzNxo/WnnvF1p3JPJE9KgfGnqCVLlLyybar/IBl8XmXeZCxnCjS+RfDTga+FtS1AWrmM4+
l+enM0i+JRzbgyEoc07U2vlOPQ6UC7Y4lwqZtposAAm4hu9gGLtNlujZy1ZfRn8CycARUOHZoWKU
bTG6Gtkwx0a8WxsfACKBxEea9Vh3/0grg3LPiGEejEWeRpiutJcYt2F9SB9X0Be1Mp6IqKQzyr1w
wSCbazPbdLoiiP1KeTCB9mCkA7hzfY6q8EUQAPnXM9Q6jxLysQ1OvJHI3U+M1YZ5U0Hww/Yds2Xk
CSi8SYDWWyR2nqb9VIIaI8rh3KKKtOFIlJafUMzEIa+Vt8Fv2ssFHTSeV3gG9ANjLBc6Eo8WkSNE
GARWghSyrrHbYeVGrELeXSFe5K43wB+R/RzzbvmwLWosDEJ3QXwSu3Zg1NBvXXBuGAuE0WiXNkp3
zGLCIplqD9lH6F5Fnd/yri+u4+tuH+Ze2jc7btR+GBWkTZnIW4ZxeK4Ja3rzsK6nNU/ZwYVg5FCO
GzW9vv2iXlQiv1hKSq50Qx6fsFrTm7j3GQMdpQVXmuUmFpy//Sej5EEYgEy26Lm2X7aISLrzhLeq
QdoCIe1WzfXkD16cr8FFCxP/02kBz6hts9hcnX6/9CNZg1TXxWCJF7CTz4GqkW4+3Y5qvNnpGjo5
4pqP41ettAsVUYVE8SY4a+C7H7GTRFtz00KSdkb2qvHWIN/Zn7T/LrT8x8SMNLLlINRMgJ0OtlWd
jIhJSnL4opFd87AtsPxPatg93ZLlGIoekEPJFdovZXHKKISZbV/Jx9PTC12m04/0e1kpGLR216Jm
D2lkgrXUl1rdOop9M8it0FiiTPiQE5iQYV5qtRnoxXA72sv0AbiLsPf23mzSaZk8H4mipvu8b+6U
+Kg7KX0LhRb5Grl67t0z7ItkXTB0429hRydTMFOt3OM+KkID9sikIBpUDXZ1psmqzbiYGm7vpCj2
n9nWGWyWAtpnFE7Qouf4/grgfQimsG8Q9wHKR+2cV8KhzzTt4qx2+vj8KZIfjMh393hWt0pw8AP5
fCMvrSjZNPf9J9LN3G25nPIid7uWdXsmwDc3Ci2IEdW9dxvKQ48q0YWOLPxpJKEZ0LJMxZ76mVqm
+pWzPV+qRnAVSe2ncTIZX2US4RJBlIjehUxDShU4iC/QyTJrKCe+jnmnDQsJ5cb2JWBlotkDQum+
IyQL8I+CD+9/s4gCEt422GnLCHVAdGIcRSG6DyW7MRzyMbvbJCpCCJWYGNLl3xYddXQ1AabSf+61
92A16XOlQqk8rTDHGGJGBpH4j6p9LX9SWYyMbrQq/BKiFKTsfDusFL7KJD7rLHuDZ3dy201ouND8
8nnI7u6cv0XemzridbhMABIrpwrqY+UDTOa+cDhhcvr3Q3J/DNe7PSAkwI7VkHxnjqRnld1Dnp8w
NW3W56DcQaq0HQr7ksRpCXYDbF/s74dN1SgRM2lJeWv0TcL8eIx+/E6Ev/QC0waSc5Uopz+5pAgd
urXSu1vhUD0MnfwG5QU+MuUwgcpF22c3Eqap2xaCxk4Ol0Rx5n6BygzpiAs1IQz4+2Hl/r61g7or
VR0gfx8yW3yXRg0dL7eZDSU//E1n41bmdP1Z4FzLKxXPE6d+JfkHc6pCwPEXCJugaDm5fNptBGRR
It41fKMPetv7moekK2KxZhFTyXkCJCdWZLRtKCjW3dKwihehn8dj7dTUWHx4oPckJTojqgE6syms
ACan78Pw21bXrNOgyVtEKxCOHrNQ6QLzWvRQiZinLySeIvTsYIGmBdiGyguIr1zGAo+ZK6uz7gBG
xxnnnKV1HgNtJ4qbiM7ZA1nLV0nKqBlEGzcAMusyY2AnDz6NUT2NiuoMfBYMKfMTDZqEKDAEx04n
sdGQQMtn9wPIy0pftLKLUQpfZ0EbYdmX3tbknExC5JoS2nqUHqoOamfjfRfzHW19lLLo8ZT1BWVH
AWBAbesPjX7Dq681AKbvqD6u/aeA1CRRLa9RpvudWNsQJ+T1GSlgnBKyYmjf+QQ1t+CCGD9qOLwU
g15Vfn01eYMzqyYpcOUpQwD+Bb2kjtXLAtkJWKlS5NvTagyS7y+RI5PtWLO25cU7jVuJJ7kfTk69
u8Sa6WxgQbHT+s5nw/YIkz1GWynrg8sMzweUXq4lAt4aTNEXvugDVo7kB/q7nbI/iw+ydXIpYtnV
xJvc1pINtx4uXQQmCkqUC0QG6bMea5yCotG9zA0thWfB8BL9tVuO6mOv2szvcAFGUHGLILYk9SFk
kb9HPE/fvbYSStmOH1BcrSwu7gdPD2vWSRjXr/bkcUxklLjV0y8ZW9P+eZ+kMxLgRlvvH4nBFaUA
1+T7D/dAth07SU/JbrUbG7eMdj2CwTa4tM7uqWlLPJjJu+mEQsRYxiGLXTTJl2YD6tZYj3gehhWP
4ETijYpqCVhfPOMUpdPYaZC3G6iCnDtsLvUV4dDoQegeeZruePtuvdOKWJWuyyjsysZ4l+ywWA3g
GgWNbme5ahXXgIX83SdcVoPnUZnIZxSmLG4AV78lXrY09j2quWlNnidBTb2IUi2cplRPEPy1WifK
Zp9jJpugII56axaT5Awkeeui9dbZCxZy9dXN4iqJfCYo/sMqA4l1sE4xm9Ou71xvjyNqu6II+6uD
VukoFupptRthGZNoc/dp26xJ/3UVoM+hsae3RkxRnD5PSRS5uuNdgfQTBqY4ScuHhUgkCbNX3XxB
G3YrrEW4Z8GU3/JP0j2RytaF1+08qoR64GZxc1zZOiijPhCnCrUEqIJYXAa3qc5PzuoXULfKWPD7
+ZcQ4b9j+xb+JEc0Fzip3WG0brO/xwKvJh1m1+ItCSMYfd3SdCpOlHTcE1DiUQawD3v6htpvkgXW
SgY8ZJusgRE3/LRgE5l1ncT5i/f5zPE4eaijHsgmkuLvMxpJ+efe91vLiYKSDH3YA3H3bR8Oas9V
J//Di9HmnSjzJ7pYVeOcVYiYCQG09l0pcrDCVFTXtdhAHA1kjo9z5Q5LzmRgFS9I95fiM/gHkjFQ
xCkO3Y1+RTgAO2JlN2vBsvdOB8jdaLAMz8lYDR+k5m5Wm4cxEasx1DMhEM0RNVnM2oZKUb8bgJCX
D0ejxGkZhza2Px9cCpNQHs/l54sY9qtwqz/03K72ZvbD/mQGhG1kRo5Bchi/+gY8lplfqHCwyUDA
AgV9hT25e8y/yH6dsQs8sNEna93mIOeArDE9d1Uvtw9Hx6rO17sSQbUlVCWLTyd63IbbSNseanny
xqP6M2IahC8VmEvC2l5Mh8cwuTngfqwRzbNij+TCB4r+H0v8dQqlS8dSmNRGBh4sk4wZqSCkKznu
KlrIUtQQQe6cJo+goGwAHbLdlwyOOoEyk+z4gio6I7mu5boiIwx3TeeAl4wRI5vfUprCGPesyiiE
rJ1j3DilOmC7+TCcbZ5vq0g2N+bGHSXgUzXKTR6FhilEZ4YwCS8yz/H2rzn54NoqjGmIvjZv7TOg
p5Z+MLut0HFkJjStz953DgBY2VQODqTzZIur3iA17DB0kRr3ANgbqF15k6iAaKVxYj4ZxE3OmUu7
ixKB08kgp1gJOeYmz7IUhAS7M0G9JrHE2eAaMUWWroHwEuo2w7xsDU1NYOVhiCzUCiN5IPFXxF1E
RsuMwrIsBuAVn3vXfxtkfOoN2cnnOZ9rUzad4XRu6qJ4FtlDJNv8MzqDoz6tDHA0yueSBFHb6CpT
ifsItdR+O0OP1Y0IWMyZQwXA9KIsd/9rbmXjHQdto3w6Ei3eX3puEgkXYibNsGuCsCYbFSICOS9y
FmwbKDlSoz6L2QnIqEs9z8CYGKs5N75jgYRODokBZJJ5FZlieOIGuKUqYSDlQ+1EyV4cte6tem7h
LuiJNDkSanhNJhqsI3vMhxzqQ/Xq6Yoyujp9uk6fTawkp/6ACvEhaDcS+943h7igqRf06Nw5GU2V
EyoE9USLP4k2uQeS+llerYAYQQsydWc393BW/wQcW0nLbEaxpn4ds6C4n31iH1J5cpKY4EnMsR9K
mi6m2DZ5a2WGQIIuBDKT51OTFPPUkmsddMwuc1NUUUBkMkzxEAQ3CPrDNMSK77PT8ZDaBaEWI7ue
JOSQLOhdHkbg8zi7g9YScGboNjyXDsUyH7Npf+faUradK4zA/rySz3f4XBBAWYzuZ7cTWzElH9TD
v6oxJzbZ19LxKunX9rJQdpH5jfXX4P2Aqln2XrrP2jYaiDdfDsbSgCMLX9WOSTkmvmNMOiwBhWC6
OEORtWE3hwNH9hfoS84iz1RANkDWrxQs0mCT2mj5YQydoxVgDBSivMay3ooS941qc8e0z/cAh7/J
BC4chkWRvnxbYwbdHaFl0eXgeH1sFPtM0XSyabX6hx3culeUOp1PX0WcNsBHpJU0c94mIs9V9UXN
p17E+ApIpmbHGTibFbL7zHJ4ccmc6yns1l6o/7m/NCyAHpa/c85kYNNP0/ygQx6KAeGQpmVsp1nj
NIbmTXsPCoq37oQniPJ9MDzDpDEAkIwlawGM/yneK3ejIfo7Lr3XZDxphiMn1QVTHhkhWdMO1hkY
lJ+Pevact11yo2brGZSrrS+TIspved0JGxA/E9Aat8t9S6x8t89Ir93w83FXbkdRMspwmB8cWBE8
WMoFqnDA8y4//bdRfiSRlz7YzKhFmwYZBn23KiAlM27JlCPWDmg0SGu/13fGYHKSbrCTOnHb5Lou
WRUM/6FTa/gRSYBmWCRHu/gGBgC0FYs+96BKDJLGPBaR1awSLvFNGkCOMTt7tP/S/tz+PKvoLVOe
UFyjGIuFrG19M2PJVC3sQ/pBBDaSO3U1UuYmhEAcq/GONz7kYT8VVBCNvsCjQQkXvL9YQyv9amUH
qJX5FrgvpAjqSVTrcj6T8sbhKijc10ZT4qCjRARqwskdGvcPpWnFcCxAYAayCymtay+aCFCBYy8e
FyfY+fIoEClGjmmj7rx2kRiTrxfHCvojbpS5e85Q40r7AO9mtTGT8Seeu11QekyCXcasD/638ZC7
0zdXQLPVmQXl1eiWA5QAAgGAVBOduyA0s1E91MKXVjPZjPnByqaJO3q8ejGrqdYG/r06qDk0ikJv
dNpZZecEN50HRxaB3NdicCILgjLJkyYYqEfg55qyMYZVbatMpiBckPpHy+d9GVuwBlepCEauHRWk
GsxS5ad1Kywt9Morq7hC5hNGUEQF0hxkoIfYmkrw15ZHoIboiSO4ZFCY9JMqfjN8N+p9+LG+N/Oq
YB6D/EHtTDy7PE2JnCxrZujXFCaQmBTtubimQ+edgl0mzwuJXOWpur6khOE/RzTISpEuvgzTCilE
bNLcVBgvH1S1AgywV90o/aQqdXKyoT2TlxHiVDmR3mdVR4b1ebd9iCMJKVEpbkOZvIbivQ6A/JWy
Bzn26MuteF9ZoY9QuW9Z0Aiy03qZFjsXFPAzT58WLEiSFM0hhtx55wZPTygglrKkzqfJYVdN2vCA
E0N/kvxYI/RDHbcMY3lCNVJrr88omvpag9ma6ixvNwad8jmJD5OLvithHXpkQliAapHSJdOUgg6u
v9siXj3X3lKyZ+Ql/ctcu/PeQpJZDqKDQXyXh4YHqmvgoy2wGs26MJwFD3ckcbHpyNh9sZDDVt6y
LS/q3uz4rkEDx05ZMZW+aTwjJO7J4Ip+SyIpY4YK9EIBGOdRipz1ev2Eq45m+psZEklojTbrDWpx
nrYCXVaDktkFu19Fw1p7Er3Gss1C876ngQEz99mMGQPkpI6e/5yjhrZu/xjBH49RF0l19AKXbg/U
t8ANL4W3Kdz1aWzKF4a4WrCBwjvzDhhpTeXBG3LlozwTpnauGVH9r/hU5WhZsEo9fEJu7az4MCTy
HKMi35SY6GSfkS0eOnKCCKmqmoMDc+GBSmsN/6h+9OGsyT3xBnljxvS9g3A4KSlaJrUOKWSnHIvR
yL7LBNnq8E8B/F8UVjhMTO7+df8HHK4tIE8lAqq9o9u7SEMZwgWwmOC9kkhjVzxlY4Yd1P+YWUVh
OuMCzmhQVItr2WrDzPWfNsFSdZHl+cEKJ+/2QnnZahd7wuvCU65RKtBEekumjT68dUjabV6udTSP
doc3GQiH4uIewoopzWzw3B8kyKcP+4hNVGQPfPCGd4TScKLUbwz0rmO/lotzSQijVE2ZrhI4n5NC
Bf1LzHYMBRemPVqmBQ69WLexGg/6mWXvzAklwQgR8Vu5YZZnInOza+ig/cCfFTd+Uxa5uVRs5CKn
RsYMNI5lQATxZIoa0W+eIZt3pPYqeERM8emG9Il4H5ceGRmFOgEhca1wVOr1tqS31Q5YXJa35mxU
LpExhg/I1XD0xHHkoC0v9uVJv4ILO88+kgLMjNBVzmzOQ7KsnRrY0FhMUz3A6SwDaMFJY3y72MGt
dcXbBa/VxrY8bbAvfq51X3++qSCPWyd7HgAxMFZtankAuS0OxSNBuzugw+VwAiX5480+gvFOSGNr
7MSnIxJxcnKsDZnFGQ6lnLUuCspHNKPcSSr0wq/IFDQQn1cFJgaaNBmK5GrRulX7lMuFCPy/euPG
WbTq/5PRd2RCP23mo3V5is8wNjwIH3jWYM42mCd9A4oWUS6K4+yYy4RD/TREh5J6W7DECR8fHXqn
dRkAKMTB3wAODRMWVaHMLnZJXjMKwiMULlwfu8q1TxRmZUHtJLaCfRMNYFF8xLhwEBKr3cOrlumy
gBNnPlc2sAs0AdbnSJoGS8392jLA8YGVc6XS0PEJGwUjvSorHmX26oymr1gqy6FzwcQA72xw8zlG
ZJk6hj08+s+briTzCnGLVR8p5V8F6pZ8Tcjana2oZ6xjZBDJYQaTM+T4cTjmLWc2Qd8hSCRPQALf
Envi6kW7fWfdBymdJo1p7hSQCvHbhc00nv9b0iIf8yTYus4qM7E1lAYPW0W3ZUoqu7mEcfr3MR1/
9mUtJC4L5ei63zf/l85F2FguX0MxcZmTRgRWc/58sh19ZuNd7xN7tkuBhNUkSbiPVusB3DWxjjvu
4xRJIEqcGp+HH8sb1CFkKQi5ML3y9Yv+aD36gvqO+pGxX2aa5bBjR7PCyY9gMc46BHk7TJVBeK5j
NLnVmP1Q7r5iA55Jzltm+S6gYcExg/tTl/yVfJxRTp/EoREa1ftYCDYHmZvax5p/mCdOV3my5tJr
EWNcVBXbBAKfTuqsP5t4m5LVozzsTTrJKXcrwR1O0i5etfPUxHIGgtp84t1AoFpFzJuUmnnsCe5p
0C2t+aDzfuBjPnO3RfJ5OpwAT/K/NSUZIEh846yPuj/HGLBZbTs0C4PrH69c6kpDr9+Vb+GqOEE8
zWBexWzN+sra+ouqhcfAlHJJOg8dYGW2BwY59UUpeFt0xIVxKJsXY6aIP6I2ynVN9iOj0P+tJCcX
N+CB7ypgc0sdJTsOjPfUPumGq8MI4a438gcE8J9mnTpAd5EJCVm/CybrpciCKmcZITV0/18T6sSS
z4mOFSLWGjvoOsG3EOxPLxKl/HVGtfjRMMaTdiF4uo2iGx+a7HuvyPwPoZu/JH5U7r34xfsDFH0L
+KuNjeMGBEEuRfTN4uTkd89TU142Wng6NDFOR/f9PM1J+RgBWPh7XP/qfdHaLo0AZG4/CNAI92sz
ImG8fJF0/dVNoLbsspQ0fZuxbRKJVYio/6zj7wFoTqNqBpevMFw5znz6sjNdxkFNqZnPB/ok04AE
loVlVc6bDzCXeVxUuVZOr6IqeEqAAH6MqGJAC1+ksYh/I0+AHM6mzS6lBYt4w7VMNQphsoOLL3ys
iqtoWN1yuWaqg4/2diSNOXWrGsQ56MTfI+/EH38YovLwl5pdARu0LUA2c51fVKVXkYjFmVRo6NWy
myIKAj1ph8+6j1akV155gIoJmGmY4GTATq+Ntv+0OL5jwoUsBbDFx+bwM6ouGXdpTEO/001QeZac
LeoIb4i86fqFfZiJprqK5lHOjo583IgDPjqZF7Ch06Smzppu3PRpzOMiCrgN/JXtxjnEFQVRDczC
BuEx0QAdK0tRBgr9FRqzelZpK3Ps5rkNcKtyi5s570uRdK1VcL2uZVCLUTRxRuQEsR7S3dKSUXdN
qgsxGZMij2asRn4LhkgkUBkbwSqwJUcrDlgApfnk52BYLOji6mQImP1cfKnihmm+YXHg2xgmfgXp
4e9dzCRHc+/CMSVdSMiOaZ/vdFpD/NpaExVuEktYplL7DXBG836GCYAGx1FjSbkWunoE4a0hJ/pQ
JwIT6AEDbHitgY++ATAuVvwwgz7NKulwUtFuTFfhyi3Pzi4lNv0EtnWGoaEgp3Tx1jDa1Abgk6II
oBuFql3OFQLlZVBIAHGeKzV9zeI4Lrp75Jfw1ifHg5ZYBiSIdQPE3nN1p+tfoYRdJrDHgqjgP+Tm
W8Ho9dUtIFRrPK2hGwZULR6OFklIl54LtrRpPWwTUd9YcOYDi/c0UDaTiGlAoPTcNQ60lq09dtyk
m3wOHg51sZXkEHqcvIHdO+vI9SIFFe+4usHMTJ4j2oUm6sf+aHSPZdMk17UpEaDGlm6jWsNQpdSb
oiZjaswxs+PVZ1sbezV1gXC3xFWzSsLfIsbzx5/SQDRu7XURWh0MTlkhBVXtVoQYuI3PIUPpf/HU
bM5qjZ7oFP1MVI1kTfzcwO+dMU7q8ZRSDkaE5xwS5t1JO4eT0Iz+J+i49rC9/BUsUfCYdFtvPE85
kBoxfMT+LqroORi0DVCVPOoae5nuitos6F76HuTrVfif1YNjuGqJMjVkXdS8Z7dumsymzbPDouxW
/Y7OUA4pvIgoQpn4djW1aUyeBx8G+SaD4IZ1EBj9xy3WXYh0nbeTkXnU0uCvfqwE1t0MVbrgknEG
deZGKWqTuMyIPhmK/mwuDHXcgKxp203qOssjUWbA0+V7sdK9GtE1QIhtqmGzNTN8FGlyVR7qIMuZ
Mvqshb4YpyhX4zUmJUvAAaMei1lNr5r37RfFWzNCFXqSAMIYDR/oLIae4o0UKY/ZVGknCp/YoIJk
NUokBvnl0+zCenNpBoYLEr9oHQRkL2u9rfnCKwI3paIbCjXjsOC3I4PePSnSIp/cf1tfwzUmGQKn
VxVyHQ3TEL9jqEX0QPvD9IVg7hEa/04I/pOXO/Q3uFVSWZMlxkgUTopa7DsQPXsAp9bXoyITf6It
S0t7HkTW2BbB0bwAoJfLWO07ZawKmwWsfi00zWJX48fMzbV1ol286yOsRsh7+jz/p0LOmcwxfgYb
QSc1RxKBUmP15hkSNldArj4AIYcD05KKtQnAwGd8xy3+zE/SPVNlCPM9BEW6W2+zp9OLm0Sj94vb
FEpYKyQtjxw/61scdFpNn/evFN5j9TiRB5UAO39+JoZ8x9dzWTRGshks2DMbS5/B1wQdghO+Vd7Z
dRP4aFyvNy/0e8Bg7GHSBZzJI4ZRlueUH47A/5Y2eiIHYfnVVpuE+r5puhHTIoMv7mN2VFYTq8L2
/4QH+oYqlWpb1Jl2JEDc+zVIU/lskj56XxzHZEzSFHTItOT4IIxC+1YPKX7A1zFWbJc4728SQN0W
wd0x6zqoTDyuYetecXXymykynV02f+D+FBPX4lUGxlYOkrCBVi46pzKB3q4kbKTCxBJCx53cH8Cn
BR+jV+CrF/ov9Y8wQ+ApKaBIToOQQRU2suUmqP4D02w4lkDYK5Z+mssvYC80OdYVDjvImhaHz8U2
9A3eT3bO4xk+OnbYFZnJu6eAkczTpo3Vq7/rK5TPVfTbPcaLG4YrsYVvvWqMcwH0WUKv7azdP+ZW
DR0vVjU0yk39QxcmrnM/lG6qr9lpULLaCC2Snh6yUO/MfMSYSttrEBnAEzWWyc3gyilXAZBfVLnL
elNBnLjZamb4W5uWn8gvohYGIw/sd9CCczJuu2ru62OZ9P9WLWhHVyJCoYObv/5Qsv0mOGrhFbrH
ynzP1BgUcZuklI14pJ4RZSQkayzFUZczWxf9x8J0jNfNJUFAujorMCtQpeqgMgDiA9yhtbbE87tI
4wLiLJ4eAyHVJgX3JgO3cGPUbMLA33xAkwmS4Ssly8ey5wcZBLyac2AbG2QlTV7215gFNHc6GmWM
5+WLcwQDNkfEc5RcB++YzcvLlgQvPrNsRz062RhHwRuZPcEZcZYhZnxilGktkAIXCAXTHEyNRimZ
ujqka+O3EA6eC4yCuLEI1baJU36Jng2PYS19vt2m9fUXlwo74Iia/kxQJaCkwNuPNneA1WxWNjsN
adxaRoQFfSr/l/WZSArOV6ZxWFe4uMrw4vGa0LBMucXoqouSXnDbtKgYdI5Oprzwsjj8KGM6201X
y+sZFVcVE2w+BfxIZrutQoTt7uY/FDDkyV6JXnLOPsi3iLYN7lE4d8JOPbsMC6bYDV47MD3bbKr7
qeh2Fv8uzdLjrlXHfff+XZGS5oPCGSoppnWscLR7Osk4h8QMw3ANiox9GNP5Wy9yy13sdg5Xql7J
uqMeVCWekJO3W9Soz3GOypS18qPZHJOiB0ISGP+6iXS7Gmug7KfQYt+aGCgQ3WxNyCDNh0W0KqLW
8XStb5/3VYkKSwcgqr2ha57LsTB4EJR7Vajx1hbE/CRyRxotpHtw8bwo8sSeHbyYwOBJkOWhz4ZL
l1+fZ1aUgj9rh8bDCU06VkSRUDFDaoq9xUK9aZyoohSfu1cxxvXHaATyj8X8DqEq1wjWxcgXA49h
M+Db+95ltJKbgM4QBk6Okx1e+zgolBSy1i/QyLfi+CKGTyM5e0pWAKLVQ5K5b1TfQWpffd++sexw
SneHAYQh4RTvu1IEith4WruNI/ft6iyw1o6iOYjPEa4oaP7VjUFWBhiA+MgAeKCxI1KfZ0EZ2Uf6
5soqK8SONrhE3H2ZZb8LzrglqnkXOOsEkGmKF+esucBuRQ0+YDx679IxMQ2UDbFR2G8iwQJluU7s
bwAbLe2dkGjcAyYDjsF0zCPHue5SacjUzlWfEHhgfPxedSFOYSJ5VdvqBYF+ZrUWgr4566mYvTer
WJPCW/WEcjwPk1lR8V7WUJWyLejBn0b5u9PqHiLO+57YG1y8lS8mIy+iYrYGjb7McyDmB4Ih9aDx
u+ZyAUMjJwe7hLGqgVFO6oWPVUDfZv+gg64SLsEY/PyLIPwb04wK7juwgx3oxaxXhJvO8+lUhW9a
H7JCfkAUrmOOJhTH/cR5oLcp/5xbyiipSmB+RblauNmhVpYkdecB9Lv+KAZYcmJ76Szrl2+g4I9e
3rXI76l/eA2hNNVmDfKXwt+clbsj52zTiqbGV6aY0NknuWrAO7SN8i3YD/Gt13aJmSHfeBQ3fvL1
xIXEfys+0fQLVIlDsG1JXeNgpOQ0Swsysy9xzkGL944/yG26KFuYbm8S0GDTWtoNBv7ObHvuitpY
1xGtHBdpFNsnAhGWiiB+hAzZsCK+mv6vLvGQgTHg3rvzq7y2Us6Vli/+nYtl6eQok1RP7YXiQOxU
Nj6/4y3eVfbE+Hp11dpbgguO/l20tF2gomzrDzzA5wQ5vHjHu8E6/3Nkje0zNepItp/pcrNi+gff
310KEnDtt0WePVXijbX3UErjk0p2oBt69p948P1E4KDMQQpfuzUBMjnFYQTCTsWPfROSYKNDihVD
f3PbsYv8lNgFLSgpDPw/tPffl86FGLXsZPncPB9cwmANeHywDlCT+MGKQ6WbuUrk7UEk+OZTaDgf
+SFMOLr5fpW6mMhkobdWoNr0qiWk/wUG2FqVNxeYaaGocGpB0Zbz2IEaU5knBdJaFSWjCd48tGd2
L0ZsueMi8H7j7XB1et3cOcfl0wrkxei1CXEiOHWNJKwe5LuXjjkP3PwsLQJS3INn88ZvCNBG8/Oh
ptSaFdYZx/SaiM1K/m0hhITjlAolQPmLv0E6u+arT9+3TRPlOmpmmvKIbxJLJH9IWrewT9wBBzQR
m8lHKsMfbTrd+WQfa0mrLWJ9SjgHYN3JHQ6NQIO7HdKYg3qOYqewoT0tCusMBCd3wqG0TobgMicX
sOEd7piWI7BB4PDchk1sr2hwt/vAo5om6fzoqFTwf6u99I+fb8uJsOPFQdv8Kgm1KmCV0X4aR/yb
9kC+WLOWm9xKXtWaO4OUoVxQDCQeio3LHaeUPg+rcrlRB8/Ip1v248qqJg0Ij+ZzNS0V4XwzUYOW
q0xXUCgqU4HWrPG7edmVfwbjQITne7JjJD5d2wSISukEJOKAvXg3SiNY6oCVdpsBCrXog7y+Fa5q
PcJsb4uA3b8YPeUDf4KE2KFgg551/XtJRg0ZTdLq8gBNmV8FuFuKiiEWZAAwETUiRh9oO28glM0v
0QFm4LFKPjhTr5WDp2X4r81naPJ1deQOEGuXY2xJWugb7SI/jgmmmhsQFAFEtBj8LDNTqAhvm9CF
lb+Rk1LhYv7Oe38v0KkNwyc+yTevS7q0mfA7LvNpWzuaMu+0IbTEdoFvv+ucHw4TyoxcD0+t9Vmx
qK1EMssH9SbHz0dO8b9f0pJQNRpnPze20tN6WMPUqY0HQX1jLcYMWrqqdALIjph5h5U4y7ELPKsE
s2TrqSnf5/exparsEQyrlTXUXfc2x+uZOdgeTT6oWt7pqIW4sn9/8CQS3540pNEXJ2tXOYPSlnK/
uUq3sa5VEVAmncbr2FyjBh5mYvP/T4pe5KSO88yFxsTOCJEDJe5dqTc1TR6SsfLQOpTrg7Z9QTT4
ja5cPitj0QyAdAGWMVuo/k8vl9lYbJSmbJ1ceoQZ8BScN4zpIuVssXMmhWZuKh3FcENGVRZPQFkf
tzngcdeAXEF9c66jEBcdG/Z/RCj/KQDB8Jkb0QV7AozrPFv9YzJMOpPnN2arT/jSBPLOCeOQNZkT
X0CZyl21GTHckzm7Mv/c2xSLor24AFlqaiBivg96H6LksaIyL/+pta3TZcWxCtuMjebeaDMXi7va
hyKmqxzl44zoooVimelh6R1U+gTamisGYWZvlZtImml4ALLbovPOJ4fvBdqgmfI79yk5rR5AoOAv
eb/JtQ6EIp8vy1zdaNnVQT9URy7g9zXPvZnk/Gq3EM3/avCM9FHF52p82nTrwwnPcZPP9pqxtHFV
1lGlRQuJvXvFSt63zGf+lsi3iCkt6cKKnU2ae1/6ZsJxJT7o0dAjxzdGpDEbTjPLPAh7naKVkkPC
qYm1lVi3pgW0d+5uvnITwUb/EyW62OS9WWulcca1La1+gmzlCoUdLvpy6Yv3POSuj0dFuYK9w3O7
Kxt/jZBUttCNn1oabnIQMGFLdS8R1BVrgT3zrN0gtOrb/hoI2kmSpMyvfFRpjjvqkaa+p4wI7qNy
bWcxAs6KjifPaiz11qJHi9ov43k/l8eVmAcf7xjVTwI7AOFU+Rr7kaxDvp9Ve7pCQQSWx4ej9RdG
xFqfgfc0RU/GkSo8GHa7+RwdqhcvBLL+wKbkl3vJjzIDjyfxa/3j05O0BvJOZmAkjsIPXd6DaAPI
J+ultM4VrqgbjUIOfAbN9fcMjEIQoEq1DSrTxLhdctouYB0K6JaCeEBJZsZD6EGmdPx/bDTqZXm5
xfK1NelTy962B9m22EMM1svtedSc1vx8V96lMtya6GjmPVSTZUjnhV4vNEsFt5WBFDIeNgC7rX1R
E342n6ynWXN4xS8h9ZvbkGgWYAu1mnrLSW3ZBAEPvrT34WniyrWAp66SomdnUHfM4bbyK6SMkDo8
TTtz7VYmGNJmPJ/mjyWiQze8Uea2sXG1dczGL6IZm00TKhrZ1zGh7QwYZlSSRKK153ZsVbjEF9rs
LhB/KhdFQT9JU5U+Z6d84M/g9x3n2liiKdRhZ1DaiQXMtWXaG2EYic3kzi6lo6cs5g/3b/j0lgGa
9skWsWBB60bptRMXI6REf/UdXB66goNuh14xiWiuLmg3wA/eZN773TX3z5lzTaXA98THuOKWskhd
FLqoUQlbNrLcciA274e0ovTHUhtD/UXx3xo+NfKrIJUUbo6bRT4Yqjqxl0sPN8E1SoBEwSXM7aqH
wMn0ZhgCQQ9ZuhZ5n4d6GyQI4skMB0pLmnVkfciRyDI6u3eP6V4DIx1nSXVCCiFmZMN/j4uICYk3
1nPzcim5G3M60T8kjvR3JUb8oappMtyHdahKqDhZiffxcHRkpFEBuc/WRuz80hsgwgEwIclDJntA
Mb9nqJ9YVAdLjPT9F1wQ1VAhU2i0wkXgTn3rBy9Np7ulpyrr9t3rFVgtrGuTye8mIKvLf0FevxlH
6x2P/XxzyUA3NYphx/z0KPrBZIsVaNkYOU05khV6OCVdkZ9QrTUaYMBOtXrTq4096zLsFUHZacWw
SaLRQ+sT2CCW1GsDDm/XFkfw88iMHGr1ozK2TW//gvt5ufg/bG4rsExn4zMA0HiBCBDNjYt92qAy
eJru09V3sMHOuav+qojkSjnMSLJG9DCDsxSdlzs6jqplZklgSC825nrSeWOBsKE0xCN7wg0Fhcdp
iBo4u1de5XXWoqN/LeBENjf3Ta60Jf1msu556kxx60eMu4+1mljLrtxVjzeS4CmZpg7Zg+c001hZ
QWEkPSnDYPTeku1sne2DO9dl39NUlD+MK2nD2arXtY9m7q6TztZTRaIzoZ9NWG2I2k+wEPockj4Z
hgi76q/GCENTGOG8L/I+8bBSYN6Oa21DsY7XuqxVFang8gWyxCdjAhGuOi5vJ0nfaZfpBbyhdvc5
1V3pBoAJwGKYiKAaYrwCjPzWnyCciVmMZ/SI+iA0xsGJazgHOCyjR8TCBpvRb9hO7jzEp6q3JVPt
cvDqRKzd3LBNffWC8dzQGMXjOT2wkRGWOwdcYAmxYQNc12OkVBScvDw36Ccqx3+MR1qsqHs0qYpR
LC5EaMoW2OLw0CGthTjjWwfboAGPvKjxKf+fg35sctFYpTHTwjtkndSJTHlYGYnpuDwOgHAUzgsq
IVKltUldwxQn9TTr+vo58sNO34IzzmlUUSFr+Mjdl66wjX7UrjqGdXEyP38sDj+QkVlRRjFA42xf
LViZFi/PRNtR7zTQtFlfWg0Ojo5fFKwdt8v3twFFreYIlEFaFcOjuhy1wpge+xwWqkktrN51V66M
VYUyjgTJa+4hM5jZ8bsc05vOQcxC/EQx6DPoYXwUZbPNkRpoUC//L/Z7Oq1cTr2lxFbisRDU/0YM
pAUQOpGGNhCI9G7YZUOZ5t7BaLSFdVfEzXn2aFwYeOWyIwbg2xLyGDv1MLEYS9kbrryuisOta9OX
9mB6tldpx21EB7Fl9qv3bEXv3LcdRccS/H405d0k+Xy37g/mztZtLjIo/VgoDB0I19Y9kD7ashau
PgtF94fwCMsGJqVQtRPdg9POeA/A0OeXD+r8dEwzTG+j5GGTEEH/JP6qqF5nzZU8jVsMcD6aeY/0
O61Ht/wYm51maAzMwJmLD+YPNChMGsODL3iKRe7nXsOY4NNwSnkICie0faUCizHbXxtJZyOYYriB
ue1vgGsGcPC8SFjnj+2B13MwGJ/vqOwHI/yu0kKQHA3j1NCzrL99sVOtSrboU9NJunWRFqrsfMkW
u2rtFBrANtCymj+XK2QzjH0ETisXiTsT2wb4L6FkUKidtSpB6mefH47Cf8E9OLXNeNPDvm+PnsF3
d8WWajYMyhXe9Hh2Kh1+fCEhDVXSx2Cs7Jt3cKcPzkzAiy8SG4N6/O7PkasVEoocitUCL4k+my4R
DzhhFSil/GDMBtJ5XovjPOLHsNCB7yqKuFN6VV1aWsUiMSHmHD4jSYf8adpQHofRZKIMovTHxNtf
BwcEnYdHkx0iOcY5l56hEmdTF7g/zsg+wtekxIR5YpHJBprRnF8fzhaDkXFagm0cnx/w8Ay7qrl0
UiRQyNeSW46Qu40jEezcgsFnrmeFDVUQ+LKnqKoZdL2jPJGgJpirm1D0yuHAzZ9rtQWklMflTyDM
edw+0Av+6ZPKRNuJ4nBBvjMu9Xi1yYf2hN9SnRQSLLmq/iZoFMvjfDbhDy/A4f6NInXUJCu7OBKc
MX8WNDO7fcmPgdHXvbSVvGmPnFC+Qi70qt0QGRaW7LskZapZGhQxk39fEC5csnr0aKTG5fbd18IU
N2Y1pQghI5FJC5IZ7GNIot7jXz5lLsWo/MuyA2l7PiAP6A7Aa1jxMM4oCZWeV17wBgHGgpInvoXU
ATrLmZTy+IFteWGqqYp+3m6a+6rgIEp7XtZAlkR+tvRAlf8turdoKvqLEGDJ0LH9NA5EKMvQoi3S
onA/Vj6x1BlaqwJqyNuakwFN9p/BMAxajurN6u6IDB5sCVZOw5QLEpgQ62lbveQ1+LnryFoGSN2O
rQ9OMIGiD34fBuIhJDp8rlCTmvfHjWAxSCm2S2tu5Qkz0Mhxzzn5MH3vkQulXN+Q5RGiEyCtEVHP
8nkisK5xCJSEN01h0QLSm6hD4f3IVTLyFjDMle5ULJA03PDU9mO23dT/kxv/kxjcXxpoE8ylzIu3
pcLoazKEmOYISsT0ZICso2H6snJyt3Zb4JAFp/oqS30cWGfBQ2fKNdQ5g5iRVMxvvQxkAn/iH0H4
e6UxCaky8rDLqThIpDhOURWVxbylPc62W/mGkCj4a6QfQRiQ1G5JDqRxKQaiOErCZoXMAOP/V+82
2H/ywa1OaPyopVBLO9NC3928mVgfP+oE9U3j32QvKElS7/I4Pxtmvy48SoNai1TNu3cygppnOxKi
86NR4W/H+50rJn7k2Uc6pmOqzyWOP5pe35Oriu4zT6lEp8a0PfcfAzBvLFSm25l9vkx1D1APTJEP
AI53AjiEF1gwygkCVDXVglEieWEIE+MNbb14WAgQ++1gyKvLkVFu1IMgJkiiBmzhEKFyEnDTyMLh
0i2HruWtMYcnNI2Q2UNrOLZ1cxjK0llKiJQyjNVCnJlwjcEJVskIteWwhOrWnRr2SniJx5uYyC0A
3PSE6OWiZU4JT53GQ1TyWf6bmTgqroVZCbCqMFHX/NxHxHEXgoaDIJWATRlZxRBMIt006Xpwo4b8
0cr5zOPw6+F7RNdoH4YkKNHMLTa8z1K8Z6qjmtOmWGoRK10vveyqqAZS2G8sjfxxwqyi2BlzB5tb
je3X1xN1L8W8RmN6rB6o/oGCn2aUbDM+feKfu1888buPYMdrmVZ9KonY8osxAVPPf+tYEr1nxtjm
H0RvKLYf5nFMZjNPIEUcU6qfG+5tFZv/o//2M/8PwGTSmkB0Miups7vQ4UPrN7n1gzDmCgLj20ll
3iq/ZzjeblKGTjcem2oBrdKpF33NMOkxRRPNGDL2M21pHcHlKXdtAMqGSNASZN/oZnaBf8A1k7z0
Owk6gTZNRHYtKp4l8xlZAZrDFNqrhiNWkqe3CCeygfilvLKH+/X5Q9W8am6aFbgLk3HCyMF9BMNN
6GuHo9i5CS3ajCPPt+JEszfYQSSZraV0O3VTCkxjA0HUnS4nkz55vSyDfsna94kEI3CmSyL1P0V6
uCALId4l3X8GNKhpbWEYoRL/WImLhQjDJraeHW1ArYiPa4nrGaFqDBaEGvf3PeKa8QM/PgAIqcdt
mtGhEWVvMv7Cg1KJ3+y+ZMbJXm3KpsL7gHQDTV6vAIT7Jdt+fa2+LXuCVg7wn4bi/7t7dsdIty7Y
YygIogbkxowbHCHI6IsDSL0D+6s9Gg3Kwl1qagpT/VmCS2V++LHR9UJIzF2e2zRsxsgM0FBOw8Un
fU3sr/aUCiYLcGGWpJwGhuGH2QXPm3wwtzwBEl9R7atmPEKtgHizzpTOjLo5jq33isNNmSOFr55X
WsZg8L83dhEPghxTWnHKNwhuLPHiIUbSdi9VOZC7Q6HhREcKSL1SLzbvbQ5oLey00n6aG3jVNXl5
zuvsz1DJC7SeHUjK8NfTFIr08siyjCw4BKC9CYEsS2xrkB/lp2cff3RPMuN5LUilD3jUYDb2wAd6
tcoEKSN/jmEimm/vmUFDATu8TGcQzqpdUk0xBPoTTZG+kx6kJ/oKSxHa11rOJci7y2V7YkENHUvn
gT0oxO91gae1NyI9kHG/t8j2Ib22VZwj3lWT6d+qygOSFVjThgKGtyRevBmOKwLZwbluCWrJmNjX
4AJkz9+uvYhIjldwOXBUty+4I4SSY2dyv7dcu7hXBhSQZJP3UM/ocVPSEa/+vRmOtmAwWahmf1Ry
bwbt2AuDcRUXxv9oEkPRFX4sO0splIOaG321K2sF1JmqUQHi5/g1BrDcK2BbiUf8oIcs5mra97xI
HeXDHkdEh5TSdlOyNQC30VEo2JCz5QZaAdEShuWcPybv56UUCzCvCVZXfW8C0YzgKCv3goIC4WTQ
jPG2LV+eNfqdQL99PvDFLnUBmZscpVdazey8ZPhVsBEs8NCwBPRBRvZnZ8XZobO7O9Pm53Bp7xtM
GtDFxMio0TzBSCmbbG9lGxh3u9Djm20iZHazJhY8p0hmylylZ8KMBJIBClGeOfMnVQunZt8n+2+D
1ETyVxrvwYBz9LMZGwBeAZ4VqI72HRwbMP1PR6Px+jB1G2MUZkloFFG0Y0yYtSTnHdDc6Xf/qsur
pUnsoIVn44j4T0Y7Z0JUVk1V3UFHncaCxnWgq1hByQfR0j+qx2ZZQVtHzmQBuTNfxOqveHqQNkVx
2MElzsETjCVvx6IYD/yTAYb24fjgwLXNX/TMVlzIUtLcznjEDjt6G4dbwHPmU5URd5afF+U2/yAo
e7d1YERlEWBibD521G/EIk4Xk+q/B1+ABjBNPpVCsgoPMoqyBMmpL2Axb1PYRdd7JR968IcwEnEu
I/cGOPwmOd6GbnomG+0AsRZ9kLNuvDJiEEG3WBBs7Fcf8N4PEYTn21j6qYYwXAnxwkHb1I+tYiO5
ugsnID+//u5SOFoCxROQ0R8Qqn/8njuQXqj7c0380ddsCNwZCg5lLv+8JMx33Qhpm4+jfdJPOP4g
z1695rzQPX0JUDSIrZlQfmNKp0xHjuPcb39ll3KIwZMIPZI6hU3oWhAWRdnzLGX40JrmV1pq2C+u
a/Vhiq6Jt5LATVKyOh/oK7G51dbaHELQUefI8SBT6SkP8LNx3dPz4aVctj1JczWnj/OPOWVGwYHl
opQaFwz5w77wqNS3R/dhJPz+/Tf7mWNumeML56Wks6d3Wo7jaZRnvjg9NU2RRvZIk+YKR79ZDjgc
0cTTWmnlXqzmnmvTCICXFvRu8nmIQh3ZFkW1mUmTgbglDwCi6p88OAXZCZlONzfjo6XsDqX8HWxQ
OHezGo1lDwUdgor/7/cYFoUwhhTQZqtbCjqoI/iDzcclnLLInOy59T6ORo3xcsCq60c9024cb9C2
ddWdvQVu1jnjC019sdNqe+I2bfLh1R06lrbXU9AQgoG/Zsbb5JPYijs2G4N3RSa4EFRjI/+U5bcc
RfHwA9wgNlajzlpFZ2jHFDlh0VUczs5hyVrCYIRAxQhJeZ+tgVM6iDR7c4S9W2aml0VsEH45+ciw
45+Sxxe/cB4u74EPkUrtp3+6dR6zcKVmqxm8Z3maqUOUEgiSiyny8IQ1zjiWko7EgO9d6hjE8yRY
nfA5egoclB6a1jN15/w6PKe6jPyKJ3a2NWJzX+y+JsJa9Ej8uCC/+J4kvT1e0UL+7MV+2wpStFnG
aiONK/JyZeVCmkcyYWHPSbtQj38nnB8+cbMz3OH/MYr1Y0XTMYfeWZWMzLRRq9VK0cT7PSJdLUc8
0Hrbe331jIn5n63VsjVpoa4O9YwoxK0937Ej9hpyI7WK+D2ay+Dx+iagk3+IUKTONPQcNrABLSXc
b20tk5KNat2gLf2VxzJyv671jzB+BUJ2edCY0mvtUIjwHSgfFLRibgZeI1UILfTNpUY78tYRNOQW
iwMQEnHw9jhPMwohTHoYf9yOvnD/OtB1+IPtMCb62Dy75NKzOUI/AhgrjnxfhGuQwz4QvOZX8RI6
VH/eJqibTRjm2LsLIRJjAupgMgQnDGhdHDeLZmbms3LWtGwC1qvvOP0S6P6AbXJLNblj6i89WNQo
svYfZdIPV0rCJW+2UK9vqvoMAJxyVzkGtjYQ5B/dhMSZZ5KgluSjJ3jpYZO6uBQIV8DNuTDVP61z
Em3dKrDL1auTbTqE0OmS+UQAnGCbtTyDCnZiVim4MA7ceZ8zP27Y0ixx+aPK9zYDv++BBkxi5HZk
DmLhtYZd0xSGmqNjA2nUERdwikCJyxZxMBnOeVwRmlTyny8Ct7hS3m2TU9gj3QIpQCVGn27uBp2b
m+OzJTVd/GBIe9p72m9KKtqo/8paD3b4alK+VJBju1w3PuFSGZtIp8b8utP1PN451BmK3NU9+wQq
5jBVvO7A9D6k5Hzeq9fEJUnT1tUpt5c4adlTD8eAbUj/lNAoX7LwsGn/aFuM94tmCSJCKHrD4Wgs
MnsL1Q2+uAbLOxAkmpfboi/tWlJoJ7q//+vioJF5L88HeJ2OvGui3Ud//OvPHkGHgMJIWTdlniKf
hkgOzmI2TwxzSkzqD9dRYevX+yrY7cFAOzL8/53Rp+ZCcWJGPvytCktTlUM/eAXem+MGw/wy/G6b
OTVZJKIpKAonV6feM423FOWduNRvP2NKv5fBRUvE77oIxHtkc7TzYHZPFjrbpjrsb+B/uTOiKXRX
EHbioE9KTEP4w0TmxrsXd4itmRkP8DzTrvOVdKCQdW4ORZJrSHzVu5/7ZESTB+sbud/YNXje1six
96g2s02Gl53yP+QRvq8C7NBmhCQWwwWgCxdJJWDPwehHLdmehqWLYbqAlk5fKay+Cc+9bsUXTDbZ
HvEaFvUaLgKrfrLO3F6VyR5d+arMBFBKrCxdM8NMNhFlzyWZ/BUjPT7AeMM/C3uXVDetoPQnObw0
P1ATRQXef17PtqFEbsTHAvnHH1Ir777032mlKErnLNSGCMEKOBTw1+Q3ly68tV5OuGqjQrC5fFr2
2X/l2HNU/jDlzTPBWvTnLK7XBtDGN+ZCDTxxhk9XoXhZOXEMAjGjm1KXZDf8CAz4st5nQmFxrMIK
Q43NFCZ0lT18HB3veNQKX7w9SYN6F5rwtZXMky/YxVADpTlTwRXDNekrU4K30Nv/9l0ocoGkFl3A
kcYpIISgcTs73ePjpbo48k36j1dnzOVLQILZO2JN1yxBcGhbwXoYUl9rgpG4Z1sCeAs5iG5hTQQ8
tqjTHKZtKWmHZN+Tk9ADXlT7Jz+ArlgmpHFnVcy28Chv0hj8+QSVjnIr9kcBq0Ii/r0S1Gzq8Nx3
XV6Ccv+xeU1pXfGovcGuZw0k5VEs1I4MnV22LfcFzU/2BULIGwIqLzz5rfFcooVR/PgrdRCjinFv
ZwGaRsM6uDr2tPaBJQozV4W9xJHDvLd1Ug9HqmYg/0FQ6uT/f9upGpzc4tCOz8PIsRbETqyHSfln
8lo2U9E4ttL4gPJvasBDVFNoH2oQU+tyFSfPeqInVgPKY30LT8YTsSW9rUqBzCmPsyYcPqak2UJu
+FUIIrMeo2jGYXc/u6A5LDJyUWzdfyZtDoPeiKI5mlgIAmsSGNVRv6iGjCl6NUBJBbyL4QHP7j1r
MKzSYcEG+dS6d+KxuBgWTg3tdKK7OPGWHKcAX8jyOoODn2p5j0o8v2uUPJy6reiJt4V2QblMn6gO
W8TapDhq92t1DPMWcJYw3S1zboJqXhjCx+AjoS7etdrhzgXK1DO4pBdj0Ts8ZJOa/ETu7zROPBuO
rAmLfvYvAR6zTVobP+N0npEuEwxnNJOEpSqcuz8+MWbgoRrgjvgGB5PwmudGHDy4V/h29aA26yIm
MwAIXteolShJVXlKqN4pLMFjubyq0ZEmhA1pjFtkGxCVfv5lYmhPttLfM/MKwwaqUXOEPhQuw6xT
qzGo0wJTN4/x12wqtkkvlTJy1Xpqnp5KixDeNbGVFsOr/tzJToS/qgoha8RocnbtrykTKjUV7RJi
ZZD2J02jCATHtmmhPkI0lM3nJnB7sFKa5J0eWlH4fPd8OKHDj1mjksMg16z8Vqp015zfOqUKqbxg
5cqbuA+q5PhIsYz3Cvoavr7FUqoKxBNrJqsEX2s2mvT1O6WzohWJLoFacY713YrIB9nopdw6dOfV
pI5nM9/zBJK9xM7wEI8FLUdrM26tUDPfblW+L/A3Lxm+AmBmbFJtqLadig2Je0ULB9ol9pPY/kWb
BZTbsUKlhgCfQKbp1ORpcgabPPH3q8e45F7TY4PHg8PAu3szTlNZNRsaL497UrELhqbRvDYP/J/W
4MvgEO+hdREujQmQ49zXDJlFMzzjv7ShmD2W6j7Orzm/wDnWNb7U67WQJv6YsbZrIM4eL/0B1WgQ
TB7qfrRNlL7OxOpO+QX8BidWDbhubcfWW79dESWxxDfC2AlIlLBu4N9LnYi64oGUg+Ctu559Mwg5
n2ZLQLs8X7rdhZ3Pne+1EJZGWYFc5TgUpXMDyRBQCG1ZVVRn+jImCKcRPbjjUeeWb3s0PRoBoIFw
1aeXNXPydX8WpMuAM4yL9MRYsrrgJLm8b7eT1n4vUh5NPHCQlyr33sOxYeLTe5UUX2yt1KPvCvGW
JDY2mzU4iTgSTB95yGT9qaptN+4n8iL+FbyCT3uHv4m8doQGjDO1zn+2e2t/Nop621zXzdhW+hN+
UV6Zf6Hbfq5Bye3fE/ny51auIPmBSSsyuQfk7SBrgoYDiNN8M4HkVBjXu7A71wpZ6bTj7AfQjp6c
M5cV/MnFg676vSbj44+j0OG4TZ1ApdsIKlzSmsU7udbjbD3X+4u0x8HNPRCpcXj9Uqsnc+0zNEaQ
p3Ey9CwJHmHAeqLGK/Pdsp1B0/879X4VgyLViWFL28YTODHpgzWPLB2l4ggae5f+E6R5Pcl/F/ZO
/orP1Ac8RiLju8THpqy6nwWcPglEpdGh/uWzWDGPG6avHVj1t7EyOOsQujjx/VZtqXMzt7k6nqlS
2NsfAiArHeUP655mWStgukQ6ZiNVW0FuiMSaYh3DLbE0RmbkkZkeoCDF5o3/DF5Ld/A9nWwoMEVK
cEhB9DRQnqWoR5CRZes5/vIh8v0YdIjlUXUbGQgNWwctL75qfc85SDfDI6oyGHI3izkBC5tTkvXD
2UinlvogNTp0L9LQ0WAaZ84NoYMaFY+XDS/odsu/hAQqDWDNpxy/KDZcrhlx73CBqBkMzpVzecS6
uYv4pNF/pFeghkKYCCUlAe09QHP8ZFOEN5vZzOpdYTXmJ3ZWLk0EsBUoaHztRyrycpjgkRLPBEqK
E2z4x3gOJpVmnGEaI/PNY5k/fhbHzvUQ5/ypFoL1uguMgiggFlvQnhsqQCgqpuUt5Oe3oXGEbtj4
QOmmTH4G/u9TMyiU6Kc+9RJo6uTP28X7cD2sNZEasPcTXO1A79ZfD3XwLnYtTnQ/EEHa4fWIVc6m
D7nx6yl10Q7CuB3IWiZjFqEgeBGIGHOzu15GUS0/Uz4eYNXDFUtzC7nPmfg//nZ0CIm1CrOw9wKj
3oQ9e/a+NI6UJ4YDDbY3PNkbyRBURLOFqHtY2EpfyDTwy6dcOHRuDzX2gELeKL7dbLYotEVEfjfE
0OmnhPfNWZBMZ9SRt9Lv7CbprhTiJgj/qAdvqOzs8ezJ2BQlDDzQJ7TLj/WbXUNCS7oaQ/GKa8st
pJCkK+AQyzpO9myn1BxP8EPnPi1Gt7H3zjqUPXrA6R73LJq+tClde58+nGexWSqEgh7qq/9A/8XQ
/YW6Du1Up4gefSDN74Dv8xoB2HFhVfx/m6atqwsw+m4HxEjxyHnLUhkNidaM66I8jjBsn4qMBo0z
hf2Fmz+1hYpmagD6BSOd9NgJ4tK6urrpKrQ4vaSkfq9LDujnCHEunav0I1TVKPdA1Y7q2V+2YbZ0
sopdE+kfhmR7DiHHm7MItm2/U/g8RwnbjbTvqCTOv1lqb7HsI6DNJNnXULH/xcHdprcbw1juj+x4
x/6fkM5QNO4ulScSVLCV8VMdxJd9WpwpIlwKFtuZKsyuNSdz42wzrPo2WiH8tnY9sTdHtyU/NCqg
gWWpivyrcUI3HCkRFTP1WPhbpXRs0HsbJwuIcQ1ecGITEvj2dOYiQGPZC1Cc9p4rCapy5oTS1Nnq
HWA5xUV7+9vCD95QbLyviJuVYfGx58+BTVo8IwzAQgPkd/sJS+hHsEi4SLYJ/bCHZnvPf7aKZb/J
PQrGpn3WxELFyJ8zGvq9JHA7szjDzmG8QGoKsXoU4H0/HPR9wsY34FPPj0xWcs3Pp1anMsFq9aAl
oRcR9wD399jukD6wnnRPkM/evbnDqY9MdUpzX6l7Vus1vlCxvLR/M4P5PGex11wCapiawloFKIlY
suzgr1jb53CxQWtVZBrI3meptqVA7DjdnsZBsaLcthvhNAVx0DBQMMiURiQ7HJsK1p3aM0el5zCj
kaPHEQgDhoAyNUUSHGAteJupapmSjhXxHnkEYqefbQ2d0fRSmVrm9Lpv7a0b3J99REqoEam7LrRc
zuckNi9FAVi8BUsdtXf7ej1xeXaS/0RaUGVDE2ATq0IGQowFyjKiffI3NSTa3WvPXOJllptoGBGV
5+7+M0tI5sSZEf2ao/NSZPAhk3Y8KCnoFZctZT7DO9otb2qWNXzBREAIdmNPLMlW2cR5cf8sYg23
AgrvtcQ7UZyGAVHfA4mELU48GrKTDD/FJGsd8paOXCZmr+z5QyaUl8blH/Z9fKdZVtgLnKQPQzEk
y9kLByN8z2xwuai3M2xQv+Y1CXqG7HOXmzlFSvFTNxBX0hoAkXjlcXPbNZklRSFyUzHaCtsuAJaC
Uck1H1tHom4XCtViduXrNwjeZXOn3qdZxSEoyNHqc3XdXc6Fm5aXIocbIBIpSCuStANwTMbzddAe
KaOa4/py+Vz9fh3K7tObMOWDFcAx1dhO57e2VKtADoKpc/M82RCs9bxHb9wv3UlAUmbDp4J+dJzY
bWcEMDdvp9roKFPTcupgkcpeG5z1f32Q465jQffHm+Hxbunw3wHuJv1y5pIX3O8C7o9gGCMeashx
ML6lYaK6c9nHKFDK7J97uwyH6X1SKWKYaIKEub18+BFcCATZZKyUI2jh6/AWkfSgGNTw8czXBflb
HpgpFuQs0Q4xGC3B+69RCV26JdvROXkX3vfvWeUzcK+pB4OElu98a57hi8PyygKa5/JBVyjDBYkk
ZiCsPaOiJ6MrCQ7JPH78u9e7jfgUczyA0HJV3z7qoD/yfssuRGAtVIRr5H14OjF7jklDWzxSHSTk
/sMUVUKYF8ZsHL3WnuDwqIjEgP/mZVPUddgz8nIxPm92ppzONZbufhRLYTUvOmIXP4cowLJMsbnW
2rX06ZBF9YhY3aL/do/2ytUnfuT2m79iBjG9ljH1jQBfwDlW74lMLXSn3ErKmiqqfH0G0yMy9G3g
P2YwYDlhRdc7DgezPApGUlhmMPKD5KdwlGWmbZqvsx72COWbhLgNnuzO4lmeAwQEXXVcCTc9bTk+
JGK+jLWQOBu671nTJXYnlV3LeL3mjKzV8FeLq2dGBLIhzqU+BXqrIRp65mhOwnLAfHrW8hU3OiF7
ZITOZU72HpXjxKl7tWAj7ABWYb3D65JjftXF8pBpRiaHjqFRZ0Z1A8l9Ed49XTTrsXwfZrN20iM8
nK9WuVdyUTY2Icta6jniRQ/6fdeeYE6dDeGKzbeb/KgZbLH2TjO3badT/D4O7raUUNNpF1KRA0Qg
xgEwmss69C2Y/+wNwau0YxKigczrJrbv0QBZXnJxPFlYkRkMvpH7YEfhs+fwvOUtweQv/gHtDBsH
hHI9KpYfJLf1zMTcFcma1N2c9DArfrn3zZum5cdq63XRg6IE5lyz5VynBu+7+wmEFaw14tjTWfPz
RgF7NoDVxEM45zuNQyzRORcqfEDPmC0lP4Pjl9MwePcxDEP9ufM3hTkp9BHP+fpGWxMp7BxKnrU6
0oeEwp5neqtB1XqAVb8Mi9GqWiLF/e5htkx8z8yqoH2hsS6D02m8WMLtdvKOOzqtu6jO1X5G9yM5
aaQSL9usu/Mdr73Ip9enCoKr7sMJ12UPLyXhDlzGm23v3alq5UMs4QRlze55hjM/l32CQ6ZO86b+
/gCPvbGTT3eoQ716OR40oBg/M14uMRd1Ro0eg66BTqXafXeh2fJUt7Mp2O51LNO/XhMFd24eDiSy
CMtL7UljHIJpCx5GoIqnhjYBcnDI/nONUCkl4mCiNe1TjFzPYTkN0IPuDkUWhR3YBfAqKvJc7H1n
ZpoWrzDB0oMOkZ4ya6SQzdbXqqs45c3kgW3lJYN1LV0sh2ayx7ceWsYcN1hcRKrkjdbHF1JvCPEw
1Jnl4KF3xZigd7iQdK8THoBKUyRpJvNNCe5Xy+uaIQN5uLnHdiILRXGr6dYDSieWtdb+O4wbhY6l
d44SJUJAy9UUell206lKZIg0wx6CMqaHFGzOmyj6AumkGkE0os6q36CliS3rAMEwoKqv22jtEOQQ
FjtFeEwF7SBNc4195m7NTRw2HkyQuN5kC7tj9AEW6FzFnBfBpWpRlj3CXTJrOsEX/92NeCaWZLvh
YOfZby0m2FEGaR3LKsJPDRYHCmU43yuZ1lHzzjo2aVGFgtG6OKneewlwmS6aFeBW/ewJnjI1t9oQ
jKT+p0lYri+xEbpNrQDDtfapJzZ7MRwDYKhCtwOX/j4DX5X76x1sNic6bj6bItBWIep3zs0Cczbu
+O8bpcYSjLt3U+hdHYAnm6gpclpNgfstWObkxTBY38eTcpuujrEfKgGsbXrTSggfzfyM8xnqqMEU
tlmKe9YxSMhUHQf0/IXEyi+Mdxj+eoKEoHtQ9FmPjV/FOzzyWIMh4/BTK3BiXhmxRz+4fd6V2Mi0
MkjDjc78a/fL8IBfBwHEmDx7kcPxVoNjcc2OKqxS9CyhnjW1dItpAQ2MquI7EfBI6cca7Za3/LaV
pI5qJW5r+zNt9LVDwYyfOElv6ijT08cfHxzsg3lWPbI3qxWdVl/hC5DKuKGyvNTPmeSPk8GtguEz
eBAeZrHTdktO16MoZ1PgSrusvZXsYSaLVS+xzrAK6Nw/jOGcT2czatVvWNd/pfEcFzEnTvwUeR9d
JMMRjhwTMkCjVeT5LVY8wl0d+984kdqUZmn1arAMmoPPezuh0Irz/5bOJRD6iZP0XamhG4blwWNW
/ZTpe0b2ry9BifTZk4nwvnzhBw45IA98ucjTaacA/mNr68Ba+WLX91jg/xsCfeCogmyQ2/d19NiV
Nzdom2Y+wJ1/NTqJrhjCqZmrY25zxQGXV7DnDuXRbIHZw7wyB57urexS3ZJxle+JNiyEMgngpqw3
RdmsAR1dJP1aV/P5/FJ+vkuchu7bCFAawQH+TdN5xiVr6nHtgLCdyL0dhPsrnASzTerTycWGCbBD
nRbpoVh0gprnLgX6uNbCC5nWtxEbZqVAKSYmK8xAxkYyv0W37tth4yxM7g0FRF4VAYftCNd8gb58
PvSrVASa9+1MOi7r+/QE7zF+SmQh6oZEe4cs5siJWZpCShrYs6wv3P1LIvem4sUZ53Llj2iUbz+/
fSusk9QszoEVgf0aNRzu4kKpOkuctwtL5z8R8IkdvSk/DyrfV/5bCm23x/TB0uxBkr5DCqKgyIMf
R/FS86ZUuIBxFw4H3rdJagy9E2khou6AHFOR13KWvj5FmPRQAA8ZM2bDdY1AqO4QrP+4MfvHqSZx
mbrAu4n3ZMnumvqUsfGLFSr3OEQXnwkudPZORZqP5pK7ynPDp0Ja/reG1MjLijrIXzUUxdPXNnMo
Q2WbgmgMoNR6jVmx7LRSxNtzqD9EGy88A0SVHAmYeiJkBoki7Nsb8xamsf7C4XNl388BOnzlv6xr
MEEQ8V4nP2I1Eb4KOKf3WzsR1ysq4miCc5QcjsAirVlZSz9uyb5sWuZBiKNqJM/QgCehwxLxFykA
dTZCAntj72NY/6ukrRjhCmPeEErs8kuMABIi2aDf+avULsxyCnT/FEYnFYNzoN07X48BCmV6wRDE
EkWFpeQtkrUWYBjaUEMKk14p8/TyheoXJODSYZoScQu57Eb71Mfz7Dj4HQ4ZOdTzqDRQbmVl5rEu
c6TtgSwZyzLGtpZm+8hhLvxZTn4SpzzHeMEXj6ydum3OsTBBZBwGOTFLSuSSryOQxGQSAmPnTxgr
T5m5V+pRYxzWMMSMOuJLSxr+bgy6g8OJqarf1oaZX6kFgRr0GJ87fY4cmI0RxHorQyGrjl7zKIn3
UaBPQ3aABISN4J4K6sHcP6hkNHa95hdGDBrOsUtcPnjdmD/K/3lsc10bI+Cegr48pGXC4vzj7cjI
om0MRDnXRslxu3mIE/c4rgLcstsger77gZIlrPTfaCYL8GcEoMlgiD1TqvFO3ahWdj3LEW1rYm3Z
WIl0zqzWVrUqCT9xJUuUEwjDv12OULVkPTQafrpI/KRrer9hN9yMujmfMT34Maiy5/JTlo7ySAK3
vLUheUUCjLYsYGvHcxjUUn1MUwAGfvJECZ3EwM5IEPsPKfTEMrgT63NfJdIQ0t892DIwvFLgJhqm
eIwjoO5UVu5CDLlArEsnoP5Kng67gIW5HHPyR1xWxNvAoc5hvO8UibGxeE95a4A9T5+Yip42J6nA
emk1qXUnnNzcj35OokeEtBvaQ9WF+igNr4jZkNkOHkF4+oqGrlHrsVWr+kKHXB77NyAiEM7oyZH/
yDJa8jG9CBjvzBVfFZRmWk35ITXoh9txKBlGRh1UU2KPQL0eDZUVNaCz2XA95MJuG5exf0A2I9yp
vfm+yBDd2XFeRrTlrYa/YX1acvHUyhnq7uZGNMy8PAe+X87c5AmoNtVDMh1mBZGAGhzU5+Z05mSx
XFxKJ71hC4KXC2HteoYOat1w2TOL7OOYvgxmicgMUPEUZp3TcZFpcHppWoCoJHLoDwiFMwIPXAwu
jRIU+8HN4Yj7uVIAuhbT4eTCxaBMo+VZ0FvB5YuXo8kPW4objPfzzCXFoR5iwFmV7qzWXLI5ba0X
dh4XQbMdtWqJjkDkE+RgfXnxhKZIUrkEKCAzSsP0CcCl7IthBlNbp/sQK1xQMWPUuNAKDvGtaHEe
fsVJZ0bdfQDbGgSJ0Aujcab0av+ANt3o4a1byTecTCathSM7ybacCBvsTcDTYOZ61bABkbWOAnuE
M0FrfpzamxqU70kbDxWkcLwJctztsiZmYbwG9eLlC0z4DNzbJtgrYFbspgDTfUhiDndse7Yc+rEe
X3F6eUQ5vg0l5XrL0u28Qtvn4hky3q+NfhzCfnZRY1IW1idrHS4kJEhNiulXzZCgzHwgc9vQd1ce
nh9GgHVZXfdg3tw0gh0sxSYW/68TnRNNySwEy3oa1YVIFA5wuhuhQvyBFD/237+3vp9S55WieBgK
ezIb48YjQyDDfvuTDQ6NttEc9HRAdfInQQ+1Sb2zcV4uohWWLu5bdHXgwLSWgi/xGkAHfcufeDOn
Br0+cBm57ghvC5oIijpIF0ascmeZfQWB/35f8MEWSMl5xEDopxRhQ/Tu54Pq+snB2UXNxqDyVK7+
l83Yquo0VCVQ4sgTJFO99ea9l2Q6q5lyjDCAx40r2hdof4EoFMynMKUizzGidSRDoBUcg9WKr+6U
aQlOHbAf2wvR92NSgce9g+458H1gBIZnZvkujwT4VusQxpwRvAo3Hp/Fl2teCENFvg0bNdAsdgOI
YKLR85czs7qQL3V4Ln/xex57JxVW8WnjD9fgrGuQYRY+AfWkC+cDzc3HcG10CtUJbkQ5zBNowKbP
8Cz+b85XANI4ek7TOkuN0W+836yfxmodVFQvS8lCZUZOePqra+p4c7goFaF6bsafc+vuWQNILJ0O
HKcyHtxTCUJqh2zqfq9FFKjt8fporxftiB0E8Ht1BKSey+M0Xlm30bxwFoRzp+kMeSlmpzlzyC2A
EmfE4m+mBh9Q4R5cdsKdTFEn4roJ6/j36IHbaT9PLHKswSoCYRVtisJbDaxYvCP7SvcZctRI5icZ
6b1QBkKSL5oLyj3RP4eqx/1Mjud5h3xTatYCZGchRsIxs6cOVr8ICFSC/GiIssQAzDEVUDEPyFf4
3C1+rYPiO8D4dE8zNwMCC0W8oZ54FQw0IkiO/Pyxj/KVsRMyfnUP1BEywW4WMkNxQYFIKmeRcnjP
CD6A+iQBsOVjZhUIuPZxEmFTLhp+gvP8m/i4L7/dzt3H3//QPD8I5kzb117ggSMAz6rq1kIo7YWW
pR3fA2oU0/dbnXOCqeNTPZ4k70RvdBYshGhDVLpqmS5mjgEsUQTlQOqlamlQ85MVbuQTQl8zC/15
orAus+tuULUnllSbhCbsmU2gPQKNR0DIjlLsIr2R92T76Dwb3uYXuCPndL7wkliCQaVOsMCR47h7
1qZEEEKxkgfiA19I1gnwKAgXQJhnR6adSQdcp1kfGAWz9NfD2vZzmpZXCreNod3442X7Scj/59eg
4JdJrcz9+umyBw3nOSyIiW8WWu2kG4im7T4AWTghWrJATztAlbBxUYvdG1xAVsAEtqIqbkeyDlxC
zao+XiN3OlV0j8GTaqoC6QOcB4lfLa/SG/mAUOQdtGyIyIgYvr1pKlsj+gbn6SqZBb9LgiDeLpaD
hM+Vd5PnlCiTDAYrUK+mHUXaZRF++SyK1hPnVFuoGR5+9J2oFORVmn2mUzvnOi3+hwhA1JX6xZJa
+kDGxXVGWxwMYKuYqHBguceI4loYE9qJtsgRdNLeDZTdJgZ+PVehc5KWp2Kx8GNj1IRxk2Ulj27h
T4qbfD347yT+zjZx1vg50QolGYgBG4gUg3FDO/jDKIdJP1zofw0CWk3OfhXzBMRaPkZ0Icql7A4e
aPTv4jKTYKLkZu9nKef7r9lSn6NwSeiuhYkZgSIcv5rEw4pCHJgYuPHf0L4Fbk/8MzBHoyCWFski
6HyJbg9G/jp5c4DIbDZqmYec9A6kr3wFlgQmrIuTCNIYP3SaHWs0t+S7Ad+3XqOFuALMig0Hjdv1
drCMJODSlcGnILhXBaPEia//bOsmUjyTIpFk//iesgUcrA9eJxPssIeVFWNaR3qOFs1fZXDfS5NH
9zQC25ahLGWZKI8FmjrKG0LEHYmfThgqxC8r4/ACyBJD+FQ2FaI54hDHNujljtKJUPepMngNE33s
luxYIS7o5cEU2+WS7ewBkGGeSSyq5XcpGjRl9bAoM5CQX5PBaBRQAsk+0U472lolBz0Z++vd8Ava
f00H4iWEVMhvCpET1uGx1c5+vZ6HB092Dn6uo7KO7ERAMiluCGd2JKuUYy/4gWWqZ/132+UFRAT2
ObAPkieqk8qx9Hl645/cxAQzLwaXJ7XJdZmwi/iYf3vPF8LsDABB1LSlsFm8RH+g2B1YmMotwG0z
okvLHcYun8HwaoU1mK85O42c+Xz3mq8bKoJtpWKENM7KzabWOieba5ent2luVQM1ZQcBu1ZChwVD
pzUS4WNsTjcD2GH9HLSbiM58LqOisMb09F8XqAdJ4bXRE5cL9Di4Qd/1anQJFoAtb1ZOs0WEBXQ4
p3phPMjbUAAyRdCwahGckUqc14X1iDLoVTrMUZXziEei5ajje/xdD56sD2eL+iwAuDCKV6/Kgf8r
4+tzQQDFL2mV38U9pAUkDrBCSBVmeRFTl8Mp6xS1tCcomA0S3KLmH9rS5DUOSPNZ8VKhZxh+BxnK
9zjMfavJNbf0V+h+F3RKo5rI5UIWLk4Yqk1YnK8jov4KLZIGzlPGRK3liYfDlGCKVZGOw8Cqs6G4
QUGhyTG27UHBq0M/Up18zJIJCrY266MJOIIntx5OnIO6PlOLxv6WY7vM2Lk63CCTgYn+RFWw16Va
cwnZK6dvMQyRjee612l/LMouLU4jTdTmga6bK9YTUVLbEUl/V9+7V4yoE2l1ZBswcn6HtawaJug5
n2hbbksvsua4dx1f62rvR/kH5Pda38rTZCRkFSEHtHs2sI/HvaWrP7g/903v+IBS/3+mOyMbqnKy
ZoA6quyw05sGWOPuEdHoxO3Ph0lfiU2BvJ1PGF479ucKhOfz9JahsOUMHHnCOmM0XvGdYoBKmHr8
lc8e5XZOlhSPFPGJnn/21b5p6Fk1w6b1iRA1pYIGZzQT1ZCjacjrKJ46S9SkynC+wMJO3wI+7T7I
yCLs3gzEGY7wainvEOiCBjYpWteP0wCvE2qrtJin8otZ91QEP2SndYr1Q6N1wZNjisTsI/de8AKc
nCVNK8htDGuZom8UosxvC8C4CwFRTREQZKGfsF99rNkEcZaTeOhxhkuQbVuS5Z6pEGr0sUBCHtq7
zSaPXT8srDso1GDDkIaN9nwsVxQEHqvhNj17HlscgvkPszzxG8/f75heh8sHqiOazCy5RcMw2iC4
MpWguTMNuDUtL30NQEEq7K/s1VOjhwoikxX5Igw4/PUIj9IzhW1uqeoTtSM7tJ/mgzEIhJfu0Kr6
U1jINcdBTVecYyzVPy/uQ3jgIke5giQOUZ/v4NnEQI/hC9uRcWXQHyjEuNc+U0ZAR3ssXKqcnJss
ofIasHzB22OjodubDYQyxcdMTXX/0t5uMUmjPAWKnMniY/N5+hVX9KTWC8QTk9QmH9eJYiDn0Dcv
o+N+VQQk0MP6ttv3K5DLbMEMc13CzdbrjtGm+Hx3bG5ELH5FsuDeLOnSCxvWQWIzB1t5PiC+8kV3
xaOenZJuRtCRO+icgv6qwyVJ/LxqP8jfqKVCdCD6skR+uOLpiozRskkc0LZcfTxkntCncpaCHEuA
sSYU7qOcoCxTGYFwRIgc/BpHnGndmjVKS5cy22CXrNZdmxqn4c+0caWGUMuoJtiVtgvlmlG4rV+H
5S+zTLXo+LZ4NRBTQH+hDcf2PIwaqIVSY584HfN15xSKlM/CLOEp6BiijJ2i6IxDMgdL4QTgY/dn
MQRrMtg31HD5F9iQPZNMMxRtQ+2zCHzxG07fOmmvVR2xr0Q4BYdImeK+1qpZ2v9mvLV/JMdnOugt
fzxRRsoMrdyQ5nP3lfLRflBTJG8nSNr/f5kFg4AAZVysXi4fNZR3kVYZpaIAxkJ3H91xkX54FaOG
kw82sLBLmKdFQE5WzQkCFBXAjqszb1jvD9/Y5kegaHRaA2fd3iHR2H5DvPU0K/RMmBAl3SAofcX8
wJpKYgRrji+IuCFtgSykQQ3D6PVWnWcKFhlWwmg95XKsJeMgW4N/fagUTnc64FnuC6R3gFAU4J2+
lIjNrFb18/ZIZpdFAH5LyJaOiYnbr7aIgltekuG80ym1kYJ0cxy1D1JOAIyvuhL+RfOpDO2r3z80
wTjG8cOCFI4HgWZ4EIKoQjLpMTj6vdubyHaoadNjPl9FzO4lp/MOTZJJLted4IhG9+QE8aHXVFBZ
3hSaNGR4clf3fXKN49SwdvhEcO/5bFvjOEBeXJwbZaFLCca7q5FNGW+QzfF8LSEdm7jbhticbXNB
h1pIZyyky2XqL16cOnKEpiWbRUAqwt69AEJoC01ZqCfkJdeIXDGcg2Zcia6PPmBj+Crf9xEeNfha
K1UsrV8KSaXuksUf8yLxY3/dZlv7IMtoMXjUwzej5eadl1LblGEfm2h/+ZE81En/4jQ3uUnLs2Z+
AH6UPPA/V0/brS+mVewnx2Um8nAXxpFoK51yarZmIOKj2ew440lYp49VlHVkeJuwk5D1KhS3ylYw
wwO7pVTBff3r2qsHOWGjjCsGL80iSd0iqfS2hjxZDg+/F/DnqEilDqWThDvMK0HaAFG/g+mR2rMX
26gPkT9zVfywTgckSt3p/wUzNTFNn6rTj3tyg7j+fl95IMErMsp2foWVi3BxM2MSGzZOCOwXKAkX
LaXsingQU69Gjz+8t0O6kK2sUWRO2W2W+UxYRKUveaRFs1dVhEbBbxS8JUXNzlIA5glvGzmrHgJn
2RbMWDJEGpMsgrv0sxqDJ9h43IvBnDqr4K5SFAo4sTZzofmn6QZ4W0P5YHpH4fD8IkzAXeQaAcby
SOrrz55hGix7bwxPutBaO3sBb3KGKO2lr+PmzmvTLr6YwrSaqGiwaaULoMudr57iNibv5dx476wk
pgXONKJrt4mKonV9jbYl/lCK2cPOBaAaFn8do/XFCsBN/SDNF8WGfIATqUkN3cm9y2aUZHElIJcK
u4KiQ+NxLY5Z2Q16kAXuotIKEOCj9Xz6u3yTOMA3TalDGMB2kXPh/xlrD1WrYfFW176knFu08EyD
Bln9KzVcp3oK8GNzvCon9V0zjOXkJvFV5PJRPBm1ET3eK9XesSvlQnlTKKqm+F3eiRHB8l7mjRpv
3kyWGMPtnX2qMpEg1GfvAthIduIvcwhZc86qRINJldXh+8/7FZs1/f4qyNiWWYeTCn5PW7+kYuwp
l/zlVuBqXcUToED9NUkHpUEzzZbWpKEnVdVJKHw6X18tuNDqDCJhfPQrZawCRR4xpvN2vKyuqrAb
b3RvPdmhdQt03x3kpfQeHNn+9yXjsgNX57eyUnc4pnbF52oD66o5P+bBCXYZujeFtlUmxg+KxycL
Gd8zqAbumqhFvC1kUMJZ9x2Qr/qrbNpMUdmnVjO3L4DDGtfa46P05DzGWR6QQaPhR86yg5bFO6xN
qUjM7CSPPN0PzuWz2K9JHWfqOWHuu04PdaBj9WKfq/giZfYgd5YagNH6xdaMjwqJZWSrveA32G0v
0ZcgJYi+wPDk50WmRGj01oAJd/KneBLuHI2h5qwSEIhZbDypQAf5SU7QIRH068ByZOD1rG8aprdo
FSmw5T0us4ORInNk0lMfZ2yzPubCFGC1PRe7jsjdf8IvZerMFmFovzLjSXue1A92+FrG9dr7rPNq
7scmfMQr2yHuePvN//pfN/QVrbx7zansDcM4RBPN8thSlvcswdScNWrsuR3Ri9NAuh0zskvRAaG8
6nINbD0a7Al0gi9O7c1lFcga6+u1WHvErwe4+iTSdKytEGlm/sgX6qikRm7uNt9fUaNn/OG/nFSF
l1OtS4dQ4RHcGNVlxcmp1WCM7Vz8CXlpr9oVgi41hxE18ASjTei8peq7YFxc5xKmUxeaM665OdXA
JzjQCJ57uAMjul3MLwE8LEbLvPIgrlMCOGBTF2OkN5AgAGpncyV0RxIaIkIZhHM2pGyDfuaMsp+l
djsHo30+Cw9RcoaFRs+LusxK8eG7O8fnvjUNz3ZhfEpsdPFrTeKTS4rRkZlg1YP92uOUo2bZNg+c
SIUJrEJh5JWfJDSjnW7pRrAUGrotMYVOLwOvhOPdNN8qDCNI+lZtS3u3uWJNk8DQDKTXVxVHoYNl
2qt/QXgn0MUOWR4zuOSZG6IDtD6o589GNlOJTeVqIXzrkXCaCIp3QcIxUHQugPxY2TXhoDkbXfbi
i4yeairfwEhnemHbRWky8yNWMRBGuZOtnJQNK0pYMyCt8quLhyxV9Ro8BMYQOgdbCO8CDZqSi5+q
bfO0pqp+QxOVjoqCwWB2jPm391MdpgwNXolBsnOwlq2/dEOlcRlcYgJh9mypdkHeh0j0dL9BT7HE
O9NR8XaRjJ/iqBYL7ukFAO6Epu7KenS9rat+hqzKEuGPcMky0MRCa8v4lxLNc+IVnnXD/9Q//+uG
+vpVDlOYU/0I02ZuwOrylY64o4TFKZUY0egGx67qD6h/HtjUosIjYKfhcQGI8txfY3m21KAX1hy5
hSFvaeBh3yVt+2Lzs/gI7CpX6p3YHFkvJ5ns7mQxp/gn3hXu2oIwtLUgGNQOjXZ1q3aEAxOilX9L
SeW+tNUbHrITibUa2ZFEaY6WrTewcqzq9/x4A1xoqe7q5ZwwRmOKpdAc6CfKpmWqVRjp+Xc2bPOs
Y84t/ioCxW8kBeju/vGeJ29h53lRQmZL1ti9R9rRvwOurv53wVmpqoxw19IqwkJkTNroqJ6wkcyz
6ZY/lYNdlH9BtbebEiundiiKnRJTY4dViBxgT9XEYUMRKYbXBSDziJ5CMwA5dVSiOPd4n/rY3cZs
svPLRv7IXaG9bkDPX+nkrF1RwCWYfWYknlM3/o/h08LPQPxeazNVrUZ3r1UmD/SVc8ppM70XQJrl
JaO6k5xqX8fuZkKt+6nn4NWnJ3rRBpnnXHtmbnMxGGuyekAHituAolIRdP8DE6oA85XXza9ZFBra
o8dZOIJfInA2Pl3fEC3yvbOPUmjG3gRJG/IPaGihJdytBCMfYrogTnVRtIYeYUlCJhFFpR/B/kj8
ckxHHrKe4nWGSEwb3OQDqqi3QqJsSAZ2lyOpTzeMhm+qieK0jBa4Z5GBvkzAip2oxYCEyjwMsvJB
jh9rUun+W9nKKSQRIFDyUEwCNOWCV0GoeSXm5EIUFYvuqFEqeSXKf4+LQ2iXTfA9RNG5/gvNMcbs
PWCzejyhLKiPP5s07qn1R96XSFv5A86nlNKDW8eYWA42I74av8u2+dcE7ocFzq1dddE8lFWB7UzZ
+t9/skHW5yJRRPxq/K08lhIpUsLic5g8YDt0FTD9uPRnCRTZoxpx2e1JtdbAiAlhAU+3/fY5XIOE
QKwQwXh5PP6BUmATYCFLQZJnn76qtYcy64F5sLqu0vUlGZUpaiBCpikVGbKNMJqSRpf4v3vTCRZS
SfeGyK1cz3r4caxIDsiWfqrpDspUPMMhV7kAU3D9jJiu2pgTl4vyFKAdu8kDbBN9JNw57YFnFMr8
wkBZAO/7b8dnK1OUUU5EeXItRyMCe3GHu5a9kdFdzDVvTVBhRIMGMPkpE5timrezzpBLTZfKD3Hg
xdLXf3q2pl0IMnbtOV4jZwI1k1r+qt5naYKbjl//yBxz/5Wf/KUZlVFm5XswbmznRPbxZvtUb2XP
PEssHa7JPDoz9GkOYm7D4sYKXnvJIUMOPd+5c2zKwEKb5jrFwZkelQfwl82kSrn6Mc9CakO0iumG
yBc6bh0uOrWrbuk9B9yUwxM7aK380Crp4oEwou991W6yAD8/4YOZiPhKrrv2hmUQ5YOQ8LxE/PEp
lgoDmOcuQXl+IID4qMf71GkmqArmWOj88JzeKeruwOVI/4XS/bJATX5nbwB5YAE9SH9MWept7RpB
MiGOzIW53b7rIN1wSvqK7vl658pQAGOOBn5pk1Atk+gLlyW6HmksUNJsobTlwP7Av68hz08qX3aO
WXQU70Mtq/gv1wEG4mlu+NvMIsE+lBhap6UVTNAL5jZ6tVKsQupaJ+sNavaiPbrWmtIuQiBv2hOW
rqgDCwKrK0A/CdxjRpqsUCTPlAZi5EpKiPc4L1SdqzxHkprTFOUFxlJ9UcDaRluLs7CSjjZwTB++
eihS72fAIDpZVYa/xQmfVFkq1QNAD9ul9IPmyeswcHf7pamqLuiX4UTbaAkpnxVvZnCIvGw6ZiAs
JvC4nbHOK+XYHRFgi7byzNX3EshPQAlTK/V+x+9mDGxcimqlwby+tLy98tNcAN6AsX+f1UXfMRsc
ucYciwz8I1c+52EHu0EXBGENMBxFE8EMVEh8KAP8Zs01e9lfPrMyFQE7Xm7nZOiadgFODiZFWBdn
EmCPJOZjQhpnNWIRv7XkbHvhVRC9dli90NZ3T2yzv6QcxtI/FXO5YwkixHKAqlvb+UQ2VSLncCPS
hxIT9kq9gGbuUYfQy/HiOOuz6u72yABExVHD5ZE0lg43QEGHLuvJystavtculFJDVtzuIaEzmdbI
fq9yXRCk4ijLa03zic6S2qjOlfRKvdjI9EA/19qAYEX3U7WClL8xEU4K61PkTf+PT0JJuugNBZqD
bq2kphmoQYWdjaZIciZ6eFQai+TV4xUREmC8EycqViCDxgvDCH1KN17klFKsAMB042QgOd2IAvTg
v1+27/QvDinXfoYpwN/B6PdyyvJxogaksr6YwVV4FcT/pzcRTPdaYp4OVol+YsAQJDnPDkapSfXu
n6JkyarHYtPJVKbxUHzCQx/CxC/j8Exfsrv+6BlzaZ+9wKy+fB+/tODzszcsILbdTMKCBdx0DZA+
hSKKuHzvZkJKj5y3QWMv09vUGIUtDaP1mja7nebAIwHVdvNT/XPHccPuDavruxaQFkzZ665uCIF4
cYvxIDDfL9mhtyZaceHGjiUg2f+7uaF9bhte6exDCKI4Z/TYtA70qGbcPGCbrSCmAkp5rWxOrN4r
/RgNCmcJKUN2BSoLTUMUIsE+sKpTMu1J/rZ8e5YohJxhgK37NF51euVnrqrFFzJJVRhiqegzfEEC
wkr0QND+sVbyy17ZKtRzUR8js6MPq+RbXgSnpbd/BrNash1CplXGIASWX/4Yz/AQIWvwtrH/5n9I
vrpIsIbq8lhk0nP/wVxeYP8UEoVkONMb4blT6I3QYYWAPuN3gKBXARjtZAeHhvwgnqqFNYSOstRg
QmzSD+Xgbv3TU9xNNcFq8WMq/5TuUpJtl7HlDS1PYm5hApf/W8FLWBwuLdnc6LdeXACS/XaN43aZ
8Jynh6/MxlBMC0auF+S+L9fRhlcIri1JGYhMd6ykctgP6BEkt2b2LYYjpJXiFbgqU4QfWcudp5Kh
OtLK5SY4UFpqx5TvzZ7VhCRsM10hMD7qCH+PtfdQtCEwsfW2YXdKuumfNWa9v5wi2b9fgzunOcsm
RhvHtw2YuQGVm7wXNjYam8rtCQD/K7MJk0tFyyMZgKLd+Pm+jUt/j+KqMYSkey4CMQ/Q6pff8NyU
0TedpGVEv2CjL3odb5trz3JV7a76S6CzZ/Ek9sD1WYC8gwkVVSn29hd3OhZj+EWdWQIJ8+MU6ida
GC0gx30QK6QD5bSjt9uanBACiYCXzJW5NLKY2JbNDappMpafWORhTJB5Yd2CI0toExs6CJJb5YvR
hTS6b6tDgK2Pn6p9gTDVW3bCUTdVHwKwxj1A3o/VIpRdZF7BeW0hgh4uqLG1NF8NUU2DaY1cBq+9
GeZQ3h7vEhD+U4fSZdEELA68G8LsEWcbHg58HsnsXhNstNH8hop5liuNgs0xUkNQ6VsdY8aDwB0Z
AdgNla4sag8CfbStjXWUliLEjoCEyJSER3VsGNwaaKggR0lUzr36j6B3k6k/F21ifkMvYuC6VYqc
5apdbUDzbPFDicR6hj6F/08ePVId6wQoscFEKKF7SwjVG5qAeShLz2wP2xHcVRJ3XrXhQJsvlmVz
60vB3TDAv9mqpNrgLY6YT/9QUO90aUraHKGKenhLU+V+L22jc6omj+VA0vJwoMFG/lQW2hxDv8sc
DtQPkD9yeF6fkC7d4d/OkPOJM1BpbMvpagLYsfMQgOk3ESEHQ/vVIjdx3vww03GVwhaiVYpycoEK
Or6vz9jAgDfl2RYcrmllslALRTWA8veLkHRFasVDeIGoBdRx1T4BuxgV0dv9GO9Tnu3ymBqr58OU
1IPkz2eQsmYmf9y0dZJoEefUv1t3DA5cSgNY5Xq0zgx4i3Hws3ZagY2Qwu1JiEZVphJPmOpWsCNI
SH5Teu+f9jGNv/2FY2wSYltrdHML0Le+NXG6h6xsS9f2k485D3rBoU1VLxpZa8xhgPesBkKz4FDQ
Y7Iadx2+SKKjtPaVpOwIt/ZZaTbkkAGiy9uuwbyV3ZEyP0gftXa5xcajpbne06R1WMWN5q2OMMye
fIgv31G8hotr0FNg8pFc5IKFMNjY8LTFqNglKR7ArG3c8Af8qNtaWFjiLtLehAhvVoNjUpvh2c76
RgJ55f9eYjgO+b79KswAgYpZubaaWMOlunTOqQTxN2VExYDJh0Ke5PHkxoiXOHjJH6WM71X0qqMB
xlO50ylZ3Y2zqw7jK7hN3FBFglvsFfyFXbquSagPSbCywZKX6qe60wgwMC8eX7DFTxt0wc3afJ7/
8vC5DTPFw1Nh0NEWRShBPZg5Y3Hb3Oksw2TmnaLd/1JgxZ7VOn5F6FIP8hhxuqJqKEZGjre2lV6/
9HwU7oTwNkmk6qsVAotEP4nfndBHNzagYgC8iMo3v6QQHXMLUEwuBKaDG+Givo42qHzKaafNRF9E
/5F/UbNmQgin49pf4TZMrbJwZlFvCrupNKpUog/GZxIgDR4VzxEzlYYDKkk0KP/JlR9OpUPwZJbj
pwbuoyIUmrdP5DxFd3sz11t6r+jn/ZOwc9aZVZMV8T8qXy5YKJgIHnv4eGhkUDq7J4C7TaJsjsru
ODD7LcG8Ga+hven5Zylu97iiWOP36X3FoT1Ckl/zyevYutyPq6RhP8giS6kwTDTJmOThhd7eNvxz
v+xLk27iviMDmhJhjYtxe81v/ivJ/l6u8Gu01KTSENf0I7saOWKcO7OHxzB/bA920iWXIX+c+f9k
IkDBJyHST6ElZO72nKk/91K1OfEl7GYMs6qSzD60edhy/EqbREuqQWEXX31T1hhmnDqnN3rw94n3
8kLHCUsw6tJEXQFIC0P26uWyBhiKUAR2/EtOELvymYek8hPPun1faGc+VTrDdhRyLFm+mUfxCHhj
0oOR27EuR4jLvMV2HLIzC+/zIY9XPz0Mtyt5FduuCRL7BmyAzd89/1PCZyreBgbd6Cn1i5jxiIQ+
za8QmCEAg1FRQc2QPBRgMaRfEAYwGPH4nHifQAxKhBgRy+nqUlch4oLtec98YygMMK3msuSNmycm
nBII3niLFeF9kY0tir03QOuJO+MsbGxC/uDGfIdAVNK8W644tOm03/MGP825k7xIo19M1Qthov+C
CcDNkNyAcbgWqFuQfgo6OL4ayHiGkjI1YrMYeoovr58i1KdKevxjpfPuGD8cx1q2tpeE4Qzr1rQr
A1IRKsT/WSUJcJ160rnc9uofb03ZSgzcaFQUuhdDi9zQQ7oQc8Ohj+KtsiFmINlkvATd+FjUDahE
U46EKmF93Yel2QWvSfDm/QyFt0SDFvwLinrx44RWWPG/+UIHohzkHe69kJsnS2bHElBP2d74c+Tl
EdEZsandrc7QZscFLMYi5jxeT6fEMMk7tIvjR5UmXrqn68ZbvXSIVgRA722V4dX6jjZ9sU8CT5US
u/TKmBG0tbl+YOACokTmLf8BOaSEs6aBobR/qd8xR2Sc4UVUgt8O3dMaqqhQyPoZQVTOHgCkj/Cp
N0eYLWsJixJbHzgMqMwvBC3KYvst9Fjd+Q1lv4hlRdgmxS9kCyDoC3jGsRsgGhgvC1H4RcxjfKUE
X2sKcRKTYy2g/VJk6v18z0Je0PPWzBrG9RlLv4Edg6GwhCViclzFSevyFS59TzRg0mkRwByFK6i9
QXqCOD8CU3DDqYFDxtX5y1ha+PAAjo3TzSQp4X08a1Lecyz+CBKkIwtaLIc+DCWgk6ILLVnMi23X
GzQqequ+1RwZNV7DJMGlM36yf1VRDDytMq4c6s7xZE2l7kcAQ4wWkrnRkrjbQxGdsd/gB/SpAumm
yilRsqYF6pF3vVpi6qmqbT/s373BZyNazSqZqaZooq/uo8muXLn1F2BAGANl8mTA0BYS0DH+zIe1
ERXKf5Sas5lyI2DGtFMq5511ck890vyX10SEw+RsCikoERduC8LbRwIBTHkYSOJNXPepD8cjuA6G
lhVuZCU/pD3bzCHbS7KkrBJVeEEGeqMw4r0KVjFGvyQlFXPLxY3nJ+XC1CT6ipKWiRcIGxK0Cbgu
dCr22A3aYihzw6h2WQjkFsfusSJlzn73MN9S3PXpmJCdwO/71khj2GUuvUxDeURIf6WKuNnJLHtd
Qrn0Zuub3Izi8gxmBA61EXcItfda0D8Fhtre9rYq3mR8rpU41GvQojxjh0T2jfhHw77SIkPRum/C
ObADMm2oMFomhEonmOehHQR5VSQ+LtQWx/v2W5uh2nyZDpwYhY2uLYuQ3KcPlGaFlKqiO01o7X5t
VWJqtWiMuh3ily3cDkEAYFgmwjsMShY8icMhxiokshJkTMIOLqnLSDVZmxQvk9IPkpAGbyF0PPLU
Ubtq6dSpQOvgYKEV5YdSteis6GfXj3+VI/SgjI86VOwf8mBK5SIVmYRJRTrjlsjZqCeaQm3JigKw
8tDK6L3AkIgok+40MUmvGZiJ83hm/RyPu4qxcc/vXxVrpQpHpiGCT32vVDZYq7+UcDdLrIAJi8HQ
nIKuNRdVbifMWYj9vlKNUPYFPkAy9/op4+XfEdkZuU+xi1n6hdJOnnsaPGV9Q6NqVfGaSsOT9eSR
FA4tC5Ys59sJdKsMv1UMbJqG7XWH131Tm2hNKh86NUFq+OOpGKnQpSxgHB2v4AAV/CvLofzaS5Mj
vNa1b9vG35pbVUBZQkD+neyB/UVW/ysv+jRNloNout4aA40A4hRvMngj93tMOan2DtIKcc4IzTUG
+vO1L74lpNI9mtXCNzTzlv1iLukZwFvaBdHepE5UqlYPNCZI5XOLq3KzHs/ju9nAbr4Uw8zZLXNZ
11JsJ+B26ixox1u+FN45DJewOiMBoSscmUo3IoN7WhjJpo1vZqz90omF2SPzWB8GSUcv6dg1peV4
jK8jgylt7YKAiIzlRFvLGSz8Gxd0K5z8hk/YnJahyHuWgOCmH0msyMwwiX2XZnpvOotxIETKxhs2
V3OFOCFoz5pT3JiUMribOMpTJLDl7cI83/chrEBDsrgaSkR5IVi+jbpsPLpf7BhhsqTXK/bDDnHM
Jo1OphBiQg/CyQFdTFRuohLmuNsFmOtVtmNcKW97wJFbM92szPRJk7STTkGH5sfKi8MuuLT4j/a6
W4QjBioBwYbMejfpmF9yvFNT2wLrn1DPM+ATvNlZicXb3SYopic2fBvT+5k4Znpiy3KPJtc+yBMI
6T2jYsZuMrlcZ7u/1U5OcHhwi/64VORguJLUy9oOJSFp96rf7UdbI1GD7K8AWbPE9O4znnc2Ld08
0HkZ4vlxTjkC/cBDZgUGhBEQvtZ11erjuMEnnrEsxxsvf3xl17EnQgpnWCCpxH5J+qQW32rXuHXn
c5mz5VfSXufvca0z9WSPCbCmXkf9Y1ceFgVKqcQ8mRXLDInou7wbeH+CfLbZokT0RiX8FUlocYay
QOJHqC7dz7LhfCsGUDAXncG88mBmFxiO2BBJKcGquTkEuwaIw7hMoBJ8b/FV1kNHHVGo3Sv/f3KO
wJyZYI3NNxSI7RP9mRdMZKYUzq959w/G+drn3uEcYdFFJNYC/nGyMsFotmiZwt5ScB0S1z62AGIN
SRq9MPgnN3QlzXKXiTpwttti45pbJZgUc5W31k/dJcIW5vmnbUrKr74jLjK7Q6PZGMRUofwz1+e7
ntdYWjnj8uAxtuLnUYBkyYG/mr7T87gd8XLiOeKK5NGqMNfJ5qEsctULzOV8Bs+aJPxPxpPyz7cg
l5uxHxLyGamtWQLXgpCi4WHzLqQdXk2BDEpB5mEXn7M649MTxhSJog4ynfyqrU5IZLnS5PvQ2rPv
uf85/YAa6/B1Lx1LidrDfi86BeHhkWwKGbJsPMhEcDoluhmGBqxCQITAYNuNRFYub34dRbSMdJQt
Vs+3cEDAsf4wQLqsG3287YqE28DmF+d9tbj6kG1nZ8Th5m9Qzx4nU2CcZ367RHN4QVKtGK4yMrHq
pCmSKeJ3VIPOduuxS4rBqU3uPanw1zCN551pnS4aqsfHMdKgRWh1f1ZUveERb9t8HRI1xrjYA7rj
qz8XVDZ7/525r31bTAHg6HTb80CeH4vY/1RsXYajzOltbWXuWKS2tdHypFgBi4wziIrSZyB6Bnuz
S0COvv5L3vJxDlm4jaib24tVapNq4ol+QMv3STwm5NdqJ/uSpLO75+Q896K0cixBaioIQ8OgI3oY
DReAlD7zYzndbIiC4y4WntI1KDFCm2Xu9BqRf3UAkvGwNNrI7lpa1VGc9RfkAcQDO2syolbAHFz7
LiVUaPulvXXAWzPX1HWuDo29DBbiJDU1n/K4Juagc+ASb6uNF/XOLGGKsmxC0rzWgleh+fx2q9sR
6ErRQk8oNHNEJ08dHsrYnpi+48rlXbDYza+/luBoEYe5nVqPbr+MecXUbIjiUpmUzj9P/c37aLa0
fLk3RUtfM4QyKdtMP6rTsNxqGAr79AMAVMx6UKwNHdMThdprJKKeF1HUFlysL2eU6kzXBOF74Pk/
Vuo5nDDEMfovuLUDgxZZyJwXj45tPp0Ral4YhK5nqffRS6gRD49qekVat6GQbjh4muQby25wOabO
iA4pjwBsd0ItHfoiO6g/CQ3J0kgEm4pm0LJuqytpG5FuyvEuppiWACDKai+dVQwX4qxhj24HqNod
zeM+CIba394uGwQZ+lJxFr27FI04gyhqxVi8npGJbQZhHU87VG38Jvd2RaTIDlnCxgW3Rzj/N0zT
vucQJNNTmw0Gh8qxHX3W9IlJ+LhgaQ2kcf5M2ieQVtUtC5t32xGE/adPk0m83U70KvOPSUG9rzzb
2M1KNz8ASEkUegBDht4xYnTuDFQlb4xdZND2S5jPtfvdeU+cye9PsXK8wI8Wug1pgfm0VDYQFSZc
oXFXv996+ETgQU+1P4UsszbWPLq5J/5L1ffdK0vOygwrHJZj+uXz7ioWJfFz6ZwKIBVb0f7PbEKw
Yp5tb9zy+YuGZWnnT4tOUZFozIr/gDNH/crAwVZmKXaCndiaxSh8ZH/mSPvrcidFdgDQC6iompMp
QJ9f471n0RSQ6MDhpWtS2KPfMrPnG3mYdZDF7raar0i7naquJRkED6+WthK0CFWCeJeUFqxSBbUI
TKLU14phVVhprEDPb0pEpn3g2NBKdJOLWLjM7p5havnOO+4bYmf1QXqIszw7tBelEDY/iXaZnaYa
NFkknHG68MiWjI3rld+Lisgu6dW+A0YNLjFPiDb0xDhOQMedkn9KygcJRKAlYbs7QLcvAF+v1XrW
8SadMECMSIPFHY6axB9x5Fbdh4mD1xPPuWY7N7vkWxWkJwZDh1Ss14ZOt29tHaOeeBAcozFbxz2d
7JbGl0oFuNiZB5Spz06ZLU6W7TwwA3pTZXERq9b2Mnt9UWV5turfMV0QKf/oXstt1bgx2MW9kPQM
O40tDQdottgQ0N3AZ7/cWlzKEkWnhpPKiazeaB0BenUTc9Pu/oDRez0g/Pj0YlGy4941eyK/Csn/
FcpwKsOxexFJHRGfpnu4y0V0N4zVVQVIG2dZZ8Pp+gzzwbfij1Vr0KMtwKUAxKxAUCM8fBXbYCYg
KGTq1F/ngTrBjHHHF4h4chj9dgeejdrQLnJwDs4x8HlFW0Hp20pQ8riIXe7o2Noe4/OOFN+uauEv
sIwpgOtvb8HhLDmFoOcSC+niU97HGvlJ5M1roDbzq9YXkInvD2moIvYEa01BY+mZDb4qhNGeRzy1
rSK7pdXyjCW7s8a9olLaXKmX18VMq6fLKGyyPUJ9K3FJRNK3R9sUwai0pK6xYMlJxPG3LAp/q+B3
ls8Dxa+WuHFxqZ4Vkc278u/sQ7GxHyogXx+JS8YjXDF/k2k9ENM3FGrK8i4KEmfAxLCRu9c0/pl5
akfY0XJukGZIqX76TjngZC8HEjC+RtdcY+h1gaxFooN+wBwBLhX5Q82E/ykLPNpRtwqEpscQnaMp
8m9wBxeO+tJP5xEC16yh7wACJgsKdhyiODrH5KEWDJ/sFq6DSscJJ2hfBekZ0cBC+xTtkkujpI60
DMXq+Or/NhLO24TfI/RaFhKLPTUr5MW97tDESUY+Js3Dn0SEq5uqYaTHxiTQ0RXvDQQLDNRD2MCY
Bxi33cXl+57475uRJbWZTUvmLJynl76AMSY29eBC33pSE/i6m8Nb+MZ1Q4Ap0ZCB1ec7uMmOlzGE
4KCwb1VGJMGVAn6/mJueMfjF/W1Azkf0e8WZ1Q2RwUct2ekOJRj+EmFmmAtbhd2BFosX6qIqLUNj
dbZ8H+3ETn1mwhMV77LKNJzzEXHHjxLPkO1XDepNH6bUL/sOhYArag5W8dgwMcZn+PjXmjF8Wf3B
qUTmU1qrploANA2O7wkq1Id7WOWcPqQwJCNdL7P2cSGjpskZEAwIIcpL4IN7tnIqI95QkSvK3J9w
1WLF0HwNKST5NAmJH84zZ37bR3mum1/KVZCCaFpT1B4f/Kc8EYhEpJh0s93F/MNySiAd/DT8Fj0e
IxndPTUJ8ji1xODqEGRpKOw3FkTZraNNw6YEGGFHWocx3xhXlGysXy/zsvL01tdxfqGF+qbTm5HU
5PdXhBKxuT29Hq+CpTDFuZ5SOOoxfxWfFN0vxvcGNRBGEc61EuW2vNpKFuwod1bfCb9JjyG1i5EN
r2LXueRIaxiQpZs2LZjTZJ68rFC2fCQpAoHGPyAZjtixMdWSf0/c9rloRwolhW3uCS4HW/xiDxjP
I+ijNctfWddyRWRDbbNDD1m2ZkuvDHNOfVzQtVCC48QnwkORkfsufK1hb6vYpY7orQ3xY/fIohyv
2wdyMPk/3OZN74+kU+AVwEKSO2WbzVbVhRgh4oT42/C4FPMATmHJq5jP1glbcd8H7rcZa0RqMY0u
PKWoxf+A1UbjXzJK8sBAYU3j6eDIuVEnOpqvzDQB+NC3tNKgw3PInzptzoJoRM57OYcLSVsmoj8G
4RAqkr54CwAxvbrS/WluMrzuJUKOteiH/B3QrlBIyKOKCHnumrTw97oe78g69MBRDJPWRN+CsikT
6aw/e8qz7JiwTajjKXatTinQWDivPD8BqXCuhi+RUISFyakGGjfHqxiLC55gDUhfKj3gOO3W/iGA
b6AhwE3HFelm0o57k8mjzBAH1PEwi1q+gm4zl6X5NsuCpD2yApSlDnQluTA14q8gq/YG+U8s9yOX
BMytnPCaLKvM4SYxK4jWv28apeHCH8CMtJLs3I57tIyeiiYChZqqswDkyrukV2S+k+wqTfVWptLq
YkmdCiEEku6DICvGTzvLFPhREHo2bvFau0g4vjzNnCPLQYJ0Zfu4WYUFoVxDe/8PcAuLzHm7AIeg
bzsCEpx9ihMCUFybwax9XYgHSe0FBYvg7dHx8eYfNzjR9Lrm13CEAS2sS2k9Pn68obPiOZ5Ed/Dh
pOvnokgrhXi/nSj/6vD+Ul2diJJCQWDWngWEfUpKgbcBtB0xQ1DHgnzLHZQZisA2e5karXD4bdoM
uCCYqNRLAM74K6mJW+sV3m8wjZZKIDgCC6KM2ttcc5FSY4T0skM+44h3CtilC3DtufgzL4AtjyVO
76XgJ7VqBUNHnC6XfZVzqBVREmiEUwMnvyQaYzN/y96NRSGcBxzPmwGu/g051we2c+Ws2RkWn2wm
jD24BDQDDMaiYOIKY1B5Eszt4/EVBOI79dtc98wvDT4muvTWSOZmZrybnHDonGJu6WgwFibcHbvU
nHsYDDXV6MZTv6EaqPcY+gFFfUmC0HuX4uQRsl6GRkJj3cDK2xVA+cv2xjvOWo6mtVFP4B2s8bZ5
OrtufUYyDEiZE8dns4ANHCzcG1aag2jOqJ0LzzkxyIwg1VFspVyK5IoNkUUt8LN+KhJJnmXCilLu
3X4vdxYNcxFA24QrX8dua31Wm/KBBK9B3Ou0kv4EFWKF6xVuYVrPa11WW208AFCp8vLGNfXyRt3i
Tqs85YosDwsP2CNBvxrR64kF7SoeQyY2RW7ARyTjy+wmldspOhGOobMGkjGuAgVa290kv37LJJEQ
iS2bjo15O6uJNj+18VnKbEr53PKCLEAwFm4p46jX5aiCVpSo79aSQ9Q2zoPEI8Y/nxRc5N4S7Fqo
UmerO+Fa2bhvbV3t4oLsQT4KfddyRedkTKxq5XxB7q6/rUhHhKU2D8C+YBqp18O+yvCULeYt1n/U
cxs/Bv/RxH3HEMxHO3Sfdu6FxUvAM/oQdvxkeVMZXj46wjtXgjk4JLCV2oNENdlla8iQdo1X2Qi/
OB/AGyqBPwq1fHoRZw7X5Cc0feupLBDG/mJxa7Ld2ahhqg5Q6sTOk7H0dI5JM3VGXizfx9C4vX6N
J33mfSAqJVHSZqtQRCBIrZr0DFXh7tXY/3JzSMLhDT54eL9rLgg8kmy6NplmUBipBnFqF/TRhmfM
dXUkUFjqPEPz4BVNgS4NWIW6NWhj9CTQHVtS1beig7jSBVRVC4BbZXwxsu04FqIpMMGVL0k9GE/e
Qk9FPgRDnrCWP0OYVPCpgycg7/Ais27g73a5CeJioE2dBjEkB8cTMQa6fihNPmJ6qnHAJBGdFfwh
urewtZa0NMnmiZ/iQXX72GtPLVB5ym01I+3YyuMJ1by++XFrRBI1+Iv5bRgo4j54rT9ugVtJEQyH
fMJ+2K45ibDANe/Tl28udohiaDddH+N6VBXXurxWJds9stgbdJWjynQWJjoUxSv2HPQ03BhDM5W0
zBzLkP/C7dRLaFxm44v8hUD3AZEuwek83pEzRimr9/fupCmEuLXn2dotTUqDYFLKzqXPYSrqLN7K
N6OJO6HwCQKe2pltK05ocgJPiemlvytPZj8tdHulX57sexIIsvXqc0mcXs+Hv+1ceVO9ymhSHCm5
Es0y94zwsPw3aGRyN1mDsjaUm0m7vaYK0LLsuXIg/++XP7jAURwLE/o3ppI2p59p5unzbxfofd5U
mS10GLQsHJkjrKVYxJFiqhihT2r2W2iUC62/z9YvB9vP6Ej7i/5QWiYVldmRud9xQYs8qo1YRgN5
9CDqnum+Pn2DkcE8k/nXuu9bVivTVgySgSKNNybKDPTWROd0wKbC1K5MzPWlQAO7NqLp6Lwdqf6N
FtNFm05onK3iBkhlp4vfMa1I47ZVK9WFb4ZuOh0bfDpPfNqkdBt1zdK+o9Xe/l+uqYDaIl+m7EP+
77zYJ9955r1zqoBuencqfFkrBSr6cgNwvHmx4tTI4Ql/yhlxWSuH5yDpJ1Sm87d9Yxsg+dUU2GmB
8jKFQUw96BQ20sHAdzbPLFRFMif4MEl8qAH5A2WebzWP9VJXz1YqXmziVPqRapVS8EIat2AXho5A
uI9Is3pmi1vqP1PSH7Y5U9GuUWVDFQzfGPFna+HQxaJuRE+gWdBsXVkPlvg9ntFb6XQbXxDR1OMJ
9Z83LWXOsSnP4CRTBIzoGMgBZrUu1izDyDc7bQ0u63tYFo5SQu6N1/75PTCH8sE8Ckua2v4LPLhh
rK8Dpc/a8W9YN8SR0qDaDv7qjFCNYtPLoo3s+I07oApTmtx0L8HH8gB5jDV/yrIy7CPW+UK3ONSq
bK3NbCPK72JtcEGEHqXBqKv9Ii8TM3TsH7aXOCP6CFxnVExkjOChB50f2vgNumMTzZw7vZlhKm+d
4+xJ6v8Z+w3MJ8U7mB75pFbp9er/Q/mH2Hz1wjzB3sS5fCV4//8iK8bVZ3V6q7+9jdt+Xqsx8hPm
CzrJpIGMYcW2125DmU4XmGDMTefLroCY6oivlzNCNahv/7PMP3Rs/fnjPCDtxrmgp2fY9MWM3tSL
dHQaQW0EP1nIjhXftPLAyH38tB1S+KYOBqdiG08f2KAdavF7dXFDOi+zWkZ6BR0YdrUuTKvQ55eT
tHS3DZJwRr/375RQorYYcBRFkPNGqdY84D5gJkvVn4YmGMod/hydncUlxkvoxUfFW+kmmLZPWddo
Cl9u6hsHFy63sv5bYhQXwmgJ7vkkcHHY/KVuPrOQW1xMj//c0pK+Aj3vwKI5zYVDy1lbFG0j//DZ
2XPp9AmRMxDGAQLZmYMqZbMusWRj3N/pXzcY5Ks4LdkK24Ndd5WREUBF3lEFX5JbnSV5zzpxTXYD
ftPG/20/6O2PMB7BG0Qo6LGY9FmF2NRzqpmycEGUwa5FQa7iHGCmeIushLYqGQRZnn9E1NHrIMYP
ZSwKPFbQewt9pLbIQ+SI2qSdgUayQKg1bIwcks1C5U4k92XPAJ744KDvmvC9RkNVB8vhuK3tB+1x
AiA/rULgDVDBQnICrFj0Q1erGvXCTzfJAAtd9lC+wPQeEB/CY25NQOuSSU43v6Fh6JkOSiwgLftf
knGthkt8v2rnDZeNNGZg1XZeM0GPr0uvod3NbQP9FnxidpsnXGMY/n6TWE7ewnfCGRClEggrbtDV
zyK+i9038D3UJafT7emELm/JNHv9MUdEyD5rs32fg6ISzGgVIV5fkVFXzV4AagkUOgc7S0zFk2DM
nkDrA0LySJhTem8r+MJOXd2LZ6VkHVDUd1dr4W9MxkgLnuQziCrbpa9Gi1dVDCZcESSav6Mvbbh1
DxKBOGvkxkLnoDAlcxAdMvdncw4/kNS6ZupjfVWZMrLA0cNSx6Is1eILfgmJBmWqiSprrUJn8epN
HKAOWNRCdMz96tS3hx0gdhypGZyr0I6ZHDQpjoI5Mm8CHQGFrmKeFLurX7qVWJVSxvalGZhUexFv
2prq6NbYAOxrQlH4iA1ut3l1r1qahfDdnQVpJfnvtY/1+fHLGMTPsEMuh8rMgHHkMapCmWxza+WH
mun4qrhQUWb58h1B0IHrWTQzncsLZ29uAogolSS9e7hu4OC6xf1RGfpZDe73UbmSbuWlFa0W91W/
C9hERRatJgxxehQgKcUNHydkpSwX8JS+v28kHvC4V2tklXgxjgeMEG7Qlt4x5hHqMc+6Z/+CrG10
P9I2Ju4tIr5IWHLfDe8Sp2UL0pVsgjj8JeI1XOYHnO6L5Udx/QN/LQB6IS2qdwu6UpoSKIa0Bm7s
EDOJ8rb/4bdWyOZhQW/PkxJS5exwflEfKs+C2Ltp2Gxgl4eID7GNoHrZGOHEj4ZzVWNtAxUWjByC
UXGkerqLaMVgbzhfbccYmMEyWJbGfVRytLfCI11Sa4rmO106lT23eMoiF8IV/giGpxbroX2NHHiu
Qr6qcuYGPtFlqvWBNeP+CPJ5q/JTKelQmFFTEzU8JhTqo+7vcqj7F1Gnka7IWDiDVrbXBoGEilBQ
1ELFtrIjZP+Sh/UIsvbI7WboVUVHW6il/dAz9M2PSyTkAy0Lhm9Wddk+rykJ/loQ5N2mR7X+jjkB
bW+oOBo035Mhl1kZWr4KEPCbe2SbTmnokMEfsm9IGlLTh9UCGDKpx0xVz+YaHfZDqWm/jO/jsew1
kdcDMcOIl2M3Pm/ETYcKXZPTOvNHIaLFG6/6o8Cb6OFrcBswdzdzVCV5L01JXlwprM4lY0EuGTax
NHeTUBmIomrvaIwVQFW5BXuxyBrXEtDb1qd0TDdAGSoQHY1Dhl71Ku8QHoLUByv7Z9OKXRknvxwf
G365xJDShc1X44RouBgi++Hp/D5z0oDAXGk5YNp0s5KLiNRd82y+dNVQgM4jI59DZtLFI47YHUbU
2tVERGH+E2STb3JSL5kGIiRWndJSGp/XpLyFko6FwbjrxVTQUWef7g12C+x/GynE0+HZRbjI50WP
pAP+A7pFIy57tiE9VS62tLIoVUWgJIQOVDkWkuXy0bB9hkQ8OmaC8ocTNwYVR57+PS6Vl+sjuO0h
XRAlzM3mE0eJP6MO9ZOqPlvcgV+1mqZ2I9V9jHN/yfLxfqzBkVuA4XeglHSFlM+ySARPP2ZcLubV
HDLr5qo9DzjY0/g3vBmbbru0Cs99/qpK0zC0n8WMTN1goTYopve27DvUrXXHu7TpKrtnAlOwGUYS
HVQZcFJsaIUscmfJUyH53jqMdKgqfCrHZ+D6YA5eXRPe36jrOE6IDa8SYjcoJkNfLxfnoEvufplk
HgSqeoh8Hi1RKKTv5G6Z2IMW3N6kqXon/g7m1cXD0LUpHghsG1mue7SXU9b6NFSPxFAKDRrHmCM3
+6UsZKLYM2F8QCxKozIA3LpFl8vwaC0aEiM0J4ec2b75vzVozLi13GB1pnEd3pbFgLuvmErA4NSl
SpXv7g2R4tvep6HwaNxksEq7LekQ6dbwRCCP7YfxnT7FFsxWcUtlqKtZROFm531lz5Jo3CGm7hUu
Asx4HPxg/M8nW7tWi/zXJZIQbhl3LXzS2zh71Ig4aOUYa7w77wdNv0OdT4QuisuuJbsGbpYHvqty
5IhAqom86mP4l8vEmVL1z44Gl/y9C/4Xc+E5sEMhKHvkZK7OwbQ9vo9T3ALZXYSdfe9q2JJ+Lg+3
vZvZvZj0CU5VbqPek9pqWOrSwOoEOsbe0jr71WguL0HyWr+oK8/VjMptgci/i7gH4/9KMK68Jdrs
vpRNdEZF6gLDSJTMrNgaf6FcuIp61Y2lRhp2GzjEfIdlzZKkXNI6Z/kzgbdwEwV+JiICJ1YV0crp
4PLUm8ST8nhe0hoxFGWndgfl6jDViuYwwLlXjzkPka5jXW1v2iXawV+rTIMUYsXfDQ+8h888nJgX
Knwqvl+BxRJNdGvMUP7Vqe6wRiiNKtMbd3ijkucnlDzBAzZF4mtFTBUsx0ueU0oQYYirtxbE1fFj
vAvwqztV3YLtsd95iSFDWM+rf43b6rGPC9uiWPbl8TIUc1RykhwRP/eZWgDwo9sYFuPY26NZiJGC
L9ozNMO/8vYogtqP7/b3qEvTlpnFw7owcOxlOHurnFuqzdUCL+WJamIfbDgwNIZFjGHhxV+/p1HY
jr/VLbCjrmUBXGoCBtnlYVJN4QNmJ1WxayZNDAxna+y6exhoR2dNHwFO8nbUCCggyjmFiVEx45tP
FMAW3oEBu57n19+AZip2QQBLqvTH3A0hUaihnRQe6AetJsbfxDxvWML+UfyKB9+Kr6ehETZoyh6Y
HCwHZWsHeucXcSqRK+Ciis0UMb48cd1Gw2BQEe7WoH3V+TGk4SCYyFludJTI0R/jMjw5U6upd8e5
4ADYj2S4xpNKP8rrkznN9UrjSfnmPLujq8YHwXFsRRCjJ71CeBqi9RCy318zbwLbnmkEg75ecHBw
xo7Z0Ff63e3YyHOQ8koJ02ZLWMm8qMADlWXCNIM7gWdoOBgFAITLMVqKXhLAZb4DG0QW+PvW4D52
Ys+ArB5FU0H3pVSNffWidLzI5ajYEPkUO2cIvNun/ESNOHL/7N5kNVFkAlwnWXPghDQG3jl+Aiis
xlkTNpBE9mYvGNU1AF+7xi9zV6MF4/BE7g2/VHUDrVuMBTV/qGbytnYGUnqjC+z4nfnd1ql2CQzW
FTnxgwtvCAXwNvIvVp7FhWUBBJVbLJmEkmsGAvUe2eyktVXTs1g/w/4VzEFmq+b9ma68fFozdPNp
/HNYRLv4nzL/AjoPYj2PxrZFyWHApXs4jsXcA17T0e4ivageHCHJOBHgqGowFiYD50vsLNnGVvFp
UUcZsTAmihC7XVQCY5S/a5dGrrbUMSVJNopV52PvfUiGpT8gSs2PFtmD8mxkCdsg8SgIb9M0BDU8
1ybC9eUQ/kFZ17jHAB6IkkzYhXxXtQl1lWnDKtfWhoKN4Dr1+xvwBFifdIK3P1YYJhT/GRi1L12D
YFo62/UYRr6IxaDUsxQ+fYOqS61vA/czHCrvAa9F/JVDs7XF3nrog+T6zSHcT/CiHk5Kmq4IVDMd
WhcaL05jaGQ7iiZIUNMfR8jA6b/r7bt5oUksRApl79Nl+AU5lzUaXGj/rJQDwlxXb2Ykox3D6034
6i5tL8S8Z4Ms1EEIv3X3K4aKifuy39ZSDD6oTBgbnLL7CdMwX9/T4aw3LqN1XP5Ujw5NSwI8ztwB
P1VouAT1g/gGa6iJBrGiqWVG6fhaoVSFP3csy+dIoaQNDdcVCosNYXMBkBazf7aUgPE+9sKXCNg3
Z2P4v7Qdmh0ht2eqVvdmiksXSWkWyWEmx0m27kxCpdDiWM1oojzgMNXgoDdDiKePhBe9XMZ2F+4G
fQicMg4BU65vOq0DQW21nbdp2y+mlArKC9jLN9JpCAW6Y0XEcLLTmBmo9GSy4hrdfinCk2fSH6Gg
mya+1tYgC8hCbk8mbvjpwhui8JA3WPhKScbry3om327VMQUCphUzWTdE2ZfP0kgxpOS5eopDIEii
+KBuU4UnU5dDoph7NmehZFueenqy3HmFT0tK/XELjhO5BkaSDy/mn69JM/PZiI0M9yfSOplJEuOB
T6PbezUsWb+Y99jF5xe5e5aQRgqyOaDnkJiFR9oFTjIbauGZmR+moAHYAr5LlIURClnU6dmC7L2h
DfZsD8x5oWEwio0BMDhxvd7bkOhgCMsW7PxrsMT6HBhlxAg83ujwR5mMw38jnRbO1CV+5sRU+O2U
URW17/qP+BknuiAzOoDW37eGemfJuuIbKU5zrN8RJbdWxrbirmGUzDyLQr5dOofr+8s59ujU0OZu
Py9rCI+QS4GYJ/O8ajfqexsfQpKyFdDp90ISkVsUuOWCsHl1brJdVrpVLnnNW/fV9e23Ii5sBp0b
DiPglyQMfA+bwVx5EUEEnN068ksdh0RB+R1SHs5cMkEdAUU7pmgKd+jk6AEG3yKgTBeGk+PO2Hoo
NKvpcexBPDIBKFmPFjPzqU3Gv4RdVfHJLDZSA5TwkIRfRPYVEBvwKiqjBWpSyjN4YwnzdiT1NgKj
jlrrn9gs0GqVQ5tp3mNelQaJEobD+r0/lN7lL0R5PX3wMmdHWusDZvpeTzpYR4DFhK5uI1ljiqqM
6ps59czDiTCKQTadfvG8KcEn5qnbPCBMGWXkusNXO7tPVcFc0iAQYeX4v+6KJ2Q+5J3PmZ4dGeaO
MBUDZq6ujE8N6cBbDD0pNvnG97/ajV0tF7xrrTCL2c5Z3WEPMf6rODjdiryvY6XKT3iu8PhLrvu3
suA/2hHv572TWnuW2ID7ZhFBV8QrLKejUsRD5SniT3zoJ1YhStv1BxlCRtRXkYGNzDmw9IyLbd6Y
5OGoBUYwemMVhidyCzzdPczC1n5kOl9CDAGnVDrwAOM5lRJhZIfntRi4N8bwjywXQLg4oLWnfjSq
FfyoYqt1PWesT649N/h/Jg5wJtjp51jD6o/SqiJ5HLQ2HcWon07Epikusx6Kvb5ZAGHb6nmIoRXh
gDLbMBHN/GGfAJwfQUlTp8bShi6DDfZfcl9IAitnNsblufRVSFy1cbOM3APCOD8BQHdkqYMp3qaU
Qi8LfgrXW/YakLbw/9yRVynnJOknvsMCsZPGmgsut7XFwmlekn69AILpVE4ALgWyR3LKqh51DfU9
snvOqwxILxTlD3OVysCpykR87RnnYgRv3MiQprIcnz7oMc/o126f1dTJsrkTpsq0IAGRTuo3U4+v
O8Ya9KdniAp/sXQlSXcZeb36HPTF3sH8kMNUQtGz+3ugN5bYf6QAkTsd9zQxmSnZlGeaOva9I1SI
zjSka6CFnND8dmlBaTEb8mq6CnS9DyUJYiPeZIlqAlnHjgVo0Xpo/TLLNd818jRuzGzmOMRy+FB2
gssHa3KE5Sbf9vkYrSz6+HSe1Amu0bar6iOVEvNzSWWdJjoY8PDpOf1v0oZCdlLnY2HUhyr8mRW2
vWcLxOjT016h0bZiHOO1ncShV4MTG1J5FraymGh49JYnx5XqL8nOyB+QNqEYGqWaoCNehYqjhAL8
Lvh2vwyLePE3xVlbDgZZXxeOKO0gcSGOKipN/CMz1H1yNGyu/bNDrMA1K+NUcZfWbgFY4VIGxtBl
dj6JOyPLKWwPjE+6K7KD7dWnApcsMIYmYUPTG5TLwCKFlVYoiWwkaceoSgiDtl5MsXd6SYSajvWo
2PqhLAq0lVd9MITHPncsP/81Do10sY0jXEvpY6x8CNnYirQbzGaan1mLr2mxnQTOHOl7ptiRMIch
fT+CwZ6jwUaedJhymxjUK0EE9kkbHdAuMw/6+LMYsk0jIv/unEr+jhlCJniR6eflf6P0HzW3q579
VWx5FroetTIwes80XAwzaJFWFG15TFIpzq21thD5cwjUfP5TxTwWCIZQLONkbti8Qn0TfpppgFIR
qEC5ke/UTH4+uwRhzDMQn/lIRhjfI+XrT2MD0Ch9NDkDG4F48g88Ib0qXp4OHHskKP/TQjyiA5p/
MTN0mpK77wW42jn0Hw8iPg09TlAEyDNZqF/o6nnzWNOuvXNmmF6aldxaLxAfzxZmxNbpRPbcZBaf
6TVf3/mx4w4TA00U6t1BVAA/QFjeoaVTktz96L2HxJWGKHZTLcSHE2FOk3IiXAmEN443+tgdIcH8
BkwGngZ+dQUfE0W/ov44m+SKhHjvbRIguFyaMl5Br8WnvwoD2rvuP7+w+vgm7hMcrUBEcrftJ6Wt
gacp8BW3oIQQKnpb59aTKr1TRWGCiE7u1mePKqZl2BC3/7M/aE0w/L2L8CZYphte3JaeRtqnjO0R
gwEEUrVMHFfqhh2bUlgzawlucWDcroOwr4ENPE3GmEOHejpjjzVh8VKxY7HgsSoHyRPZDyEnc9EI
j8oZVbFsJ6umu/h9F8s9qTgXf9KbgFhRokFl0Ee/824cb+TYRdngAkwnehwongDKYQhQn5aReECd
dm9uI/nlAGasviatKUwMMD4l9Gu6pqaT4gWnwoijNl30BSDcol4jf3t5mJS3NhI0VsTl3MRkGZol
Yj2FsZX4kVC3t70Je7JwvTZ6Oey3fkYIXHA++/fQ52xubLU0uXRi0n+S1nQv3s6T4cH79K+lr0ZB
5Q6Y8IMpkOoiSZkvkaIKN6OpYDSNK+OAzWv/BQ/DvQNIqpSa5A4m63ntHvoS08mta1jB7ZHvAmD4
znwoDnoDzhQvmIXhLKEL+tkFi6n2JAaz7Xf6Ed25iOp+Uh6MCr2Guw2BNWz20L50QsrL0EG+eliz
zB4k8XxRoUHrZExGe+pyvZMuyG/gfwEeNqlOHWZjbPKNPyouDl928pOHAJ0jaTALjNGKrDe4J140
udlDcfG3LEHIkh2Y/pad9wdldciqtSrRbjrKkvq5HRxs+ew0HEl16BnlDgBZT26/BcRM0AMOZNFY
615fuXOF4Faj0R6nuwudgtPSYzNaknHKwD0G09RBVdzu7aZiSwCiAJj+IbmJ+0Hr1wOmm+r8+3uo
pGzqaw8kWtMfRrHw7lB78C0tK+W0np+lx5Ku2d6s/W0r55eUmqOaoBVg+nnY1S8+1OA3/FGWp0fv
0RBiMTIX0moV98vEAjcz7qkGHBtH771c+KMxQy3p7sDJ557PE43Mhn/PUT6y2k7PnOUNh4T7p2r5
SY7XYBC3eW1CXJC79dfd2a8mIFP5jRbR/XZyGZf97MjV8yWfSXzDOmPrJS0FAd2n4CmIH/vu9jlE
1vLN2S0+uA5i3PdTnNrdhDeGPfPqVQE7eJkmEgc2jWfd0eJXxIPIVG64UtfDFlMNwIL83NJ5kv7F
KAZd81qKI665SCSWL5l+P+zP8h1GdUeLR/zMtGg5bJFB2ylNjjOMbRIJVPI8v01MeEWfdqe5O/cx
8MLP5VnJ3pxdvLAxqttcbs+VOWwtST79Raf0uH0V5EjCTd018FINhZJhOllf+KA33TrCXMkHFrQP
Nrp86/wby9Zwo82QIJCpQbSCaaHWIeJsRo5LcoNXwXkt+l/R4qNieNmSf4XSq4BOenbAXqWLFTVP
10urWw3e/t6TSIuEN6KauP5Ks2xGa3hyX4wYKl5horvYWml0BHW+DHobwhtk3P8SkyOI2IKGyJ47
L3JphB501L4jc1L8sRY8YRo7tSHd0gkaKZGkX4p1j4fzD1sGARjMiYWAp5Jz+APLi0FoZGrYJMvP
I45JSBHVYd5gvJZ06w4AQC1QjsopkW2Kn0Vol8ePU7gYnDDspTZWI0xMCfeUXhQ6YmOhsTh/MMBh
L4D9o4/vbZLqJrTjkP/70SG1Re8grp4104g0NUpb9mZZ1tP+WJT/Ki4GgW2laohKETqH0K6+F3WA
B3KNlJH6ZtLg5f6upbuMO2eOC086xJiaVuHPNjwmyRDmKJkqaQYBgUGD97YGXj32TfcR7zrAl+wW
rxnO36XZw3muxkVyfrTEem0zr/tllEjEZwmMrF9Q9g7dB3K4EeluFasd6V/n0GTbcZN6yFhn4okh
XvshaQx8rTgAsUWAunK6Ukz63Rv9xYY8IrdDpxfxQWdg3DYzoImMPpeAhH28wuiYJSX/uy/dmgOW
ahLjukO0QEFSmrFtKHIC7w4j3mwxXy3cRy9Mnn+zEMkecmdDnBLHNc/2sd/WSSE390/8vInVfviN
pACFSZQKQZ6P8UyuV8yPYpcz/ucblnngm0iYTFd9Peubq+qsvbyFRxVDYRjwYsTeostlOIFC3UJK
iI99ckAC0Ftq6OrTVrxJRuGF4CVWsCR5tEKgrmK+NPO7kqR9SZWNj1pNELCdUjicZT+RyOuWaRJr
jxZkjS9co5YD3lghxbx5ulSHo0G9Tqgw296jj4AiALqakrUooxWnXHIwi7pjo+KyBkEaMQuUhVPc
j6aZuxrLYV+waQZDtDSz26xUSRMoZHSfJYRc3LFvtgCj9ptgTZmcwmSBJnoZCA+hFm3YAUByyR2r
Ca976XaQqhfTIgxjKvyrlxG+9Ip6ZXzFByN1Cozg0hSVqrU8mawG45G784db3M79qtnWQ+Jo5B3E
7clpkBmwjrlDcRBRAc2UGiVmCOab/MewvKyn1578r0K7H2KamN610OEV58iF7xBBAEJp+9W7tAl0
s0dnSP3JPcthpuLHkhIHTWll58VlNMziph05lPeCPkrHZuVgP5hz3KLr7PKCPAVGtyPdTo9Oz6OY
OGYHdsV5MhdP/jwxd17bvG1n89DAGkqkQ6wW2jzzX97e/8vif+/KiUdYE1D7yhv6KHtnOx0uVAzp
dmoQt2lQmn6+S30cpJgwaiOkgDQ2oqG4qnAoiNyrTkBIoIHEdXV/5N6V6lAoD6zo6XmxIgmqA2kt
lrR6zBxz09T+SZhCUGaKhHo41H/O0A/5Fsp5p+FX6YYcIUYEdr7fKIQkNmDQDc98FhKYMNsVVKTH
20bMriE2HBryDWOXnYw1gJt8/GUhU6I5aQwVSk7gldczlcxOZz8pqth9KeQAjeJXQowQGhbZyIeu
+qLfr6J9OJElfViiEXXAxmGL0Px7C6gQIry3Kk3iXBCATIh2fKmbqWATSnl+PV/EV9UmMBpcILh+
aw0ePEX/UP7noxYskO8KV6AXAIETfsDWFn6Z8JdzAL8zgRybfyVEl+/fZh6K7E6XOr2TdQUm9IFa
OifXtVfoBuVXMNPwFUwFv5pdbf4z8NRqXXKEFpwXhSPUk13I13cgHFV+1GtUPFKaXR1mYL9aWHVP
SY1+6GgCIT6hRmCvRQ3oXAc2sZUuzQU/dEt+3v9SdODCIh3zMZ/zn6NpFzg993IQV9rSXlsQy0Ph
4BuXh9tzN1muXf84RAovyyPk+UKVYIpHP+z3DoKBt39bLhaBpi5nDO1HScgIkhZFbg4jLLsx+sNa
mS3dPOo+u/Z8XPfpI4PsNbNnJT/OfPVDLYLSnJkW3KfptK4ZeLlhD1s8laFk6m7sz3icYebPnC7p
zwBUxNDRyCcygKGqpV+AHVNdYr1dfJrohXOfLvjv6RYsj5GwMZ5AeIjxXoyEJ0oAFFmXBO5slVf+
oR3QmAXgeHh6fOEj62oIOgDWHvXsmkthHrRZalKcjZI/6wS2SF4SdB5I1YsnbEqgBhMmLcoydZaS
z/rZr5hUfwxb+xGhS2cOdx4qNBrHNhAt7Livyml2HxYd6snB3scotb+fHOC8OpZlR6CPDDJ4xLRf
nAKRPiwHifOtzSLtPHC3uMYWo5rdWjls3hwZqmfXFQRh8sCzG2tf9LD+rKO+HX3xteaf6XDFgrpb
oGE2VhuvhI+ZzzTUYhUvyDQXiWQY1XfZKGwhGuvHCFyo9/iShJ8xag8g/DjeUcn0h32G7brc9/LW
jKnL0PhfZgtAsmlphwFzeb04PqFo2XdVccm658YmHeSa5PHD/zVkbRDrPHzJnffrlqrmF5GM0P4H
xWSBeZBWtjHVGn23u87EarsT59ual8GFmGPtuZu3fxRuntwsh7mvF/RAl5C+p6wSAYMdw5FdI7Sm
DrMjxjNXJcGXDfke2/a91NOQvNjH1pUWHMiQV2StX4oilxrJK0zS3EBsQUCE2COrGfRVrOHTJRiB
fFl2Nxy5r2j9kQx4in0rd8khtmlsVqxVNgUGciMEbp54XLqXZ+1Xe/kfJUs8B6O1G6MteNtJ5pmZ
hwVKhwVRPLgiRAOulLbV5AAc8I8OmuOz3qz8wRw1qScR4m+U5idM9WcpoC0LM6ySSiWAIsvOrfKp
4W3xUibvT3Cbc/dAPGofMcZ5und1n7cKGavHshKsOGxu2pcUL0T7ESZ/hl0mb2V8I+Oj5JdfgS3X
mX3eDC2O0DUhviRtpT18Rk3TtGjfERI7Wc7DNYsx0OLRjNmjPs4F5oFnhsbAiNGfJmRIeJUD+SPT
AeDhoIAxi/KMgTSSYTsvyODr1YDMrNM3zMQ/2LvXDVgpqyizK38sBSpKUud+XphX+bkPCAkMy+hf
hOgysoqhyhkk4mVLiE9enTbwrC2jPE6WDybVGKN4LHU2B/lWUGedkRHtQWVqypxjRzDPTpXL60oX
QBlMJruUekW2XVTpB2prTJgkV1z0fbuwdPVkqrPkHGNery3BMO4SMZhhNqLKh3BtCRBbQIc4Oujm
eaVDWhUw/zEs0FL4yAFafch1Pzc1KEOX8SwoEMnAgNOUCxeun4W6ds4vzA+g1RIHOKNHGGlJGsQC
qSjC7hFKzS1S4pcXsYu7Azxk9tH7XZKzcafkXZDiejwJi3mgKkeQpNX0P4upg0d+S1KOWlA+rDWJ
BazOc+JJC6xzziXiFaOqMzyvbOeXZN0lwMHDb2P/iWsgLsOjInhNoDAEK6fJW2CVnCD88nITpfBh
1K1ZBbtTzpv8zeH0Pis6WHbvCA5Q4j/E9W3OodN+XbnWor3U9bwPRlewlePT9cYVQ4FHfjsgHZHf
hzqDu3xXGMCgvVhRkUPjAxTYtyxOiqY74PZ/+spDjlqugeWuj+Z47BNp8O7R13A6ADano1I1DuTQ
0l5ZYnX/znkwIoq+BcdShU+c6CZybbLb0W1aej/7xtGgHGI2qVt5gTZR0HJHU7tH2PmHv40IoCHb
AWiN10BOS3PjkPQyHnvmQ1NL78nVUX/gvUa+j7+lkVMqBu5EQzOVpIIJIX+WM32oZQlbQ+gO11tV
s/+452DVae/iBE6xlXJdLqU/IldARLf7A9aHcmsU9b83fmT0tZlQM9sTDDPujN5Zxkf9YnHtr39Y
hbL7yF3ILsEEBqtQrxQQO83uBXesPgBTFUfkbSpunwgW40vWrb08dTsN0vSvYRmsWQa9QnlQsWIZ
eKfqfx/AmMA2YpzDJkFCD3vVYmynWeIJv14G2tDOh4goBMjhSer7xIyXQSfrJo/kEP3riIc3URkw
6OhxmHNHPKZWoB/JmDbcGL/epdyxNNwhYA/NtAZDAqP0j90Jj0yLdcXylttt9rblbYPS759SEpL+
6OFuGsB7LpJpukEdTSGSTGXOb8zTsCfYVAk9MCOJxW0Ik8rZzPUGPZAMYouiuFAiumIVMNpsVZUB
HE8XQpUlO+gvtdPhvRuTQPtanHN03BbkzQdC4QhiakbGmLuZ54Jd7svLilaHymYi9NW4XjU0jUF+
EBGGTTrwIKSyxhQfU8u+rIcezG9rho6WjD1nuzeGgo8W2cG7NXgWW7lHzXK8jbEYt13b8RHw3KW8
WQfaotwXluHXGyKm34EhA3D9MjYQU9swPPIBlwtvaUj/mMlfhTkVOTEMhBku0Zm0TYN9k7pxNsgM
ZbAuO1lxRBydFdetCQsfxbl0d+xyzkDjuRPNzRNf68Rnn1ecrbg7NnZgQzYSUKT8AJjHaajBZZb/
OGJ6AbmmRWPou0rbPMFgUbHP1oZSqlInCw1hn/3jWxKAJwysxJfs5JDzdKK4EI0dSuqxF0snKUj0
d9KtmydA6YdFShYrMyg0fS/2oX+yWpNHj5YXWWZOI3K3Rbu0LZS9Am4Mjo6ZrFPXX1fF+EYoT5w5
BAi1LBNyZApAKRxsV7IOv6pDzfXB7EwJpwJWIy9feQp5kACJOAwnoTQvi3kjXhd2N1SRz/OjUbBZ
/C5+8Roj/THOIxx8k+nZYXq2p83wRsUr655RL6RC9WxhFSzyWuQTsgUgK+sRWWeBmH8A7Xvwgt9g
sfjMCNYUdaBVwJE1lljQr0jF7Qq+Z8B+s9XEuOKwy8bupygwMUa7sNszHex/WO7HPhgHoE6o08ze
Umkh0Yb2Zo4mbVhaA9WWry7ZCaoM0mih9b5aurfIVfEQ2Wp0Kc+t4EKxfS0B8TtAqwMMQA1MDnSK
CPTmyYqrBWWnmt21caTW3+hzxHRgo7BCBhHayEFEnScMpzFFhpGnUJsrVAWUn0fLBjN5DamAXSfq
DKY2h3L8zkOvIbq54+vTEibILfHglVlY7TXMMOxkCDL8eRdSXCjXaY89+3kSUYA2chaC4OYWjfSv
Mi3+m4qR5du+gYp7tE7HJXS/1UrihFDXtBVE1viafwISsyPpHVhgNYT8OUYlBMJIYCGSqXPIgkbh
RqFjfnd1hc20zpDrlKEvZ1/fdkhBp9/1A1gKLC2oOZ+kfaxBU/b36sK+ugzhuTEI9IrDMTmanLGc
bEQYitLnjSq5XpT0GpYoSQ6bLWOanC9k0e+SkzkN1zIXYYFoRjEUlqo7NiSvCHYCw3OUuTFUn2o2
YpMun4Si27N6kmthxyO2p8rwBJ2IXpsnMANqOwfiKTLK+Bw1mDuqEhxUd/hTceT1ftJ9KnLQxTmL
tIhTQgxtU9ZHNkff4iIMRMDROSvdERCC0OW1lIiiv6rRh2Fa0Xsk9w9I2zuMU3Rxm5tBCwDsyMEa
IVU6FPopBT2T1kqXZjWZJ2JerxU+X01JCtWzMspJJkK0nZbx+Ol70rucsQDm5LeQF5ha1mc+EgYj
Qhs9IkKwMMT1r5KYD8YjikdI7s65GvRNKfltnj6jfK0gWh3hch6amR/CWdmLy1Ps3XyDJz+cWUic
zmFNrJq7Jzsi1YBXKZ42aV0le3WErOYqFB9+U4UBiiVMvPsVGI+4KlM4nid7A+0L1HAAGwYV1oXN
o448dxhKj+o8T2bW34RuQaOMXPjERR/JW0vGVzR3QLJoX8X/6+g4zPGS2J9jLtbOKVIvZtozVOVc
biVDkCYYT04KdNxG9qM48/fR1cUBkwr1U51mvC9El4RPgN/hl6UG5E4SJUO/Nycj+9M5sk3xo6z9
o9Ys2u/JNtL5VqTedo+4sgc12oPYVkSHpaBjcpv/+xLvROh/wxrQXqbs3dJ1S232FqK2KZ1gJuv1
5+1gZ5C0hMEl2/5EHeuroEixcuhZ7KkU7GmPlczZeqKwVaoKOaBmbe7KklmaB+YHnj7z52WBXawl
umMTCvaS8Q/K414F/M1lKf2dQlDQ6kLpEDcqogBg50PtlnjQDdop4Cikmx/wgeFBVrMMS0IUv1v9
2Vf42Re6Lm+9y2SckTaPpv0OOpvs6GLG0vYgwe18oZJJxfDgA26sfl6569RAhCKbd+i5NMEOq9G+
hTuiuGOfq5yBw6gZLAuxi9VWkgI2+ni+7X0T1Cimawl7pXe7qOd27+I6j2eJgTGu/G+HISyI5n0X
L/oj8HMuU50W4LwX4oskNxpQTeYwcBxss9VW0AH3MAYwM8qI00nDF7ejsVgRZnmBNFvdssvt9csb
JV9RWojZuYyhZMWFNGRTC/v42P28+OU76M37W6Xt1FEG4cj8HfkCafyL0yApqw2/pXIHJVKCXu1+
zPhLZwNGx4In2GZYRqVpWigt0swj83/X/Y3morC84+YM3k774kFBUTRAN87wHbyUPNxJlWohEVbn
MsVOC09HFpU8ITZ2pqeKiD8B9ov4l0r49KyHqu2gMLywXbUdk1A7FSjlObBXOnvJ/kJxSnaLm4uw
KIcRrUMYIJlTunUWKZOzNHNSDI2Zwh+E/II11gBPtUC+eFzNRcupy4zQpZ4h/hFIK1jTtVaDWUEL
U6HD91oN36rtjKRqBTMZdTECVJRnPBZ7lJvF660WwYsSs7A5EvbgdGZ/XhEJXu4sMs/JfVMC9DT9
sId3oVyEZkH8/hMzy7H0UPx9tJUcHVvreOu6pCHytqVSHmdOO6ouSA1Yef5cy8ssYXyydwtn9kfJ
pp1BbrKwt09P63nEr+ek2YGhSWwz3pK0MAT5jstQPHuhBPwWM+36kSYSQdByN/z6Y0NH9GYfBHFq
/y56dI8kdx5pGyI3qSJHn45uaj6TdMgUmNSOxpL9y7h89GZgnaQ4WLEzYv0ZxGoWgyLdLsJYyjv6
kTq6DNctEj5JHBT3H5O7eQtjJ1hFtDV2rMXJDTgdRNraPSIdDZpSaEpq2SgEWd3GDGMZIGjBQp6Q
/A7nEqTHcnbMrWdO8/ApiZmyD2iNPH8aeDhJTeEzm8/SF0SkgdYI7M+GmlVsNwxUhVQQydGAEjN/
Aayp5/i5FzBDWcZZYsOdexYcYPm+GbMuvkDScV3vlfOONdLhvHJzrj+Gil8Q0+7DgDvX4A4KFvua
U2QUDvVjj6RWKdG/3d82bAtfNcZ80QYmTCAUBsVFp+x+SVq34EDLL9TrH/L5cTyLeFn27suCbayz
6dup6es6INHc92pASjmsVcDhVGgiECwpEbQ8ffKMt5koMok6B1KkpzZ7vFEnGWU/lage7mqg2LjT
DR2l8nGCwE8B0nZUg38iEMbvRfMQUgBriGhSLJlTQW7qPQctbUnniPaFSyghc2y55XB7Ef49biJ5
fZ4BwqS+C2pHTmJhk2IOx+pFk+KOQ+D2CSQfgM8gkNVNPHR27jkliZtj17lxIgrs8/MweCsJYAa2
vZt+HtZF9XeFU6etTlVvKWVqR2b6a1Zp5XNSuQ/vwPSuYshwTB9eBDgKjkjJeJh7lt+deSJ4Qeld
eDFQZ9u871GDoraJE14SuA80o9AXoQD9UwTLAwFWUBFjv8SqqKO77/qmrSse3aVM0aruxUDRJT0P
MWLQU+KhPT++l+S6GqgeOFwzQOTYTFrf8Wz0rQwH8E8nz5xVI/bkLH0Sk81aFOmc0Vt88KfWh8uj
Mr9WE5TRsE2e6zdCi8xeyzOm1rnM0n526r6y/ygr3jKgBCPFjAh9POlvUNZqavNmc79ZwGWUgsYJ
xFgvBsiiEo0cmKplQ0T7AY54oa6kceDeCwqq8zbKvkduOJVFrC2qMsFPuNaud9jyxve4AahJkCrr
6JYu/oJpD29muSbjidMtFRj2eHlNWlVV5UWIrbKAl1iN54DVtJLHygd378dxvP5K+MmV8g45Oar/
brQVBE0At+5VFmgpvALzvUvUnnoylfArSKVWkHP55QP5K7z12IJ6rSWVpYg853KoxqxdIIhLNgOF
dla0e7BYNxcmmrsQJcFLuWnUe2sTBtv2Pm631PV2oI8cXqCbJbmYYiJTjRCRAPSWGjOl8/L4UDPN
+SrGjO5JVa7XEfxRewETmpvLH2ODklM6ielFfOqaC2E51ZTtKWgyVWTpCJW2BDdNQYKcnPsmj8MN
K8lDW29pm3sJN/cbC0ktM72q6gUE6sdTLFuPLwxv7bNvvakVOaUjx9Ous3gllFLAWDIlMWb8wnXg
4yPM8uUEDdK6UeZ/AX9I6XSybMMsFJSO1khcaxIZvlouplxfN32wBhUSSR6fyBMGRutmyuJ+0egS
YEukkTBmWsfOIdD08WQcj/YdK5OS+fUQKO+i0Y3aIGSXTFWssa+lFUkO27U5H1fYp8yp3W9lk45n
OInPc1eL5gKLnwzeUUUiwWyaodnjEI8qsrhPNZ5ze+N7AT1nvyIF70QeAn43BQbT4zkJ+HBXByXq
OADVM5PjdJ4ea4djt82+e7Sf8Bt7167ZnlgEuKRXmnOv4t+dyzj64KOZ4Bvr6FppUIKfwQK0XDJ7
tt32bBrITM+MAE79WuzKK+CNQhJbru+vFvgVB9gKu0NSnM9XAu1WGy+YHf0TxojC/IDXH3Xw811I
rM+FkqBCFx01s5nRbLcO2VY0leV8Exc/4wyudLMntlcEiLKm2+xnv7qRFI1DzYquUcL81zdg4Bdd
pebW5BoBBpV5cvqjBG4bx/hJOuObDEOutY9rntYCu18kwJBXFqX5wpFG+v74z3GkEOGs5yu5d9oE
N2xThsIwzZM/HkWIIa9cYo64vq5GEBZ8SI0A126K+TzsUcJeAvQCoeLte1H60q1L6a7W6OOHNRBj
WzHp57GZ6wOXAwDpspx/3w42CDHOU4ipEP/apgEqJ9+LIQ3/iIFybRVvWXLNyI1LakjJeKOZq5Ul
goNuptY3adhMC1SMhEBBNifWmlvU867pcpk56JLMh1nExs0Ijd3fb3eyhEEBVT8yTmNIrxS++P8K
ItkteuAgTDl+Mt1gdz7tOBvMwPIypNhzjBFtw+sMrYZUZZhXMGpouzxWU5WiGQC4TcFj2GeSVNdT
mMrqkc+9YeSQxRXrEhkTh1KgcetUdC7yvjWkwZOSyCEep60iv6+stJ23xevHk2oMhMwIJgzCYBkd
50i6V5xim1ZMet+20InFEdb6OzpuLYGt+4egKJu8oFd5qRa0YpZpPht5eFx6Rg9Uqj4bkg6eZ/Ft
Kbf8VdGuglQY13gxSrDYwFVoZB5ltdgMBrZTq/hHOK2bgMqG/5Uv3tv87yA2g5YkvtqeojFDfnPC
zUrT7nsUh/LtlXQtEo4x5QCxJuZc1XlJ72uI8cil37LxH0STUr7kyKqMGcZKYtPJFfmqQgsmSJcV
NhHDK5XQSv94wGU6n1WEW5VxevjK+Ll/p3eK4rRwe+isiyhSUl1eeV1SGfo2N5XzLflR6Rgj+S3R
2CTt+cDGfhNFXF1WqExe7DGpHY47HFTxoBHvYQ/ghWfqs4qr1qCoON7adZO7QDu5nMCO48PbNVMD
pxclMfr3dx1idOfebUBqR32CO/PEOOUZkCcx+jTV7EEFtuNw4ofiRKMwBM6DdgXRAA4J5FrC+5wk
RmZ1QE5lWOoN5meCRAEC2pqx/eVT5UggAsTYSR5ROY1M+sybmPNJYRaGdjBdmu4J0fJuCgERwvg7
Z+UPT5qtn3x21ggv1J8hueozBVPIvLCfmIiAi6ENcocuIcsE1pNdLVqLx/wDwoxgbMwV+yT7DwQn
ZyA7IkI1bHgoXGTVI2KSHebtCYuC+MKDcj1i1XERrWEOo31tlZy41swKM/+bQLa8pR2gSqnvPAGH
qv2zRHZvBeb7k3gnYhPQZD+EjUZBRrGFw9r1ohKkzn8NAuN4Ah0TmmUH+Y62dtBY9W6BMskdnBhM
DANYhEcCIFwYCdZuRdCntgxrgYoIKN6+6oL0ywOFf7BCHBtLYQdEdiPWJ/qBxFwd1dMuUyJ/6Ouh
QO04xlmWaj9DZ/mumr/UJj99N6DEMnXqARNomOE3HHsyzx9aGWTOUd6hhBPpSGwaZtG5r3YaAJvm
+jNWTKEgCDERDFQMwoayXs7MzSdRfxJDHwODJ9eVM03EeXCAPMAk1tLqoHNmbtKEekUe75XMPQcJ
VbmgPwp6iGxSYc2Vw4hv0gCWPRUNlRtHcfz0iRwKeMR+qn0LGB6EitvGhGoKSvJB87ZzGMMf7wyv
L11XnUjp9hLCXNOiYQBHgaTXhTt/xE4o5/F7VVrvUZAEqYU06x7VP/inqKJ0Jw/ZrAZ9QFZkKSdT
ccMusPTUaAnOUWEOS98fNn4NlwTp9ObDKLnf5fHTx1XxCox+JcRx75Dcjyie20S9uXybN5+6eXJy
vo4rCbLmviaGMy99WEtdch+cb2L2IRtayt1bESFSKjuX8vf+aA1GWl9Cp0YRI474LByggu8oNSqz
AljveJWwH9wIn3SdaI2I7Htn9ciTaVf+R0FUxoH7640Ul+MC+Vh49A5MxaZGNiZcUfTuDqZHzZke
7ZtXVvjVfzbxWCy9yUXZBETFugDwxzj8NB4HmCxehiDAVZci8tbvK8uEc7aJJNKom6jkXg+xO8in
iZi99vluBU9bv5EYZlkdEXwxoU8DOs8gK5GFbH0somolBmnBgcRsfCfZVMUbskZhA8Ul070q9GxX
HhQpLgPVhlnBIxVK6HdGY5hK5UjErbI2A5P93nf3x4QOcQbMR665UFKVgiK/RUXNEeVgBKwAp3Bk
my7qxvKlPwZSEh7Wjk1oPE8XYj44QIbklql+Vg5Fij08MDTkg20cMQz8J+jMqqsTriUuyCVDJpoG
KAsBKmoALcVPyKEjGM6fwgBnoeypQJrtaZwYS5A2LNVEL9l8cuWu4ejkpJnodpSMiID8jhpiO3iU
NCnBj9QiZoW5YvRjUfdnIRfjIQsIAThr/aIne0yikNVGOJbgyq0KKii4sPQ5g9t23dZkYBFDTdtL
xUXHjcAbBhd2RKtI8V3RISdZwKMeza/BHu0CCwBW8RL1zU4yS1lUhytQ0wDC9bAWU2eD8sHQEE0q
1K0MLO70UOqu7IPQ0KYjj8BnLC+OTe3JCN2rv+DVKUa7FtacKEe3JIgDHnnvLRBq3tA5yV2PXSgP
1kvEuP4qc3cIsMnOKDmlyfcoFrIgZZyg291Zo+VoB3pwc2TTIU49xViXbdnwlaARoQU5OTs7o56v
N151wedwIoLal67/QUkiHLyRBlR2lTKDddBzGQMvAK6sqjRX5PzaAZjms5il2wDSIc8+891nWI2G
wnQ0X+WQ9Lhml4sAYi7Eb0zSP0PkjrtWd5O+T/jkKM0WOm+PrTvR9wEjlvHB0IWkKG/CUTGotVDx
m8sOlpizP3UoaVfVmWrYga+YXKnyqiHPx1EwBPRmyab8hsK/1VafH684zwSe3YH33YIDW+n4hMyP
0Ub6145Pe6qB2E+Hdx2Uk1pj+efz4RZrIZPoyD2JE2Oetd5QSmggkEhJRhRWpTo6MqGKQUMOjgGk
QUB9IVPBjS4qarNopXNHpGucpNz8nHJpIt7huAGJUkEonYV0FavJS8UqCwn8MHfGR3u5dS1xbBGq
zLNN2BgMpPhcd/KFYtHVdtjC/HlKa2kBR68PRM6nSEujbbOuoOT1XfYrm3WOWdGIkLMvw6ysT7R6
UVOJ32JyYAht1QOvGvPyTR1mzKbZ35y9Fy7BJoEuRHlFJF2VUkDHK+AAaMgAwxG6f4KOm4Q3Xw5s
m6jeEjiwwXagAkNM2G6EvePgmUSLkNp5y82Guj8WOEPVtC6RvfMJyro7xkZpH1VXIWx4BVstrv/b
mnBgeK9EDXf83pHlKbgu147nzfDHJ8FUaqo+G53VdYVr51IFG/n0QdlAMa1qBdlogPs20NvlqLjX
zUijRCP728C/4F69pkD6/wtC/wtmS4wCLzQq+JXXBDwZjDTi4t05gM+862lZCMKH4hIyBAxpBxoR
fDykRZOrzKFMy8YV/fi304tTF36/HTc2ZuXE4Cqb5aV8L89GOa4N8kOHjofbxZnn/ZZNhspUVbZh
yLy1uHWbH8mLonLZ8aF2f3+p7IRMYZ8yVRgVi4UCmJWmWqtpJmSQs4E3QUlGYPYOyy5zvZKTytdW
C0eRRDxprdhfGaEQ0aSTJeXuLGOelTa57Po/1Y7V18TyKONFY78SsPVHJBPWM3udrB42HFvqe/WR
vBDIw51bjKLVYUbqC4YK9qNB6yyGq2uKO6rhpD2CQJtTERxMNLwifoNtzKKu74ISlaX2sE7oKobu
kLLHmyevkCp5/X6aC1k3pHFprihz4uL0mQE293MGtD95LdufLV3SdHcoIKk/BfAiqvQKK1ppAZBx
2GcX+cLvYu7G2uTLgeK7pRuI8rMZTlEw2yL1KRFZOY8CNc+FOO4IQL6/aANx+cRk6jgJ/PiWUNbt
kJctG1u3dDl/vlIarT/69DKcoS/IvAlg5bfcCvgne6rWYTDNdM+s3qjHhQ7dx8jS9uMXZcPKIU86
H0K3h8H6D/Oxocwrem/xtu5mS4hDRV1wtstd8RwjlNTQnWWPOFJ+QFI98Zd5jyHPYq1f5LrSNW/F
1YbJ/H4Rnvp7J4V1xRfND+sxidcGpQVTYTzTeXDhZPAPQVVuw2RGPhQhjZ5OEy9Pc+w4tlGQ07ay
p2/s48PI948HJYo6/PqvJ8ptXXzWmuwjRdE8abiYKO9i7D4+nwKh2OGP6V8Rf430zrKokmxWaDtd
uThQ2umo5Wf4Kd7tFRyKy7Z2qkvrpt7qnsAQ3CXI5wLrjrP6cy4JTWvNdkonYTPcihKpNHq41R6s
vu6Uc1ejxMmnK6++JgowXJjPmsss9TkJeFElVDXU5UELjH0Ogkk1h/qu2trth0FQiThdTiULtO1I
iLvxNQWESn6XHrY6Su6e865Cy/BXX/n3B9tMBKusGEI71IvKpExYHQqGNBiZ43d65ZW37pwMuor8
9W86OkroKpmn0f9W4gWWmFPEKg1jdxAVf553XX876kyKCIct69dJSsD5WvPsNhaoHOTkFffmszlz
0ZrLns+BD2oRfPHU0WWMpvGKAkPm94pnE8NHRm54Q6Jj2YzjUVnQiElw/dE6b9zqFRwSgxsJIkti
u/c265eqVf8uKod2HxUsicslKcRWoIH2BigU9opf2AtVujjV9LBIBZFDXR5SrTNfahH+5HzydO8y
Sf8XsBMNXM+LoYatgdRhtkee6//wSohzvwUZrOON+UqjT7KKAc2o4Itf7IqAoJnnI+6P8NYaVugB
BFhBYCA+rtBwbYpu/Jg+t8H7rsUnaoAGaIv+mZvZqwMrmcwAWKutSkBlt4dZo2BAJd8fKm8d//I/
3MVHj/TCAfqvvl/sYZNqD9sWyTHjAZtGt/uEtC3q4mbXgHGw0zkMS28fGGYdkVcvfulMjGhIc31S
QHDzWXitb7Zb/NpNMNFUo9IlUscAP1bxip8VnmsrRi9zsOk8RroOn9wnsiYulrmb/GuGCYpOmhwd
U9M3bpva81iK5ZtPBZqsD0p6x5ZUmGhyWApRzJDdlVym52IMtIFv4axWMIVM9Xik9FjPSURleemz
AP9hK/BZBoi8GDbFnJ21JCPMxv/laD8alQpazfI8fSW53Cky4ocPqKvIyOHQ3lPtWbZA4kffni1V
PBaAakjc4FW1aLlyLCDIaxCjyiKQnZgXom1eqMTcOJWHn2r4YLPsuQYu3bWyJtyrUL6rQ3tUH4t8
R7bn6sswNxYjY7h6ZM5vyBvMbLcl0S1f6GEsZM8bhRPdwS8HRZ5bOCYysfa1w+MKVsOG3QH8iMic
wkL9C1DwiOy7yx+iCqWdtR1Z38adFejU/vi61ar0K9xpiN5bLLrNe0vN/58R0D5mOF21CgweB06b
knpFNY5yF0dvdCLxVoeHT+MSPOUFsbi/D9wG7HxiFmXjl8sP2gOjZQVffzIJQP283SQ/iK+os57W
8gROGLv/q6lb2mm0jGfxR6iS64crdkQk76OenjryWVL09LIIlnJNTjJnB8KZFGACURDmAc36G143
eXVB2OHhQ5PpvNSS01oE0M+CzKZ0dAARdvyxeiVdpR7SbFbjTmZ4kFKV8iuj46er02MeVSq1hmQY
/ZI8Mk0rgh+Y1FGWtgfh+gmr3SCAfA63RMZblxaQnqoSmjK0dRm/lzavzHI+Ayz1Haw9yjtqLsUZ
cvWsW9/qwyUaQgjA9LPKpvB7J8uafrLrGkbMeilaIiSu7wDFZ8XkyBcrD69YfZ9jgSqU8U7qe/d/
3MGzs5Ph0dU6D/RKXgGbvIHaA3OrMcisCnrruez28XvNAHRly7+08BKSV+dNoJkc6LBHb/vu5HxN
KHcGTsGrj7W6g6gGGYPEuLalKvUw7AnPYQBR21MK3N7lIJFkCAu2IYJR7eIqxJRcPKzUsy2nwZ/z
iG4tVjH18PlbzMFCXc0dxP7rH3Mm+8EhC1P6uogN1lYFoiU08l7gVsT+8NfG0VSvTaIdVWBScYt4
lVF/xW0a2hszc2Dsdsz+qyNS4ivXyOPY4XHbhtLyK9zidPS5tppE/itjxDkBE2ra7qL4G01Rci6x
qKET2Is/SCxbY1lm/f12OGiHhFFE2cLAXKQuCZT5bSNBW1mSMEEaHNQp1ksc2HeyI1iETMX+s7EC
YJ4/7isVxxacRYlDjn36K8IBi4HA0WLKdfu67VBYuHcDZLGNk+zsN+lsmJJMnfTYAGl99u4trcpw
Lbws2/nNQFTCJUSfWDCoppopSbWCAdO6x9C6STJV3zLAWwVT1gZucpKUwNuaalmL7iY6w0tWZOBR
7vJc+jAGiwfzNV4RPYzf2ZD9sjApLkc+6ZWxON/MoPFQe9LDIs+3NTmfsYFCytAHdMsNy3XU1Sfb
OjZDY/0rx9Oy7CxLvCz7dnsSITfUtYQ9BhCbjunZmxTZ7lBK4xC0aN2FCfuKKIZmEFtSKfYbWMmt
TPY63n2YRuH607E7LfXjEPJxnpRVH8ZIUO9bdDUjWeQaH5voWZyWJ3/i4T/4/DH4tEHuQGk96tvW
0e3WU7AaQA6nlT08DjpEWR5h13VYE3baeNYup2ygT8UVOoekSs0pkfSrbBqZBV0pHC5WiJSmavcl
RuF87QYLmBZA9LUNurQUZy2/b4RCgxx5I1hCc0E37w0yXLXRfCfTlhpNAeWodIoYNswEPecRELoT
nfeVzHFms3ERLwArzqyCKu/zddFHiCSZ52Iv8/RfZioWdV5lIwITCAJxrL8yS5OkqQMG8HqPlHm8
YOJmAyCHde264s3XmRPhUzvH/o0FkT7bduLqewLnd43jURVxQUFnb0npGwb4OsDzHHquZ4M97IGU
owbsUXOutf0Bkx4J9GfU6ervoQUaNgFq9mRjjb592cg/7EObXGsTdgKc091Ej5rIyuq6QZD9dqXc
B/Xn8gnS6nN25GencJrHHwl+vyTs0yHHrx5SW7yASoASHloNi/lLGENEt0DxoVx9QuNaZ0Nicylp
CSG4igorK/nVfJSmdspQWynAyKC6d8yzeKDvCgxVNpru8YomAKXaTB33b8y6A313tD8RMGxWSdgo
khKpmz1Hr2JVBuRBrYMUvLugfw5Y01GHn1wRcWp/C45OBW2oxdM2AZNUl7rbKhpjiyABPrMWajd+
7Z47MSgGOx2mCzzITgb4KRp2T2WSdANuUNZJ5/qYEbgos0byLGPdpQaePYFRKFhAf9rAbIsM4zIX
Yq00i4b0zOa/ORRtXkPLqgL+areQq3eucZpTS5IwzLU79b8vpMWJf+5QriBOaQJyc/rq5BhySNN4
p6kKBBj0/GAlTbKQhdA6LG5w0knFHG2V0Q17L7cIB9jXqOcg4fa0OPn9YZVtsx96BzI01+ku+zBy
uqhfq6RtZ4lpYWdiRoLhrmc/ToaDwEK3MTms0mxL69ARSuX8I3HWjY7hdPujXX7UigJTo+MgHnq0
4Voyc0Pu8hRZ1UZQuZg3klARVRsPRrNmk6k746g6yv6torcKwZMLwtIojzlGennu3Uv9CbBVNAkd
6YVxInuhhuKHLm8aaNdfmGrt32xH3rchVcpiijPsLcG5oM/L080zn3S6cV2Fo+d+mZx07E26zv/5
93aukgoOicns/E13VgGxOBth5zABzIO6eMO1VrZivpBkVghr9MqxH3e9pLVHdfGirjadIFeGPGID
UYpBASy7/9L3158z3CTou/MCE3vbJqKwVrKbTRrbkDaifyIjiijmuk1hUGcgC8Gmgc9QiHPo7cx6
FaFIU/Xja6Eklyqgwi+4oW5TTLmdWNf6kRqmkVjn2A0RuyJU/Q4YI3cTBXVvPtMNBGtbMaHnGXkf
FCgKgKntM45WHeA0fCqWUrCRUKn8U5kGA07IPxGHIBOesAesroU//P3xQEkzZEI1fqO/pC97zfhy
DQjQ9XB8JesaORNlrTZRzhmRYR2+F9hch8lJPwr4tNV2z7j55idmCOjSWmP6zxHJrBOwClXY9AMX
MDJsZeH+agWzEb0MbhmzzF7unqM049NLEjTmWu8fzey/RbJMolsTtJmnfaimqZ+IHsAYjaVQFeHU
MSWtRbidP134EeO5TPP0ympdF56f6Ke9xpXFEL+mHljx+diI8bZdPUMzInyuo2g8+TlddzAVNhRv
FXdEKR0Xh8HEuT1GTRzRdrCw8LgrptLnMfzDp6dY+pIJb2/FqS8FpxMsp0AWXTF9PO/MpWZGRyQ4
2YlQEfe1+ag9oNOzY7jz22xBNuV9MTnVaduJH7Nr/hUDTh09hlEP/Nu105Nx0wrU5cR9oa4Ry/38
J4gwufgTbMnGIndxYrCoZQSiwwQ1FbNiUefS4MRlaQX5nocuFW6K1/RsulYluWqc7RurjMRztGaX
/IZsACuiBRgQ7NurfUurQrWzomMHLAcV7sDiVZgleAaYDK781ep7DOVc0ve7DDnA4lxO+J8/DzyH
Bgl+QqfHUI1XF/7kYp6BGVrnXXHnJU9FF+s96h6uVTAcv/+s78xr7FXUc0JT1ZB13VKJbSedC2Uz
9C4X62xSrdwXy4y964gsvJxE+g7381Up7JGspJeJoS/NiYZJZ9Rm3aHI+QB2wlwiJxGDSs7N5U4W
qYswlSjBJPAUVKt4NbbulCmsGm6D5xEE2b77+BuCImcwYizbS7ZKWYbbM4AEh5B7PTQw90RSSbOW
otMEKOpNsMH3I+cx9pG+NWkIABzgVSq02wMQzeywa27CKYpTaQ3Jj7LRQZtz5gCe5txjGPweEHYr
4eW2UHoDtZ21RW74zfTuZ8hTxboIvTTLgBBUQtAHOjcrpYdWcdfSDw4XU1WXEYd6/1NKm9ympMAo
/wNua6dH9/JlNt0ozSCqtQWBDbIVQE5Edt3eEYNKocTtor9YTbEMYVl51OmFsjPOKdGLcvl3yCor
OtynJhD8LBmHWp3TkgoN62POmeyb1wtf8qwbaElQU3713ssBJ64nC0pvhS+IKElx4ygH26p+1/7E
ZYLa++WH5hafIcZecezVcCNI0lzoJSItg8V5cMWvkboariPedv78CnihPZTYRzvY6Vb4AHyU5F7x
AJG/+tCtUYvSPSzMHur8W4kw0Ff3HkZgjwGblk6U3FcrJsHpB3Y4bmof42Kw2IezYFwFI2OOuxq8
/PF6z6o99Dj33cGR0lz1CGFQ5jGJSQ9J3yZi4wpPxX/n4ZO5n4wv+sdGZnT2VBE5jZBI+ZK7xUaO
/Tp6sgcPNtebvTg1kIee9b4XxY8MiKsJmDQuJnAI6Y3oDSzNOxeLWQ/Qhy48nZWB+ZBIZLsi7mqa
/i/h/Rb1amSJHiiDtDSphVoJECzjMwIWY+i7fm4t8p5Zh1rixkK+QyeYJH8dpGCuOyyaeaTbBklB
aR3TAYlVA4qxk3+fgrYhz1q4ZjujzRl/xc7+/0Ce3iZwjRIKsNhtPX4N/iBXlbsxNTctOx1Os/K/
/42KDi9Rlk/oPT/gUwjOSiDb8O5kVJ+GxOmkprslsnHzjS30eqkPnratsLywd9z++1/FTdEJa7c8
BCx9Q5SDPRd7L3l0pll/aSrjQss4/eTmGbxeT3wb1hjw7fzngaLnNAKqXruZb7AgY2tw2v4VD844
cqEDrM5aXT/w8ClOp2EUGrGghUurw3i6ym6NU3HJMIwdkdLQiMBvFL9OiNJGuQNNoMk8JxdG6oP1
CEfvjlOPh1Rg3ZQ0WnMegWe39xtWWhjLR7L7vBycjviMfZUdlCttINMvjW9r6oC7mwuENEG9L+O6
eMXxlqB9YA0jHol5/MMnvSEqxHt85smCX8vtav8J5sTN6V9gfEAq5kDB9RldNI/shMNY0chcvgbe
p8C7VhA3Gyhc012p+MGTFA/ZoJCJpM0miHVbWGC4aLkPaLeFtHYJNHBVcr8l8iw7xY8kWxWqXF5t
4Y2+Qj5NmLzZLFXiXquOj0WReoG7QrFhQiRiXI0PixqXuAjoaW/pZyIemKJsSRUu7qneDqrv4ud5
R4K73Q4UfZg62bcJPH7cbcj7/6VxXHEHr9PFC0S/VjcbdeA3eNO87/x2DC0twla3ob3ffwaNKTol
NPC7YUSA7R/ggXFT7thIJq+5qhLcPi6aq9tY7o1cuL0Psz9nngWXSfma1ov+QlYHPHe44D6AHCNz
Trk9LMmaRTco57kezdH+JUFxczRdc54BSXYIPGw7aTP8w59WGst4YwtiomQtnVMfKaGejL7G7FRI
Hup0ntxPfkaF2ym8yiZ7B26qDN5kE18x1UqNVgK8+ej25YHVAEEkGC/371BXUwmuMyZlExYhT4+7
ouT6JC3BdmxxK0NqwQLYb/Qiq7X9z7rWhqX5t5rCtj45pAFrXBmbVevFlXB7pUIidLWDl9hCdWU1
2f2zNs5QkNe2H1U4fd1dk3p/roXJQSJW8i5RKXqY1sUXRZ/ggJcfpanmrJTvOkMvYrYh46f1cu5G
k4a3ywHSa603qof3OP5ToQVbWGf5K1O5/bWihOyydfw3DRjEn9WxlBWxet2uoF2P2AJezOjK/76Q
2T0lh8ac/pzJUSagJQ+ma8w2gNkvN+3B/tULq2By772sbddrTFEcn0C9wbjYbTOm3/czQU0O7LVY
68S2CVRC6ukDekyNmhbeL4o+WuAra8D1AFfGKJQ93Bh70Ogz6MysM+nvpiYFR5/Pdvc+i0GfuYiA
8sJzEJ8zmPZlOKBwcLtn5QPJ+h2hzZddz0+H5YtR19CB+5Jd5ZVXByBeaJZ9Bp0aAmfI5dLT2oho
+l9M7gjwRpX/0ePMEAqPawZKC5HEIK4nkrnIf5z5vBshoOXKBlA9keGIDzb6yj6E4wNFqlvsteD0
ig7XMGiV2Chgtx1sCyMiU1NLhTFEs8xz+xiPovDr+CxHR+fOQlnDxyV+raBHqzedwrvYBdnrMvyA
+rqsxaSDpFmrSBBP+ARVatnkFa1Iqyq6ipK5psSD7MB5dt/SIo9mYdJE5dZqSOn78e956SDbvKWi
5nW9VILvPmDW69KvACHH0fnNmOFAh5C1BPGp5s1Xl9W0Io9edjgAlQ6qqd9RbpSOL/GmxW+LW5BV
vmxdUrwNhXDcqZ95p7Du8gzvSObacQwmDLy07eC00i2zjZ32nmdiXkd16l3btVMadMqGlpLbOF/H
rzWr/xZrM7VN5GIxi5wFgDbXNiwCNeiNexQzR954KTwUOore/TMtmKrJwIH2cTXUxs6Xrds4nZlv
25PnNHA6WSO6MWbkBAmFRzTjVypy078UtCSFL2zSDK5aJAWnh4BfyfIg3FoEk6rryYgQTfzFkTjr
jlPHcsKQAMZ/wq2AnjKq5gwWVl9w7QaRLXKdOqkSBGxD6eoc72BvRqEVLU70AbHjmkpmFHJ2SXGL
cpkM6ZQRVx0gVYo+slajbF3ryGfiam8B6LKwdhn8yYhB+XSZ9sELPc4P/zOtssjOjCO/Zjuk4lYz
jzTmcdMcx4LsQZ2mZLYiTiFXB3Df9iVhVUgvBIqRhovLax4wfK849pVbnbaE5TWI90xa5y8mtvQV
h6sHoiRTfrIltacEjYRp3uVnhLiExnmQXK2j15Dxw46v+YZ2oHAqexTnOhMaterLE67Vqv7CQEEr
Tq2y4UzKgYWdR9GcVJJQ9bA2HRyg1oOQKn5F7RVjsu3mJ55OlExWaxJ+kmLN7NTHF6LHFpz0IRWj
U+rju4bYstv783o0uytLD1AteV7RqznbYK8NseNRmUqTH9MQWJcEbmgrBnSIhUwUT39TeLFQDadf
t3ws/BR1Uvk/kSqnqs458RiiU8TEQcFvDpStaXh9vhb4w3rOZve46p2yTsPCVxrbe0BV2aTh0FPH
FrGp20o7G8Cvmuc+hxQQP2cBT6MbETROZo9dt9D34i3KWt0OL7pAwCW7qDrL7B+effa+W1qSAsaI
aCZD1h5t1klevADpjMRSAuQIkNtmOKzbTDy+9xyNzNWFgFzMfbqVw4tH/JvMfNw3XhP6BOpFfkKA
gOhVSItVE24KQdm2flCdc56ynAsHkew/M4z5cIzKYnLfrhqdhAPhP0bXhLBwnU2mBV2NuBZtWiCq
gAa9tCuKBBA9/UqJeGrXg+bIGnMRxPo+c/1vLmE50bqok3m7sbCB9FPifsfJQk0bK0enSVQfVZhj
KnhcJGmebp2g7SrZF4KDeVu1MSCa060IKYG/SAh0hWkE78nhQCp2442NshQaYzS6Icnles84elOX
6jmOPLbP4i0erm6m8ehobG91Lpw3dvqRf6xydhmNQPYN9mGoUgFm+HbRPb9ECeorBO9akC6UZ0zp
IynsvQ+iJsY37fNiYgZ/WTS9FkERE0YqSHa94j7nOvHtZjkmuj5IOGEAsNaSzH3kazENlzwQdr2F
yhIUcRPli1uK52Py4G1qbhsPxqW3LDuwAW1+I95AVXKdpWjf9xPfT1TKVpPesbTpj5PBlpMOJPKJ
3SO6+V/07+7ybOdDqJDjLsP5uN4y3M6TlxSOblF5xPRGpMZP6aNRtVsS8mooMxWFcL+PlUip/e6L
ljMzeVfTMNKf6L2i5rw/8zs0GDi7GdRZrHs70CNe5TKRjBfwa4CAPKzK2B85jno8nOZifVSOJ7wG
W6MB9hkL9LhvxeYGb4lZAGRVmBYG5LJpIUx9hlbKt8fJ0070CgXN3RQdv5g9edisp//PuP5xexPN
rNOlp7/uKejPW2G7rYWZOeeSqWy88B11J8RRWe7OybLf9Fbs2nG0EJYU/11QLpC2pHjllwHOF3jC
YObiyeYZB62aYiQyotHq9vtXyewc4IeECfLmN1zYOIK9buSeqCQVpSHVOz26PJ+t3XGCYATetHbu
ZlfzsSj32yMGXxIY6OVD9CoTRx87Pksri0JUfuO3Vm7AIIhDuEy0BTtp/i7cxcK9Fqxu3rPBJDYB
F3JW0dNyWyNxxrocHF1/jhBz4oqspqbIBPoEsZR1O2Id49RtHNYJg4nZV7NNbhpPQtJuCQdQ/Pxv
eAnqideYTZiVawO9pBCYC7w96UzqhSaqWTT5TuK7SqzMkLXk2JBQuIJiuIdnHr3TPaeG5va8wK2q
jS5jVvyfrDaUrZ9AQ7R+HS16DU8b8y84pybWHdAKjH6Use9G4ZfB8Vu6F4BC3tCibL0hf7lGU1ph
/on/hD55Plulsi/BhCy8fZuu0BVAQZI7Mw5/jiFKMgIJ78WEdk2sNEW2yTQYK6uix8iQ68xv2YaL
th85N5/mNR+ka0KS7iQa1CuFJaaKKaDYLgfpuAm2ZUiEhoFrD3g/x4ZxAMwv5urhGb8ffNk1ew1e
I1AquEGi24OtZZ45/9bXrbUgMlIrzMoKvrr7hyc6k1Nu0SoCOOAUWESI86fledUyS6328GihGPCS
CyciJmuoFmJFfXiHX73aQzKtSHP4/EuCOQ29nvVNVGYep3n3/e/9yk57vqFtRuCwlVjJeNk0ut2S
6QAlt7sAqrdPbApoGLlGdcBwf/lMFDncgV10vAC6ZuK6zJL3bkYRTrmLDUmUygf9G62WZOcTnGKg
ZV0qSq+2ukkuS8oWoHnRMFVz7oQmFEdTridSMszKr6qeXrMteVbribwgyiTTEvoc9VVE2jFFjzIb
plojIam1ps8UTWaiWE0BzKJ3cnl+2uBeB8Dyc1NzxRJsfHJTy4jD3OH2E558jLi2wHKPR5TM8Klq
yGYKpwnbJN9E7MqkTlnjoOOCTuj7uT5xix5nloGhhsIts1ojqpp8iCGPMgGcKbTMGW/mMsZ+oV2Y
5aIbsxiOnw3fAugSF8zs6DI/rEhVUjT6EtZFwgudaamW/7TvKm+a6aNjTwKqpeex4r6RV1lH8x0j
KSkknoaNCxbkxQasHYj/aQDUEr5b7rNf8qSGBiuzbiGEMn7TD5XTRfWVd2TzCxoIJtTSNC2JdwHN
3LvT5HQX+bz7bfz94TL7q3rMyoo6yyLCd3f4Ha5I90YZhvr4a4Gp3lYgfILFhAWFHsNIr5TIUilW
7XoowrYnRc4EHFYFalfFUIOaBu9vt/80hIOoMY0L2We4AEKtJWIQPkneOqLQvqgZJD8KAIxhMYgP
l+PCRPYPg/xnD+TVOKTO3PqsZh+0xPangAav4pDyUU3CBujT34CgMvAtuk+WOkG2XreNgvgrZSCw
JxlrrTDrfRAViz+Idn4ZekjBbd/CfBAIS3g1obE7VevYq80mdL8AMglBkTMNkCwobnQtXb5cahbH
Mck9g21thYlCSkO3cXuBYp+kpx6jQ4YlO0Csgd9s5zv49JfIfkQaRHWHtzD7lKh1W5mmBrLv9V1Z
rCru2LlrPizJh31YFJ9qzaJK73m03aaSxGu4RpGSOuLvg7605I7zGWVVrQejHVY/4mu6j81Jrg1P
xJEiSHwZQk2bStoStdj2pAidIy3nuomgM/4iap4puyY/Ykz/JmPjWisfaEMKgoG4frgs+DDDXxOP
emBlRJvNDwpzuVJ1/2+nAVf5ODnynawgcne1hbFYMddhrL//XUcTxu56T6m+r3rPqBKdpyS5xJhl
TRoeW5VoLMvF2B8VIM7sWuocN1WcuHgXgWyUz639t/UyWIrfdf/rVz25xFZpsZuhMkaqQECMKrst
sdsnHqRBKd8icAU2lZZjC/04rMESuWvVHFNCRB0wvc4qJS1j5UMOh2pS50uJ4CjBDLeXa6M62ZQz
99Lv6kYISJgqJUGA5Yy/RCtkdZRC8/wo1j0v2vC30R99K95OhzR0nk2w8ZCtZFvyTFTm3jxePZy8
Z+QiuNJRaCVIBAJKTNawgQ1O1Ujr2XKKDw1mrFzWbOvPQfmDVeXhiAAulFyikM4rNJMjQWmTYwDK
eHqWXmfzavljKLhWKg3VFoualXSuLPTmvO68Dc5H1m6v86HfjeTQes/mf8JdtbhARGXsiwmWl3x9
pNCuDPJhdAwwwKce/N4tuQOsI5pdC5WU5UYqzDG6d8H2aVs1cWAMlTh55Vz4zJP9otxmDa5AELQQ
yg9SnLI0K5WHvmAkERoNLc7kWeto+Eopi92DkLpzFycc8nsNN2bSaq949wQ8aAhzCo3ytB+hSQH/
tvAAioLs4aasjbcYP+MKryLhnoJ3bGYB/vtZ32B/eK1sWYVDi9imtbt/R4kK6aQB7032SrHGx+M3
OIlWJGA5IUS6QL2MyzUmuXWwkY/hP8RUWgAC/KKWqjaZ/VPy3uhy2L3pOFAeXmFV0zNHAzzEStDN
QIyTWT9CMT1z4mvYEL3R5CmbkLCfUJM5SAJORIpsmDLN4OKXIK0iIG0Rz+I2ucFQ5AQn1moGgMIP
WxBvHGM/YDe9Te+OvDjiYHxO/ytki11idVfqY4bZHak9nDyBNfQrlORFta7Jdu7q3brCbG/R9mNp
cdsTqsdsEH31Z1hsLwPRHF5oqV3w5ZrXRNHX4JdqQtRbiIgPXf98QAKkoJLMoAl4y1BLBgAsQBPx
NAoy20AdYF9SUGrh4/hTg9vvCsEMcax4PIBRQN24+NHjdYRheFjOoRps/5rvwFlwJT1FQlyG8bmC
SGnJIwl6jXsZhRjvIx3MFsxIe3KZijLwo4Q652sGpSSBW5c6yWKjYY84ZT9d7KFBrnveVbaO3+o7
mvgvqSf0jr1h47EKYetm5SSrIwnIM6ULHy6RAhVLx83V3Is5l9yy4cSKND3azzBAUyJttZfPSzDF
Dy4GVR8+Mj6Adxoy77p0hNpfepHVO+21K/yRrMmJPMXDLMxXS6JiqOf1xJ/8rvm4cwxhozbekrcK
++irgU/k7bXDtjuwlEiua6+IuAf7rfeh3G8cFKOFjN8XRJWbWNyDXvQOoIh4o18Tm6+4hN8FZdNp
i7CNJCbYkWSkhdCyEWLyHJEs7IVvhXWo24M/4iUQJjfeXy8I2a1sBfUm3Vk6wpQcAU4UErBSY91M
ktUKTJ5/TkczNMsfx8bZ2KgNY06VE+B/5q36gSNo4UD2c3xT0ZZbVx6oLLrljE1kLUlZXd3nSro0
dXaQxBnubOGYuRkb0WhRPzErYSz6BFFuu97qSd3N5wZDOfv2MZ1HAY7NF6ua3/PZjSer5zk5i0uT
MzximYjpfqZp/jjHWcCCkKMXB80XGqTVGL3zbczudimeosSRtKgej6g9O5Th6AIDu/MRS/5dQrH6
NxLaT7WBEAMrcsSE8rNWZp3nyTH5B8dWjRogk6RBziTMANknOExTFGelRnP8AdKkke6+Sm7uHleh
FGjkRg95855S++lr68Bc0An+TtuJyRBWBs4X5ycljTDQBi1U144ZZ8yTYW+VhK3PlOd8ge12cvHf
1depArcBQNOgb3oaPchSIatmrFB3YzXiLbMdL6mODefxdWeZYa/OxRV0f8L2W6n5xkHyPvnzmVg1
gilgonzLafDGdjKxT2sRNmvIZH5SEKcDq97NS4d3nYBRtk7giS5plKZINLCV/Zm8fSNAUYWz8+6J
HHJZ/zvbGp5cL0PgIIcbGysFPO518P7kUVN1ZXtAUutGkIK6SXJeGPG4Ucj5buDN2jFZxlUvm7lp
9xmBjuaYW+QMlo3o8Je0YlurIn6QZVaXT0PQrP8Ew1giyZmTN9P/zFWIVxzfJdrAuIBPM3yZAXFN
dKDk0L8fvKsF0RwBDGSkMmODsV42bGRniASMyy7wP4uKcR0xHLrUbxfMnxXLI/KUHLukeB90FjR5
irPRYeW3H0kDKDJJ/I8W0zSG1kx/eEyQOPw8m+FZBzYhcvAdSQEKNntr4lWKBQiM0Cids/Zrqk/7
Wza56Uw+C1adf8v4mG4/eo+kCHbOkq4BAmp38zIYH0uL4WEEXs7MaX7uci2l/2r188SYVeSNUslZ
ech+clNUPdeeEJ1Sh3L7dNiwHiCCFaD3j1izKn2diPzFKcfTOg41G4vW0mpl7flka9chTnevxJeq
se8ABrGxVPf1gnnk02b3OojmpxVH8Oql7jwrQQuZaAtgJZXoN1ohe+hZu7wXWNFSmES+0nsvFDvL
f8A1X9uMy4dIUQ0TI42hw96WpmePdqjmuTTaZmKW3WmSlMMOqDNPTlMdABQxCeqMmflAsSNoI3fK
vLBbWPu8dMpzywShJKmyOznvir5/zapkoLPofqK1YirCxsP10/EFfhlFLsE6Xp6XQdgRZdqG5E5Q
WiL6d/bMP4CiJXOxg/ZDE8pBUM6ZowEOKbxNmlEmv12/G6X8mRqw39m/vC6c0GokxKi6GbisTvpY
dhsKq4fo0T6QoZt7vVJ+kwerZSyFgyNDryLRZ8Qj6sX6nstV4nuuHmzn6mBVZZM2iCSTVDRbvwPr
M745N6ZcZbFqJhEGJo3KArNQ29wTJSMvLYW9fRX8AnNNCS2m+whdX0RR31ZkIhfpJPclJzwoIHLX
KCAQ1J0eyXn1Il/InWBsHnbQc6mhR/gnj+WIcXnxmb9PYVO0e3jGXSGXNiFPRngmvijI1byZ0Clp
mq/4sTDoOGyL1Ycqvs8NIsVB2jeMWU8eFnSxRA4T42NnHHYxo8luNxp7uEqI09LOLCHH0C3z2s54
PQRSWJTb9uBN5kad3LmvsD5UgFUvegx2XV4Y5NLXN0Ws4lgbCyWivttAlHh7ZDdcRonolbgpJdp4
dsHaePkOztS0iBKvUT8+Rnk1/6UoqiY9YY3RpzxJKRajCzYi19kZwliA8flB3o33Xt+SIIQL0Z3q
ibDIPi5pyiy+oxftEREcKH3HlxgKYKDCMsbTgeHEIqopQfbvUD0AhdqwRgxMaeC4S8fpn6CYPYtW
x/2a/rQ07Vsd+yJSV8jH3Q+suEWffUcoOnetzZDuVuy2xLQxpnTs93tEaUKgyzsi6clvWlG+d0ft
jfXJiX1Arbjr4ZsAeuKnMihy9yflGjcne0WdWvTbfBrLnvhUYQISIlZatsFU1C//hLxIfvlOZv1j
mBLwSWJY26sNY8jzBMGnA1ne+Yj8Pt4qHQG3gbPNyVnquV+6A15zhjp9iBx467ivhzqy7BmiDw/T
G8IWjjjfK4cH8xHl5nF5Aio6AKeB9R47tvOpQPxyFdVC6k7yx/7WcDzpXtXth24dE7q0aMNp8Crd
iGVNElfCxjMnz2tWolh0Rl2c68iZ29Npk/0UQJ2n832IIoU0ul4x2GScaKM1yoc6Uw7Z0s+HcwvT
I05hBJEu1bMI1+Bpfz7XXS7gUm8mv7/PZ/SJgysDI+sggvnM9vi+VP70uk24ubHCUXdMXEHRaRBo
+B7+mbDQCECNtRJZN/N2cpYZSHwwGCw/iAxsj1l0fwf+/sjedWYDe7i+2uVORrTbYgPqFlXIR5qb
0hYasB/0miYG3SQjLIFUX0aRCL57NJimVN1QeyqPhbgg8KhQyrUo+yynZBt2VcmfDvV+5CmdYRai
Bhf12hKrr8xe0cglA2+eU8vhJMoMAkAi+JD39tIuy+nO5V99YhPQCYrA3v20OJuvw3AWv1iU/Y5A
pIougakHakLY3TfIrQhbimIt0rHTXWJFy1VVSk8lTYGecq3mzd58yJgw8c+PXIQfaJWSQ7nUYQJo
CiMHYqLTeQGSK/CtySSfsCQgikRSV6WjH4CI6eJfyKBbw3xT7nRIgUGgSDYHSPkqnideEXynr+mx
oGMUjxxmQNlB7yOCe0pmyQCq3j6HlMYas8xTmxeLw5mOfdaCXmg4xD0T1MCxgl84bTx0c88FHuSa
08HTlqWwH7ZEe4DoYKJrVgWjZONMuBHIcbLB71bFITDx5Yp0cZgIUfk+p/P8qYCxOIdIczBtapKm
7xIwQV3eJgtB+sARhYfaA3UX1pb0eplEMpvjiC9lGKS/d0iYGpPhjNuA3C11EcsPF8pp8jcyX/1o
yRaN1axiN3mgM/mrd8CfPJQi5oHNgyNMVnG1HQE4vQjZf0rNBDrOdQtZinWH1RONxDX19H8weHjo
mF5Bx2lUirUK0mEuPYV20f9ih6/csLgq1Wx55B+EVm6KSj9+UQizmAb0nhDyVzuS1OtGOTIDrTaw
nbFHyaalQa4DqGwtKasiZx9u5uhkQ5I1MpPWYNW79IDZw/Qk7RHfCl5S7o85cl4FUxUxfEzfpTFX
nHYAimKtaouZfGPapw9vsohEK0pUozqL3mNhM8nDznBq5K07CTNtrSARoPRc6dqaDbpRj3l9AJa+
63gKJkKRTxwi0SDTZJwCFnNpIJxmYPJEfovEtrw8rVTVKluswaGJwUGYvIsl37CNgzoHbM+y6M9t
fUd050Y/Wt10lnMVI/ogL+JJCiZhazQUrwJ8ljF0KXqwVZKiECgZotqS4kdUAXtqGY1F7JZTtlpz
jNq/uB+QUbFQ8PLOT9/izCwtwkoIXsY62orQmWDFd/ovoVZwII+0pmkAfn0eXCiIZp4w7BHlVAWc
6eUdwzYW1OQ+Fxy7Q5IFSKIbTWDHus5G5PJQ6OUL3T0swqgAbIicUbArQRlZ64jHfJKav0dHX+mC
4Qrb7WVGLMhXiEykRqSEIAZjzp9lRhIY1mntHb3AbKT166CWbj/My5/lSUOuPxaeUvR6HzHNbhBe
mOPaTwfch/M/Usg4GdmjZjsMjiv8o9dV1JegnGqSiA9uukQ6uqv0ExMtHGW5Bss2NSe3GlHlyVGY
dDK5Tr4RqX0KJIRfYrGGTorD7EEUuLxKcsq06KbvKTx/JtOusHin5EjT0jjj7Z4HoIpWNZ5BffvV
M3rHrM+SAZvaPggoqB9k/bRLovPQAGchxlWcVVvgYb9Sv/MzbFhSIjV3ibIPsgLf1K41+xeCXQNa
ujYmpMpSlk2wQ3k2PpByEALNc7SaIqkRTEIihvED5dU257bidnVEcDK3dx/joXyXCqstzjMNLlpN
ZEHWF5sp52TKvKUp50jXn2r2sO9ohxYxECzIXrs/7GS/eOmEOX8JbljlEizA7X0d7I0Z6w+Uv1YT
PmNPVGdeDh7WJIFLP7OJ8vhCkqhRCCU5yS/eRR3kNS6HPKhHBX84JtSdzyUuDSxHHYh3hrJTiA8s
5Rsx5fyc9F7zbm5Y1hJeewnF6zH55ahK9owBID/n7haUNddcrS9s4IfyYHNaUTFKMnmKCVV6BtjV
RtrgYTVdhT0waypdfFVoL+TH5NOrj9N8vZta5Q2bHNSXDjf3DSyU9MID7JFmt+DwdzLAsoHwbhFe
I3njZ08HM9ZQ1GBZb0JDAuxicK5RoLO09GEc/p4XZOzTtGkV72y6g+e8ZFo1Nd0MUIPeD75bOspy
NM9xPsM/4tRmxl0SFeSkRMzVt8E3g3/Wm6BNJ47NhPHvSerV8/60eFPRQjBfjqjueBAzl3G3ul5S
mrW/aycCjpD6uLfzPVtoprA8sEPc7HH7JT+aGQT2MOknI4YF4WuNNH8Cn896Uw91NspiE53Ba2NP
aq3+OeymS+O5Gh10x37vklkZHNcOFTTeG3dcNbY/Rjk1KJGdjGGy+h2qZPkuYXNIgnJ/SAQ4D+Sb
NijhmT+VdQP+8/rhwQC/T+WBsA6LROkF9oio2XkQY+r15MjxzH+8c0yUbP54PJFJXcCNdL6YEUFP
UVC++23U46hkDAZCn7VSkc58vH2khKirxyQRFTJ1DboYxyYU9sXiT9LC1p8nXuuhGo0ZG2pJWYwX
5SzbW3tENzvEpHVfDuOZxy/HS4wKfXHIsULSc3dmrKKvpxIb+/xdVweWSzzybfcTasbTaMs1sKgZ
Bql48TX5i9NMP6TSjisQ7r8nRKTlxH8yJ+uBLDUdZdTCF4HsxcEH1FfTR2ZOkqZNPyretm9ag+o+
2ccR7hDBdHoxWuWfjyoo09LFkiRNNCSXVvF/nEB6ZYMMYuV1S4nCnQWVcBWE8jxr0e4L8WXhE9B2
Kunfko0RCvXjSL+4A5ghHfw4+Hw22lRn7f6w8DSLZOwlyHmTXNBfjvjse5JtXU9rIA8xs6UqmZZ1
YYGQ9G6QAtOVXvgoQ1xleT3eYTF/r7aDB7R+rJQTlGtGtEQ3f/6TuNZucF+IqnIc8iLeeFhSAMTz
VuZDLpjniteK4C99rWUUR3OZKHluVHXNaA1gfxiPm1yuyWZhyGGCzgL/aTbelyyH2RbZzBvcBaLT
rmJELwid6/hAEeCqhGZndiXTOprzalT3/S09QVI042J7Jqx3zzetC5CmtYn4T8ppeq0IcpJvFvvr
zhKGuHOLbXeTFdeI+Z9Qq/2jf9eTfR31HewE6IWxFQUZHhkIk29hXsxaZIXtEuWf+Z5TJ4/lP4wq
coAmkgMwPIOameTBeOAZzQwhT9NXMPb8g4Oo3z/xPvzLV6VHwVcyJdW2ZIkVIV4Kl+vnxPVvXmSC
WRP/kHRtz6U1nidku3Syw58lAARkQDWsYmVMRF8tzDWJYwAbasTS2opz/ug2VJTT2VXEqGn870gA
6VzB2Og6nJ2MUPMG94Y/dVDvPafOSJuZIcRDEuivh74OJf1Lo869WPGjEOTIepNCPl7B29pt1FUV
gaPv4SFrgKGyvBcKBbpEpH2q9u9ETxM/bgZiCMUwKaJpPrRYreJiimmVaqV4BremCJFJ/7ylvWX4
Vh5GmQcJevLsxd37peJ0JXm3seb64A1Nyv+9Dlw42Y0um5WedRwgnQnnw4KIi8zlhamihf78Ucnh
K2fgZrbEiolBRwLpeHt3EUOqCZ3x7HLMlXRTv1bZy0zgVo157CubcHUEZpEiuZLmBrCbdhxHdBe2
O/+RTAoL2bho/9VQGlqqQI44B/LFvo6tKZoFml5YvQlBKcE9OWq205jH/ab4aUSsD0MGqrZwF0dm
dq1dN8xs88MJNC9prXozD9vBg/B3atFEePNjEN+HDkjeZ86yfUjRDdvnyJK6GsZtws4/bR4JNeYc
xqSnKB5R3/2w2woHaR9Dge8v3A9EPxwxPFYuel3yykfl6UCKQD1vdDFuuCYtNslOdJRPoOXxjI2d
iaogy6YYqU7GzfzBL+h6p444p9Zj43jsQhyT/geNOOqVr4/7wi3Q/wQutinC0keJqgSsIjyPyKSV
TsyTxEIukBl1C3rYzxYAvqezLP8Yyb7KcKRKzK4A8IjjGn/OIiYXvXsAJI/O9OOKWZDVSbogbk4V
KdAJZvcCgLnQlGbWqvUrKsVQ8bw3E9DoVaqPdIdWicDTKuubzr15e4Neo8m5seEAld56yBN/xTz9
ennAkdJFlOGdc8tdzJXJNRXEDKtSt5AL/vaMIDf+h9Ggf8IxMD58Y6na9bTG3pKan/yQJPrOBGH8
PqUxkJlA1CQryxKIXt0vTRLR2K3m3V2tPWKGLzTejRwG5ix2QYk9tkbcPMOiYE3bnH9vietnn0Ax
TANTfmiGE4hrNh/6n5ypDbSjQ7pcbadaB/yDz2yYlqhNuY8ZTgD2LmiZYY+KP72SVmIRMm/qRToo
L/Ifzt156v+gfEer/B1ifnxGWBe0PZ5441O7fYfXZOVsc/VJex3jygLvvIaafFZVxTN/yeO8ezkx
9fJ+EfjafN+SPJJLs51+IhwiYol3eACb3/19MwmZGxH+qTqFHklvjOUzQClL+wUiHVoANShVrjvW
89LwlcS5GZBBO/sX1CxAHI8XeEHwePC25mZ6ttxHWOydObpEj5c04hFPr5+XQeqmKr+QSXK6XskO
a4JOeHnpNIBgTOZHqouHKTLY1HAwqpLaWBhYKag9HUdPC6R3jwST8mE0nNNtVY9UciCCZ9IZ38VX
Onpybe5xtiSpmB6zFbcvxSHoukP6sK6qehHD6M8CoOKIivtW7KsRWWJHD9vHQjV/XWa2lKxhBm7C
TAHMmPjOSpBVN4LBDHqqFPafjmWTxZ5HHvemCt163eIdweC67hCJByRMpyTLVafN1TLwVZ668LWs
oOAEZguoqX/PnIHf5FrGR/IqOq/3j+Nnik4m4uGSORUHyfY+HCedqvhC21ba/QA0gPenbaVY1kKA
1jkZh2SmIc6gjUIF0ETeL6fsJEKe9OSv041oJf2dfT2UvgwjYgxXX/GFS+F/K4cU4Tn6nIazLf0G
+B/LkPI3bfELZqOO0dnp6+ajLStZTSEJ6SJySFvBDCfteY+uukY5X/ShnxLLLIAuiaZFHHT/UCeq
qEPc9h7MS5YjGaAa16wIkSxY9b+SSJw764Mv1PcoU64IZILHFSiiEtvKYn27cKi+yqzeAh2BCW5o
j/BI3hygN6JiuOv7bdnRRoZqZJAUf3xNoPVhNjl3et/TKp6vWY8TDkcAtikh43gYOXWl68MCeo+7
EHsUxkEI4uEiS1sFYqd/UxfM5b4J7v4EYNXNkpx+qGAVNN+wGfMFidPfPGnipaEyKKcszP+gdbDQ
WC+0bNtZ8Z44LnC+LZzYfcY4YtJ30vEya9ic7jkNwxwvKGnI5fPSzPgQNNVCiAhOognWOlHU5RcJ
L+nXzqzfWKjr+/eAqVU3meJedB5tD2oNoGYokH0fZwoIxLsPadn0y4J+8gKWrmDCwpCiMSPENZe9
ya+lmi5BhLDT3ttyaBOIl6XdM/TWGtWvSQcRhIywjAVf3UF7hdV5vmdymGNmP2zqzd49sEdl43O6
4tpW+c7J2dT1Pf4+8D26alDrdbmxmVYweoMy2IZ9dCi24GAcCX6ZVO7C7AyGG29TaqYofGaypIrf
0PvIVYIPb0FKfpT1k4A96n4FJ+RAzfIPjwplo5xt4fo4kKofHuVA6QkUFsoJZZp0PcPnhiojvONA
uvO5l/Y3sn8HqJpLBAB9SV03gpuhwisGDdcldQBxnU2maq8BevcmA3ombXJ1e6m26aGFIX5ti9AY
WrGPWTRF8HW90kWb2qBths9N/WzRSFE2fBj4C2o2aJRtcLoIKxGlvHPlfbcNQSG6IlxJ2DQCG0kc
pFM2iFX+J/XW0r0SUJ1adjXx3teIHKKT2FWfMsoM3CN+6NOO30XkkCtwYZShcSVw7ndrcmRwcfNY
JWL265PZmqnSoXXV0+v8RDz6hEzJS6grK9rtkNLKgYEt0OPiedVEKWyZuIEb23HeNAYahS07YoHD
E21Pd5DmPLQ+Q1iNCqZ9JZl0PILvuKX8S34jlPNj2R85tZzloxA+QjnFoq4+Cftvqyltq4Agx+69
lul6xvyqBQnDy4UNW4UQJRfRX/c6bHrwT67rtEArr8bhpaHCx8Nsuo7rFV+7HkwjrHugvQmmWTKE
dLcpyto7sRl7bqIA0+aaHIU5PMHqSdQlOVBI8G+lVVT1h7EskwlUwhIQtj3Dp3DyDKfmsPVJOlQc
MmM+A7fkDMns2Byc4hmO8RXuPnbxnC9O8SBtG+dou+eiB+xBgJbmZJu4dW4ezPRGMtqgyomhLZX8
x2HuCmPKcugmtpkMharRhvGxU4doqGeJE+j9xqOiUci2ulM=
`pragma protect end_protected

// 
