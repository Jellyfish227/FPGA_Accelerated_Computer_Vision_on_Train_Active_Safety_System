/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3104)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnKXH8K7XVxfmuTx9fAi8IDzAobQvovQq1S4XhIbEOaYT9MdiNh0mBnGP
vjqo4SScQtJ2bzDIAmTLjat2G/s3K++IN0IDWF4SZtQ77NlzoDJz4trkHlrDRcO7LHp6uyt+w4Ok
sRamt2aXPaRoUDSrESuZOmIqCbVOwGtLFuuSyYN0TOjIcfH3VpLg0pYT3JbbJO+tbPeprJF8xRRS
qeUnr2DDGDBZA9fg6Yy3/ILC9nUZtNkQj1SbLKGVbIDqgA1dL9gTiaqVut1i4YWSAD7t9YTnpbTv
+lGrRmqJaKQ9arpB055CoogtiDvQ1n+wslr1t+jyuFR4saYDiDosqMliXsBwSLx6yQ3ro63H1HjD
p/reNYCjDH4FFWnso1odM7M3Y92LE9EfMx0dI/iJD4/chSZWIYQtwH2tBhq9m4HcMGX/By6742x0
VKWZkIwEVXoLwl9ZCxhqdq78vhlw7svEFH5JnHB4crGsObjqrc4ULKy6I1vK5axfxzJBFnpyE9IS
2VsO4TOGmu/XjCWJ29OmCxty0oe5qOMTjfikWKHleH+V6gpiocws6lq5m+Z8YnqfPfrFqnjiosWY
5HItG9fAujo3QQV7eDx6p7cmKDNsqyuTIih6sThJrtjDWMJcE2U7ZxN/lhe315YFBlWOj3plvIfR
1yNU/5ryFyzvLgWeDqO551501BUGvOTupS4x9eZK6iz8BMC2r59ipS/F5Lv/CJuGplFqsFEtZRy6
/qe/RFnrV5Vokc7xUOGoKt1VZYzbBbZhP8QT1POaB60nYmfjA/KCxhEfuAGF05EZGXt9s5KD3ItA
ntAILMP1dfaQyz9PguZwNZ+W+K8Yl3hf+MGCJq5wiciU0rIrpka59t5Q0IWOrZByRc5zpY97vnNa
MS8ur6FlaOuvZiK/3awRbUNC1O+Mf7wnBvhe2/BNC7ahSZQhZgfZCmevfjoXBZwFbevr2OzbmqiP
Du1D8Zp+EBdB51ZFyCHCXpbmBgRnI5KrzmNLZz/MPDbrPBrWpqniorG5m7K0tYRovO4AoRIbmLzl
p+pnuYVS/XuPir6FthhlUHJ7DmTkMTbLpCLumScSu+Vwx2GeG8dYUAZVWIRY5xTsRvx81vT0IUAw
FBM9P5FGDtEsvuZeNHpRBNHuk0HBVxAAoi3h/WrVsPW7W2aM/RZJXOb701CMdx0+RCFygR7FnYIA
eU21zcKIpUeN7FI9gijxJBGqi3+mzh+HY9Z0FDZTvFYkHLEGfuZXFxuxif7H1dCWViZoSCKBrOHU
6x9Z0Lp6NLuMGHqFOkk4/2xtzkSI5PuloepJqZkHyfx2+0QtWNK/D3D3N2mxK7UDX7UpBOcTjWI1
S5GsPFbrbD0lLET2gG3JUy4rO2byu6VxhpptFdMgIMv1M5WBUlxcZq3Mp4WdzR8QC+p5hBllb1PQ
fk466fNAp5F7RGv4qZL4DR839SU8rKMnJBO7uIzjeFTRSb+SzQaEosl+N6WoGIi4JcSzGE0GoRPS
VhmxEypgGoFIrGkDlStM+JGD0w5/kZ3t/X9ili9HXdi4vkPtSon7rVUdwXZOzXhGMp2s50n7QvCK
y7BfcGHmHq9VOAv+8wriDI+Ml/i/DEf5tbyinrXLUHyJLgNIVInA5lIq+AxsAxg6gWuMB36ALC/w
jPMYFFycHlrTDbpx/nXHrbS3kqyQ293E7prngIZTZJTjlM/8RfU5Rd9a9oNSkkmIcn63lQKv5i1W
qjFO2uu/Rxo6U8y3RXTynWchXuPWCJvLy9Q1UgldZDTW3B4j8auMwHp7NwJau16f8E0NJj7ZEZIl
PlLB65MZg+b3GvhS7LgEzGGKyWvVJqxDclx8Zy1mk8wU+cVXR2ETCZhggoM3ue5kk/WxIEcx2Do2
Sj5UeAEX47YtrYq749MpVy8eNmm87Dy1R1VQJBO5ElHuSyn0bRS81/P5NBm/mbzmb2wljzvHfraH
W73H8EoxObCmU/8gTUXQkqqtFVpN5uxESwZTr05+rSVsXc3UgeFYmw+vH+tQ5BPl/QTv65w3+HLC
2C2pz92nsq67BjH3PRMhvvYFn4N5p8n5x+ofAQ7GmeB5SNL0+43CiShVZXnX8DEedOEEcGLaZDRY
tQJsSjNYHbbl15eYsXhOy9S9la5ITU1lUsjNGT7sHWIFrOwHXozfEMjN6qL/DaS3KPwc9xa5GnWC
jjDZDrwxpKfdgZLcJ3AK98pRzVe5Qdp37nMJDg8K+1rztZucT/YnvtZaUWrt3EHO0BKG3wchiuKm
L9t/0VVU7DGzD69Mf1jnG7ysR5zQwE+pD676A1tc1wiLXDcNJxB0MTbDMkAKtuwIMqZ7SK1eABg6
ic+GHE3kyfJqtOaxYmA+AsX1o9Ef+Yt25ONIp9ARVKBzHgcsn3/u7avruZC5odj5un8OwCjAhAXq
8TWcV6PIK8743nosZoFYk3CwLtkrUANjPApqCB8k17YJ63gtEJJpGEbpc253hPw6GncCLG5wpH8h
6uPf5OzGzABw1KSqLsDQOynYXTl/6ctNOblmN9bxT09Zy0vincO+NMQkTGS1qajtY6NaRw3/4Of8
jFSIPAg4cq2kiWKCyElJWHuK5F0uweyaqTJQiqxrHiYf0uEv4Ta2+zsEiJZfRq5xy5ISrX8JqjVw
/+yOXwC/lGzdKfIxVaHBtGM9zKup+E4q6+8WugoW/UUjy4sEmd49PdEv3m5xCvu/m6bqeZI9be+W
Y2OA4VufYMwwwAez5781agVvl4V7Vq/DqQCCEZdiSaPKzYV6Gw8xvLoVpuD8G69YD+/3Hq9Z05c2
+/Y7O2Vy438u2zQsQ4nqZ302bLP57u6sB92FdiQVzqlBMA6eWhuUQXfceL3VC0fJKt4tSwJvi4Tt
DXfiNronLal1LGeeeSn76a6SCqcx5EZ2fbXV+4npS1bLi7YE2JnT3Lb4BS9WeV1Zmxf1YMIOFemJ
9/PHKGWKyFenOtcS8MsVjtw8cYWbdJsWZAh2rnR0s4Zngl59S/Wu5mg9pXAs4G0O/4bZD3rO51Tu
MnWWXTo57T9w3JDCT1XMME6cJxw4i/Gq30TPvhnXgzW/lEjWF03JIb2p5hm6n4vtdNy+/1gUoy9Y
PUsxmaERKCBAguAuSv7gqLjLDPE4eIiZADsuP/1XVcNtLULqhao6+yS3rOemUwlo/3+/WPCF1/5l
jHtfk1O3mEy4REj+I9Rp18pNLS7K0gK/2ihZhnD8d03cqqXYh5asvt2HcC+8HOi1C/ZuWml9ipd7
W1yfNfn1fKYF4smmH+s2o+Weaf6AXODWOy2+bluJ6alHoBv9IV0Fs8PdqP3YrzsrVhnh/uKzxW2Y
qXSuRFg0E2ZC4SoDM+uXJaWvR5itqW4ImdRcLcZwOtPkiPdFFgldZKCM9dt9i7RfdiJY2pAmRyIz
5wwNetuZahwokeO51QjaYFzlSwckh3gx+yurzVMQvNsWKlMCZS45/1swZNSTDPsWaxf3hgKeT4Wv
hWo1PJXUuh9rcbF4GjELqR4r8gTyW9t6lTyas+F3q7tGYUFOPh0gyUlqvpZ8KE5Zzb7ZWLOoWfwF
pnqKzKhD9BE9/xEM7w9dClSfTlywZ2qC6cguTOWa5Wl2k8QvOUWdlY9I1UdYKTQS/9+3CZM0wVU/
FGWmSbFyBuGbDmk0SSj47m41IObv5TZUkMjuiGJO9QCXjtbIUhB5WBOfuJjWGkeDknGUnMVFndBp
93jq6syk+Lrs8/WAXkwFx1QTvqMTEP8Nq/yAOy9UPU5jHxCqf7xcxhxv0Gyy4+fhojJ5dfUbDpCB
dtk0wd04e4RF5XlrjsCCK8AjCel99DBlTZhiIs5OAeQ7W0BwKirGUzDjqtilGAQTpRZpMeI7FpUK
7z5Jqzk09voRwlprn+F2/atyuG8aDmJqsCSZwY3NiIjQvkxYAsjWJJFF63N8qsIrD2PMLbYFHQLU
a8WaxaiQ3LuTbsXyvdBDTiGEhJeZZjGEMLlyYC8LZ7ZSD6TYIqyJmUYf5UtT3REiCGXelf4OHUFw
exY17rZAa1aj729V5734JZTo/eMZh076u0adSuBGGDb4eqB5VKYJJeis/blOSz0thMFjhzlHYZcn
0dSnv8wqQ+P7MAN+q22EfTHnlLp8kfMJucw=
`pragma protect end_protected

// 
