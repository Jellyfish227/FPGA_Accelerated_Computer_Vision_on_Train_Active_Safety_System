/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
FA2iPyPB/2tpztCLxyaqpOqdYWzKk8FkR3dpvX92DJoJOYQ9Qc0Nucd2MFWr7H1/txXVOsHKujyl
umXt7y7/ECsfh3TH7FKmx8Q8ND425QPPioMfmAV+2AzyFJyb7fFOjakIOmAszEoXpXE/g9ssblhS
pfdRFgjSafTue+UvztGSTJFfzVQXZMNIrrzjH5rQ0Ao2dAS7SdPoRYKOOdDUZ8NCMp47RoRWyEcz
0hsW1G8HyMXRK9cinGAcQPqIoO5cb+JhKU0J/ePfJuhND+UKVMoLKQ7dp0SxMuqEFU4hOtJHXHet
vYzXNFhHLliR79jLoW44AGt00xN6HJLmt2b9zA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="SowHfWTRpH/Eq/YbabpQJUEqKOBSTyQqcnpNEvDZDmI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1236672)
`pragma protect data_block
RRZG7MjqAe1rc7xfGwypnOflgQFnrN9anhp8Z9g/DPaEgJwT3ZaYPNV6WQ+vLRPZrttbNotAskB2
FD26A+7zT016s/gst+FQEtlz2vnwCRKds0kFJMcH20olPNiGa51CFAtaqhTOK6/M7AgQ9shbYmrD
aWNA0XU6oT8LPYi4Y2YGiBE79Az8OIdk3qltF99K6AaLMC/Sw12EYvtPaCt+FlMmgTZ5FxJ/a1u7
TDdbRp3isoQJ8sR2ddJekkFprjEmqxnc0Mb6FHT3Myh652vzEVRTnqEy6X3Swgh5fC++k9Njy6+G
sBVlY6h8vKXYaEoiLwm9dOTpml+Jrs2a76OBaStRhm3KYvwmuOAqMABoidvGMbC6R2x8qZhlER4B
R/p5mEpnryk+zWCiVwY8h32/ivJ6+ma5Cz3rtnpD+Vva0qWo6CNJDPS8pFgo8V2LNHi/sXT+IRMG
5zXPXY3c/6C2x7f7DPyz+2pKrW3UG7d/zI9EBPJkTttx1aInT+avkwDKIr3Nj74vmxrAHBYfCSqB
9AXsKd/kQ105gntNUIi0qyEtxbDD8jh+ACIQMFR3vaIUTtXsdFUDhnb3RvarqtFJEJDAQ1mU90iA
pz+CSZHVUrjyHYaVAC+85CLsyABtL+qIlJ5zwMcmrqYaTYD9cz/FRVOXnbCg21trFX/5bYtKlYSY
lqb0pW8z/hcrUT8xzj+w9zkIObt79IeMVm0jQFhn32twbfrmn3nZvjpJupVD+pqTaIFjrSZS0BJA
QRZggp9yKZcNqxKd2YfOOF1dzEDwNlYocdQZbqI9/YKoN8PQdLvB1KVx7awfXfLccXbIU2cm6dQO
dQ83l01UNouB9ok6SBuunM+XszQrT7smYHo4QNHDC7RxLXH1Jf0CmvHlgHkNgTzv6tTWvn2EweFD
djjoAr+wpcNSJ2+4kRuRcQIkSG6pBvMPtz85Ql1An8o86qRjWMtBSj62q8BNiTeasaiqnHSZgcfa
oBCI/rvw5tXEKaHWSze6enR6dSJOVkt7rmTAb6Pi4CE9t5eIo0tXEldIEuXuWFtYmnMWbyA/JJuC
xKNveSzsuwDTpjlRyMILQ2UrPX3uuQy7/S7tccxlnwNhbfkWGGLZlttutG2Sxtzv2tk8OjENdWgO
wV7smT2YQQXSUgQkNBi58guUQqJZ21cAys/QEWxjeyzF+uIjPp6o9OJQ0F4CWyBlIH3DuaxOvB6f
0QmQA9rF2lIKIy5mNZWcC2MR3GtZ4RQwlElpFa78YAi0hIbQY+d+TFX7fBhOm4xWOtwAZw4+tDdV
0yd1aLHTYMEnHsypF+fFem+D0aCBxiCN1jH4dQKgZo81c0MS4z0qGYnQFWn6eSXEVrhkB9ilCJu7
kcrQbJOOywlCf8d6eP2mWoaN5qAd19BmLfmKJ+b2Xa3Oh3+jI7nHIsR+buu8iBqqPHFWE8Pi72R5
/B2vmPrlRimG4Unm9ba8mzMINLv3EiUR3ohDogcI+UioXBh2cs1ACkLlE4kH/rRh7ATHBJMJvJsz
PbJRPk3oCMsjj57meL4u5xHp9WWMrQ2ybJYgqLGQ9Jjcsj8IX1JTQd/5BYv/N1wT+JCVQmNVIpTn
XcJz0K1mbYMxh5+w3EjWv4ghGLVwumTsbKuOPes0/YQyJdRrld9xIKF2QzrrnzfaQ9gVxy+XZKQJ
qw1DXIVapSSW62c1hLsHf0ESwbeFqygrIoDL/V5lqfj/ma/rv/FsmWboT79pE4hIrupE6jmLqBml
oOj0IwroC47eoDsdzKnunIe99o8vcI81BgOZC6HMEACT9k5BRACIdDqf8RjD5C3y2zogOZxN7LAQ
dcissMkvl/XrQXX5t1DlfbbZekmGfjvE6SRdgMVXOlDa4CGiy7dsejG8o9w0/2+4MkE8zi5HmItZ
2r8msiJEYk0zxxH3xpZpxrEZbLuYpuMIK6ge94A1JsGGrBeulMVJHljwcBRQ0OvV/vgPHOW7Wd16
pDPAbq9f0j3sa8noUVnblMpHFf4lOawaePNirYqxfnEzskUrUt/m1Jqp7tyaQhY+L68MIr8wDkVa
/hJi7BxBOA/22d0TluUcyby19pSbsbxiDgri8JGyiKjc/dm7Q08fJPPei/WarF8KDKwx9W+uEJpj
F1NJjSt01/EII60B/fgAhxpM5mgHQOVeFSbX5JGMgqJNFfyVvUHeOHkQbHJU8OmXfpllpkFsNm3W
uLvMDfzBI8vP8GHorNOGJmG6DpvfjPlxH9GlhydIiXrmK27xCseHSHMpiSL9hwdqfvRFdq5nzCDT
6oeEVVR9ALjfTatGjthYKpmlGFBe1kTMI+02KMZeB1VnKMO0VL9hIO1PgVWrlKBfu6dx7PEzgKQM
bHm23bdkxZnzCZ5YujT+Orx9hlpLZdw/Wel2AtNvMc0uImTdBzf/kvCo1l0ncpd5+Qu9xQ+W+h5r
vwbEPXWcUFv25R0H6caJAneMteZEVL7nHIAT8vxqZrylnDV6e7VpyFsFL7fa3hmqjeJMNIgejni/
U6H38BYQzxp5R8IWpSzN2LRDhvm9Dps8xV+6uMZCNHNvzCVZHPuccELa8JrsopTq/SRdCWNXHWav
AAvSx4KgJg7EmRBG+IhrQRspWEC0rEpV8SMwFLVpkdilIsVChVHAidBHN7tdCScygD+fyjnlIodn
ZCbH9iAHJLVHUlD5yvEXhz865zX1EncJEf1h0RWB3KEvpCUwNuV1wfHhsqKWRqJ4OEzJq/15bjT2
rdzKWw5Hxh8dKuSg4gUwpVwrVCPup1xeAhpHaDhKxUfhRW7+ZKia/2fxCAXs/cbUoZDdzVCa3hQX
B6AsybYS5Teede9+udMRHQPPCxroPYJb72yV+nnyuwWUcQyGh0HtACwG37XK+QW7uAGpqxq1fzqR
ze3dQGDfuxriyY4OairANSmMyhOW4/83oHP05NVBYdyuwFy1OvP8Cb5N0dJFcsSkTjRjgOobzGFu
l8CajwupJSfhHpUOtWbKIp8xkT0+rTawrLHTX1uKoxPPU/nih6DUuLqVlyoWxZKkMR+zUrVtrUxY
5i6DNjo1Lt7VPLASebbj+SZQw/4R10ZPm6pFdWWJIdalo5trB5SfdSxZcMj/VayBqRX/qB5CHTqm
nkioBVmdnbc404CVUyJuODdrxDwuqju/wqKdAeD0a7Z4XAO/40Oj1OJ9kt5tNXNS9g7wixS/L/X0
8PSxhVtx5sQGff9szmT9xFvW3lLXIJZ+ZspNf2b/iWBKF7CIO+5niINn5DXSHrIP/6GI3EZWIG2/
X3BS0LRwS/VG8FC1jBrnzutvotMtvDA3tbEWrbCkGdUzHrmNW4BTFIYL7Q9gu6XSp7a4gCzuUlQP
cyCqggRwiXBchRtA03KHaSqLkIrUizY0S6Wyk+WoHUFhrbiDuh86NGgO6LiTJX2vfPLqFsWwWmlF
Y4L7Dl1yo7b4I3/+dac/MEM/KVagTKZY5iQtsV2ak2LOdL4jaCj4mnWe8LdyX7Ui8xB8b2DxcODQ
XS58xMCI9NSzRkpxenCLoa4iXqE61QKErH0U3LbmJldSnuFamGKVxfBrXvC0Jp5m2wCPptbhah7Q
VQPMksQJmRYjzmdA839miXbrwutVYTcUvx3fGAHaRKKx83d2UWaBvgHmLhPK8QRa0VbeGRLWPp2B
UHtiSaVURSNDc06YGM5zoUwDs3W6EUy3DTKGb9rV7C85V4B1JaRl1sYFGYyLYppZvHm8D5mwiMnA
cZ4QdVTriMfpdU2kby8YdJtJAYwFFwtsuy0/AQikZGRqcv8yrNTymFrCGcbTTBnHNGoOsr5dT6Vc
Id3G2sWu2U25FE0ec2Rrn5qUpW9ANkDsCtmPy46IOGC35wWDJwCCsKB+BO/JSMypPVNr/GK8cWAA
oPFlyqHNTZRSRVV1WgwGltypP6LYAuy0wn1kpfYpojxYQYNWcKtIEOwzdJPfvnb6gy/5fjtw0dm+
5BgO2mpxvbIF0Dy3jpjF/D6Hr0p63JpA5c2hfh5F/whqT3gofIEN5GcLF04f148J8iyK87YFCU00
O4wrn62EPn/Ofsy/nPfGggWp/qAhqgtlbs+JJc7Ijh71efL223zVwUA9VNEp63amkWj6vNLBDV/B
XqieWWHNB6BzF8hm+28heIZqsIC66Gg+skEUp8I5R0yOSVNqoI8NR8cGfwYJ+pAf4gIvmCU/Yyhg
FluWr7VGC6dHFHVD/+AS8CatzQWqxBYN/EcFOa84ZszMb3N2I1kQEe6UbxAU9ZDGn7138ggb/41o
vAg3EfbTFaSXlLrGY+eQq1KqSP09R2fJztCYuTmg/niUw1904ySNMC/FBSv5BlVKckygvDZa8Kss
qNmkI9MGDfMXHT42deHpDp+yVqmtD7nWRL3YqRvYY38EdAtstJOT9UOx650hYhJ3bVGLYCuMYKeL
WbUpu/YBTSPHXQ3WCNq8pJG2JSgqAFvHgO//G9D5AAEjYg/Ji+8UOD60o5qjbQg2XRj3Gvn89E3z
eIzDrM2JkFd/N4J6hnOuNf8VcUkD/mjpF4S2cDMS4pMGF3H6QePPNbKgCoKFcjRGtoWkuoOB7WFm
rNAiJAmS+Ad603zxcNRiH8g8AFlH8XNyeMMGnQPULN6zFml6/d1dYV5qSAY6xE0jzuZisMOP114A
jlrd5ics6eaSiEcClxyi//YwMwkUrFjGfJLR84LpbARvCqJTYoEbKIOhr+Li0LJMb2zPq11pyjFt
uQvSA0kCKD0NfYJq51eWWE6REdzI/9Kc40JXPKORK0LpBHiQOtjxJRDL3J94EuiDc+jJzBMT7jNc
LBXqQnSfe0b9jL5lu/z7GPp969i8x35LOXbH7suG1vV6Wm7ZJwYKZu25agsDoPEQRnDy2LSpWzfI
fyRQc/pm6vZPiidn1FdgD2lDjT1NtcvRyDLk0s4B+F6VYuBRiChKf1j01GDFLK4c3QW3fOOfqS6Z
2Sb7ZDhxf9pGU8Q8qH6ttabt5U9CSAXH0VZOmK7BCl8/Fm0KmQjpP43uadLQ+wQPO6bx0cmuz4bM
np4LQl0HXjuk/oXQ0eInMQBL1nd7uVtOWLWVOZAxreePh1CLCMAg0gHsQLlA1zgurDLCn6NOk9bQ
pnvqoQb6iG8C+SNEvnG7vwM7QveLUCIa2sjSq3vCfI2yyvvzZo/6MlPo6OJuQ48Jdv2J5a6V8sYP
hLOi/87CH94361g6IUXouci9nhDfgcY1lmjBlaDLwDoHEOWCaK8o8+I/T5x5KjmwSIvdjlA+u2wf
ooV1EMKEXnpETsW7RiSRqHFoJ7TYCENrboDEIpbQD6AgU8/AevX+wKsSvKj7Fq5PcR+O0ABjeP3m
fViMBfSsGEuLCIAWoK0KX/L3lhrTQlY+yUCe8awb2K1eoCOCVM85EnPSQ163feinTOjVukNk8Tl6
HBj66v+GrOG29rUAwCJ2XFeWiVeUIb4IbkcPbsZB0U3PT4abQxPKqV/MGdH3kik6QurEEMzgpcqg
acl5Gr9+r/qQOEXmGROkHxdudBRW9vjbAaJz6HberVIICkxl5nVPPEn1buwZm94+JSouFddB1mct
kaXpdsu5lVve+8LWOoY9emDYs9pURBsXFoYkHC6oHqDM6Uam11P08HqTzH8wQB7kqSf9EOHnaITq
/qGyhCb+RalHYGdlFdN4zmLyE8DWpJOdyl26l4izSZ7m/ffdewcoU+kx7ZkyIRDPRBAQNnTmg4vH
y0lZehiXcc6rYXGXcgnpJcvABaUWB0bhTE9wEcktVjySHaLAr7qiTeJA3ytlYNuwA9HowS4RS2AD
qYqtd8W+sRbuKv8fdxT1lr0h7vW5wGlpND6Wh2NhUTukNxCUl1f1tJ8tPVsZSB6xKLZE5cPG8PRy
ejUur0h1p8AehJMO8Lt9IxkHlHXGCAYw/znecMf3N9jqx4FoPD8i4x207vDgIfRpGeXwNkHalBkr
T2A8YqmPIlOsomYcV49ABviPF1jZ2zetO5ATfUogdmgxMsh60MSI3VPPvGg1F4lZ1Tbpu0/pAKQL
UToOmx1Irw0YwRhzbC9LuRTHVUigWUXJE9Eivms7MRey5CV+Z1C7WS7nzSjtuMnKqmZ0x5UxQWB4
9ZBe0KC8l3G3mkLcQV7P9JWzMXXBrFN/3xWWhbTBvKGQVJgUxDH51vUWiHe1rd7z5/0/gOp7WBZh
2M4j32WRYcVEAxhOyiCt10AgWziOQWDtKzF1q9CoKmiaION5er5X9CwVn/6lP7UekLfwB64eb3r1
ksjbZEv6E9Xn8gpclox5VeyE9C/oBhk9g7fL/bS6b7DD1hgt81aoQRtwY+gu6uEzH+vZmSJuUqor
cMrnWFNxUD9NkNIW/oxpCPpkuGkDljRc7TNMXowrB2JSjRe0Z2XkHMx7ThuHduKg9FwF5TDRt5mY
i1c+XwiK2bRizC1EtOPCpMklhnooxCAtk0LbBe7qNd58YzJeyb7IPn2rPHCCaFHvZtQgLKxnU89i
6lxqGFPfi92ZZjHOMyzzkqPoIwZj+POAD7QLCtBrU8g5g7Hsu8xoQ50NXq71vy6SkGMnpZ5tlrgs
lk5dU9KEpkwnz8lDknnYaKqPJWyZkYZasy/jBX3V79/DLLEtLYq6vzVts/TH/19+X6kwiSQ36nqd
mpLgCZduNHdvZeMEpZKboXKxLheiQdRtLg6mG3g+qsNepyc8yvt9R0HRNn89RJj2Gz/bs42bfE+s
0ZCsP2xNBoqEhiygfPqLoPrIXsSMMV3aC4OZ6vOKzBiJSmI80MH0pP4upH/BePMvuGh/RfWqX6MM
vSoVtrIuV8k2eyIC7SkfgQbU1dQXx5uA/Dyw3CqyE/Ela5O1Y/BfoX6OLoHQvN7cphwDztUg/Nmy
4KZakJxFkjYqwx7uvixSUDqWcN6gjMwmVfx2yaaQs8m1/Ga2GKCOO7IZC7lyeVTnPEGfHK9TMid8
WJ1H0NUkwBeOkFJDFupQEzE2ONn2wgQPz/lxAEMo6fVMvG8sSzKyGXpNqD2N7Zb3hHi9ktS/0VAb
hbwc32mUucIlUm2ILgHEihNlQUJKC2+C7M1qXOEFf2Di8AiICktaBrtre/mj+c23PmKHUmI3OVrd
Z/tWGuVYxk6dpT8KJEOE46yeVBVRjphcuDxtkfWd1sx1APcYNZvtSDVdVhkUoQBiK3n6hOeu6+P3
d4Gtadr6pLa52K/aSsFtzrQL6Iv5yZecIvoJm4Zq7iESbSNgkeZIHWBW2pA2Z9pujMhP6EPHAp0p
PLktFhmscfEm9T14jr2H1UyvTEM4hf4tiYp7E8ELRjMNgmH0jSx8WVtmMbKeiShmzkWEdLMz2XGz
D0Opo/EZh6wkr/YZxdiN3AThAXsROtTPOEAfVUVg/J6dtkDIZqsAZ6Vv2rJGBrsT1ohPHX/Mh/HG
oBxvbET11qy4VQ5I1jMSeCRc7V9eAhnROehnqRKcI06y8xP87adOAjUu8uurkwHCDpvpws/l6alI
36NKxJJ21/O0Aa/6DPFiiGn53X48Pahl4yvlLIlbkIRZUbTIr4FOxMKoAo45qGo0u3EpMXWU3I4B
hegmbyNl+ImfTwbiXkq2QHiCoHDvi+1TmgWkqN978M7etDibe7eDOz064CxIb3euz3ShKXBymnn5
TfZDI0//SYjmV+E0nYb3aCWST45nFLENMMyJQfZrFArmZFjDRPVpcVRael0zEym2wk4kMpMBoyli
c5BQ4Ga5fzZOJD1A0O4szE1d4mwyaZYmIajvaF9wQmApNTO0HHtXIx2Nv6k7qnZSBtPR2BozQ7/k
O3AEOIg+4jsztEWQaWr8f4Hl0h0oSLOQVgieFmW8F8jb2nu3VHBUQGvQ8sOvHSH9zYJml6GzeY1C
OTpURQq/IhHeZL3CgAc7h0Cwg1zxBINGxpKYScBfBDV6s9ksNE1BOkISwfLz20waR1ic2BaTtMHD
OInNrtA/YOzsrjtamZosmcJbFjpoM+ayp5MbKPYhIomse316jhBqFWZNsNbVVV3TSVYfftLk7xJI
xLDh9Ie+gsDf3F7YauWYJMYTCSQHNSvr3TvADVQ14sLk17MU4yZEZTPHfRKvTFF2scm/JbMb2r+K
z54bbwFNbZXN0UJETxgnJPpbCLNoVb0vkCkvbwumSN0cYeoFFpTr2qE+DvcLh1cks+hEom/FhWmA
EcdacLTEcj0XBMjbs/ZSuOqosyiwmquvqAKR5NvYcM3YXd/lb4w+nR/EK7doiJ//ogZFldLNlI8r
H28Z5GCkF4meEQkPGGmGHFvyH/sEIAwl9nkcyQLY2RF4Wn2YwI5KyUb1dihihrH4MU+unv3xTwc6
DZJeBc1zkIRUKULrFJ3zqq65tLwyIPUVdYYF/Wk8ebOIGhbmAVK7MfQMIm3lJnEmpIyG0zILBWEc
ihEKG2r3g6O07sjERp6+Z2GEqznF6zx3RhroeSUL4DJM51aAvkOEN/8Z3cejpXV24yCHSI1/JU8F
fUTZ1Ildo+plOczVU8lAd4lxcmj02rliRPbtcCYUIVdwLAKBCeYzl5oN5wW169/Nb+I9woWFTR3h
yBTmfEsLXnR4MFI+Sys5V53Whbr0Q853VfCmBHxFvWSQIHDDNJ6ZL81HJowsds3fU8BBm0fr1GpO
x5nSYsYmOgtKu3aYzK1hx6eovfP6uz/z3KJWtOXLhgWJmLUgEQHGhrslUKboymMCINN0/KwtJe/5
+6QtROIznTRVyJyARDuvFfxst1GiWVrJfqoMc2BHSEDvXHHFBr+BCqklGnmzzV12afFGuXU37iiQ
ISWVpJfkuH3tWvzytVTlNeTnveL7zDuzz5JWruMDdwtRR5xlgPPFMxJAhB4R2i+fROGTTMC8evxX
bit26/ftDziGQTEJkoko4qYsPQH0V/WYcoD1oVT2iG0RpfyMhhd5tVYJt2u5j9u5u/RoBbH/Kfi5
26LrSDFGmLso0cD/k7w8hZqQvm8lDTHVPaCUGfNXVQ1yoPXZq+x7WL503Y+qTgkFG3okrXjdq93p
jkKxlJwdVAa/xd8W9/LqjTHmB+s75ffwXC5k2hd1ivSSM1juZVQK9m6+z9iXLiZjMqRb1PCKpCMA
ezwOsp0T2+Ls4OuRma/u/mloVceBHDWger6HFC9+nIFdfy/flzwLTcg8PDl5i538yOUUQynHke57
1YQMK6eGv7+2LHKmxepB1928+P/amHLQ8w0kYML86c66vMsaCWTXV0TTkEPzUwiX+hmc8RrqzPIl
3kc2Q2XWA3mXgb1jfBBrsovOK0v+RFvPetcoZ0mZVPTYv5AFQ756c+O18x5FCCeg/aB8TJln4BMY
vvG/OFfvoftnEexamKg9/6+I4C7NEUaz5gTl8eAs/aMZBqKXx0Op4NOTnaPKseFofLJFZAi51lzD
4SFHPXpPOvkpMq846pJub0gFCI0VDO9qsB2VUlgAByOvut8BT93HqS5qhPyCeBCJXRYGaD5asBJp
30PIqfxLMz5AKKvITAm6hXVgdo96ePQLMQiHfO/Fbgx3TGGdcZM7EkG/xZuPPKxMZcpIyTYhLa6r
9vbCkuB/oJpk4YxLVXAwzvLb+3+OIp36t4RzXpMXfSuH5dX7MeIUtixAq6WyA70OmO3WUI6Rd/2f
27tDzMYOZZPSRMeMlrAuQ7MJstPnc++W3O2YkaFDduK367QRFmSOwMwwEJQ5udSK3b7sTcEEd9nf
T0lYvAs3l4D+U9eORN2flkz4ZELpDQ/CY9zhHC1nf38JKFC2Z9fzCeo2XHjGdLMHl9ZXtTNG15Na
/M4ntzTqiEI8CzhSghadu6cb0R33GCW+pCHInErpjIISmJn/TCvNO5/hkSYXIoCb2BlvwL7f/Onr
KAsghOkR3AN8548I0VZfbwvGtXpt98tXJKsevnc4mmtP8LtgpnrJ2cAqqjyqzqrH63FP/SHcjFWA
h2RFdxgpZrp69Uao0q78Mlu+ob/+tqTNF9YeiSU8QJqOIlLrO/lGw/qjCI23pp2i0unFCkAfF4ej
E1Sr0CsxUuER7mrxpSJ7hV0jjTTYoiVvq4ATjV1NMm+YoftBuDkLODFJY/+p8Kz/QWRBjZ2vqKug
ul2stMx1MnZtoU/q9A981rz9jNvrVNMxM2KSojIa5Obn08m8519GUwLkgnHP59sqtaHOwtmVGGTU
n9XUB3yujlNwBYKNRwxslnBtdKYjGRSoALkGfGnBudlFu7KQa5/X174rzNrN2MrVlIUpGFgBC6ny
0i6WMYGXqE/9kQY4+SFVcZWDv4EkXjZsF+KtqL42udOjKyBtFxyI8ZUC0q5PEfXVtj1lkO1PMfym
jfLu+xYDUYEHefgzXdSmcA1Mx5fMYkRGqf2t7isnskOHqa0gjnvE+88efwkpO517vT57yPKi8HFd
YmDFi1dsfaWBDNWjVvi6X0AuNO4Yk+xOSEG/Z7Jm38XG04ePTdTaYmc99ZMIy+KXlLmPO1ATp1AI
rgK2jDI/g22ISkd852ttCZhC5y29fcO6Qi5S5UVanaEWg8Fcc0tS5eDwIAMAzDZAf/3dJHwhgSQJ
SSPMYyCps3vyGRSA2OyP0E9pyzpBQuxiFkfbP+IxBZjz2T++ZXODVz+gRzw1sHNm6uH3HQCvEPFk
sZCG73QdLFb7v8eIT8P/sJl+g1eu0yhZqLdkrq8FHQWTWQVA5o+1N6pvmL7aMnai2vJiZSAQnUZK
GFGy3HU0jiw/xUUMjaVKf4d6dBUaDNzD3OePFR/YE8CQcvy+n+Y2ImBWdxSHfJ9gjkQ1GJY+Uqba
6/OKotP8PgGvTf0Nhh+DOxy5K69a4No5jGiiCbv84tbxTzoW2FlEQY1yUGwbO6Ogl4Wx7tYTrX4B
1EtIznF5G2BQLw8SccBKyXFWe4DAvper049dg4r4Jbf9fuPvRQ+3pk02lWIX931G3AC5PVIXaBk8
2Yj9Y/+czoy/I+n6SC0TxNV9HtoLMDYmoI25pOnRWW/tdb0oMtP6D5BWIn/3y/yBzI+M98ZfZ2jU
0qBYoxeAt3wBpOZd8e6fulE6O1JyLwfLEkqR19rkH5uV5PODgOaNVd5l7rO98nvChQHUHHbnDxu5
A0OB3qKNjaGrl3qVztf3C2Tu6JOiRYR5hsYptT0BEvdCOChzAqZ4o/3recZxVbtsFrDtqCM/YTTh
MarsRycdqkXu7TVk6CaScIxgbFfqaXxIYAcT0EQd1+4wZ6Sb5nobSRa2zJGOcwBYyOJObh8759df
mMckhfkboDZqSBEFRUsblxoEsVFVq5ib976iMEn++lYWsSWm5l7yhLdYhj4JGIoAe7Jh0uIwcyZO
u3RJ25+6qUjr/59lE+9EpnWg8iXfVh3uzrc6/hmO5+24VK1w6UymEB1NKlIYjQKsh4H/KGvTHiq6
ir4VVuojp7AKdMJSohD54Bj/p2Oy9mQW3HiXXGFX6K2GcKFeFoXAq3Na8xlFNJ8x/HVWDOiygFHG
vYoKDFHDKvOGfdifiPdxPSQ2Gm1kcsEEan8XkiwJ6m99r5FY7ZhtNq8h8ZTM+4WkEkOyUBXj+oj+
M9tDBc2kaWQcWgU3JsXK9rpM1XtVrnJY7IgtA+jg9bdJ9CEtjcvRrSEe9tRjHBn09/MFJfd4Bdpp
p9Rf29CAfbcMpqxsQbQ67/xH9ppjpbXzQZFVct/KR5ZX+WNZCkmuXWCOqjueaDz2v2DvY8RwYar2
2zEf12IM79RIwvOmMGWq3NuDI5sOdIWCUzwlTc0QEwQZN39yMcyrtwLUwMygngVLgbMEBrAB9rFo
UqTR5mApBlGOlysIzc5dMJGLVhflwsMXXRvQI9YeAslruQ60ZkME/1NdwjMxUMx3dbseR/GqK0de
KAshQJ93ft0EwkmOO0MMx/fJ76MFqWfQS8N3aUT5QVMQbVU8+Ujrbr9DkBm9blbtvB6u8qvJLq+i
IxM5VjhQT6DFS1dSAp/b5L8a8qy/GErkf6rg1ZKlQTRTw0WNW5+gHLUiZKVURz4H0t2rD5M9vQxA
tDZhZrPdGmnahnwSfbanaoxWvvXWft1Odr9tCx2GKS6536jDb1jyQGWIJzNyXazPmN0kw6o98eqB
yC96iBlTqEuZi86vZwp8eave3bCsMHv2177ghkrXx8MqwNPtjokgPu42uzHXrIfvFABZMa2eQi+g
PDRrcHbxmdsZmiHeHfW6OrBuv/rryVZUyUNPVnUEPZiiC1hcVXKjBYyIabsMIzfhyKtPWq75ED6A
yjEfVMTCqCgK/1B+b5nuFCeU4/oD0Ee6PDdpIrfCGSsHTWnh8jB81FIHPGN7T0TB4Az1Q8VSlUPc
09BcceIAooXD1nqvkWpm+xoJ36GBrrikwlSshkMgm6ixDrT/2Vik96wztb2oWk21ZywsMB002sXg
GQ2Qq1mujQzvTV9Eg1m8nfH+Vl8vIKfUcCyjXhJcTGfqCRmNlH9TADRn6h7ankLMEaezPpvs32k8
JLToOhe6BLVraXgO8J/4aD7bJ9dPTuxtasRhcybwCvN3aNrOTID5yV+N9Fwz527y5IWRxY6/xS6u
AzEfqiPm/vbAP063YFT2kwQl7gC8o5ma+6RZMkb2SEm516CSTQxbQP/Y7Y9m6oqo72UAPwImUlbu
MImwxX+iBCRb1LXnyj/5v2mnUFsccp/Uw+PcDaTf0pPftMa2MQibYO0lO1RDD9IO/TWiVN8l3uob
ubJdjyBjljxqLNxF/DHzY3xEGIx3ZQss54zfPZrZz5nmzXuyNjxwaX/b6ZFAoAAcSHqNjQH6pFFo
q5bOLxDM0HiymO7LmkBbk2yoVeYRz2TmKdZ8ohpWjD0PxM7xYbEW7XFUYDCPCA90rsxAKjAEl+sj
NU2uR63EKmfVege1QMUHluGGPnkGgaTAhKA4+WjngfJsDEyi+t4P+PiCBQKsvlx1X3Ucy+Bb+Bod
mpagAJIDUB62jMH7SrpjB48jnad73aXPLOS61WMtX5eFfn9JvfuTtNVLZEOOU8/Hd0P9PGWC8Kbf
HqiEtsORdKAE1CjrRlrxplrcfMwHnwRX8IVhdMYzS8wd74YJUSp1qMMJN+kAM6VBk0ROCbg5Y5Kh
NDn/5wRVZSNltuEAudMVgqIyVmK2hQy5RxaMmmxv/jdvbiCiaZrU7QfEUA0q5nQBgSFQqFu4eVp4
Q1OFayl7OS3oOAF4BUZJnmltsSo4PAj+h8/4vebZ3hbxmrujEw9DS3XZ8AmPZ+s23BXVZ0oXaW3h
k3nfSOnsyXVJmzqtqf3VaHVQZqeI013y31YGo43grUvqPQd5W33wFFiHbYzd93wP8fO0ZrxlIYPr
r4bZuWk+cWvY+DTVIjzLUPBCuQhvUeUtiK4+xXlmcxT7jPXCwzQSOuxq2XiCRpya9uKSE0VRHcTl
diO75xxSAso3uo3K8nIYk+lYkG6HeyrcwTHpOSrNI4iyahKx59XVIznAwFFyHM5/KRMOB0on1Ziw
PVm8tdl0UbVxH7g7zM03GKy7zYhaWGRCtoIwgwvP79+aViqoUJ5rnAODgUiIAlxS2LtoEe3rKEPK
/njOASCc/y1HX4cmnJgZVUEmvKID1gv9trsd9KIkP/XmO/974y34+XHjhs445T56zvY/Flktx/3u
dz9gsUxVhjh0p+MiAOvN5w52U7R09QkYiuiidlZUNOvVkIaAmYZmeXavyax1BUhF3JOGpwB1v+0f
Uh9tdnyR4Wl3VHj48SIZORB/xwZ+FX6/Qz+V0b1Zx68A2ej1NGFJZxqH6eIW4QmqY8zpqwclogFS
O0u8fLV5AiXLJ7BzUfQjuTMGarYDO9cNj336gpLdlkzrmGx9HCc1E7IxMTOO3Kx7pFUWil22Mj3M
0RcURxHX3kyohDLx6vNoGfN/XLAXKPRJpKpIAL9fD120AVcghav3/cXprst6BNH6Hjvtpc97FwnW
FrC3Keo1RJgkylUZfvc5lSqcSs+a2S3eH03QU5RqhGfComHkEoXLdyGWK8N1toeJVnEMze7oNGIQ
u6fEyM2StskX6tosN8n3RMXC6oNjyMSY/M49ik2Onyqz6XDYgTcmNd4pAY76WVCqH7ozODUgYV46
Ob9eyI9KJPOtYn71QlJ+3V9Bk0B8Kc3TAtED3Zom6O0xA0vb06fJCqLhOfxo7YcGWCCFe/q4N1JQ
0K19V4VY1vnIfg5gYbe5Aeqidt7GANx2G6drwrkBhRRPPHvBCT7RiSC1Xn7/ZLPN9bTUzdkNn0TW
1+Z5ZUNUDb562X97UjKbHkPuc2I+j/wGZDFcOVqnEoS2BQhOT9wCMOknp9ElKcVctWFFclBthmKa
UCiNmmtoL3fMaEHA272s3aH6mNkfUeYOZ1sTKiC4b/W0Ej3Ow4aYPO1fOZBKFpz4ZSvt3ROpmGIX
ZuCEcOzPsvIPtNwUyz+HXRdZKVyLAZt2gtfqmQsJJIWVKKS/relYCkxHAzvFxCwssksL1FFCSis0
y29jk8faZ/cpLtoAISPl2l8LdXT+GzF1M1LphPvswdjlKoExrfN1wzdyE9jPFhnFTXeAwcikQT6c
OZse0/006PVnUgdFlUjJ68gkYaGSVU2uXVBqAZv8i21uATKjxZrx6m5k66yg2ilsv79iSuB3pJM8
SkHolXSNkSJZKs/wLL58CnAfsh2AMkFUsUkF0n+JUCR8d2jNkzg9Oztfae/OU8lLQcnQ4yGI9SMM
GssroDyLGJ27d2cu+vkOfaIAIRmy81oej2MtlCOYqdGXQkYDbCseRwcBoC0n1bbduYamScr6yVAs
V2xQH0y5OnZAGQFx2E68zB2WucM7cwYruJpay6WNO8ruz/K6pxTbQcPTScD424MEkLOLL56Y1uiQ
qOQDwZrs1QcWKqOHXBDIMS7SrQLxIyUuV6qR/ljIakurEtLCGhQWVEsjxF+XHdSqGQHbUEWeQALq
9pazyviZmrSuIFiP+jC4stfbqbtboJiYmefoFfK+l2szfXVbtrBH7mevtmrADDKoXGZuccAaDTz3
8XTiZkAUDNxpFOQYPAAZBz/vVXcbuB9aTV6Gd1J2dRLrHj2IeFXiVHMp4OgphvNOhHXSOieXFlln
u+HswEZ9Y8w+bQFuC5YV4TrePX1EFz0kWNPH0EAxKuFykebyBOXLK7Rrotf+N+dHNniSrFst8isu
ZLdbTFmXSJyvZM/9CWjZYVNITZxQgLPB3rJ65yM6Uw2tn6XI3qB2cOqeT+IvfLPQqXN3U2t58PIN
WRLN6SJZHy0S38EXL4wuON9h4HAUrUUHL3L4E2EPzysTFUwj6lsMW0Fi7na1qwkbYRZfW3oWI7sa
CxR5JGB4QOQoWVzNtRvap3ntpanHmrcaN90+CubX3JzC5xm2flKQepVKginH4EQ+Pk6nZtAKuxxK
d5qyZRlasffiGdZ8d6oRrMA85KMEq05SiQadOM4wsaN+dheQvtwvek3TfnY/PDYN92E2TUzS+RKC
JofZjPFvypD74cx/4vD+56hgpWGuq8T63krP17VMkP+m3Vo3nGhayBlel1GzT4p96CjoLv7de7MI
ZkDHtSTMTTtTlOalkKMQnkJFXOO9ZM4/CAgMv+MHXiGlrE2qHR/Xxgzm+ED62ckldzFa4870svV5
vhaReyIVYN7tTUkDF22SfuiWTxErT97EyCtUkt38fj6jo6xKcpSZjjiOHmTkeg6NvcM8ojNURmLr
gsnIeB1Ffd+RMeqiW33ddGtLRIcgcO1Q545LEgX4BOqd6BAsH/yyQ8liLCP1zVpWq3ezT//HA8dg
9+l1sBtViSkRCXLaFmONGcHCTR2KOjkm2Z5LNY2cetphD+JYIEy5FlynYuBj8w1l996EXj0w8OW8
QBwBgyVzWFdMB4G8TzCcUXznxVjQk/L7OrsVCMR0HObyjt3bwg1ZQgMSeW3YT2RKuURdpkiM8JVA
Qjo3o+XUik0j+6T6QkwYEZ1iHvdDh2TD/h/MpeOa0bC0jVGks8dLpuOxoI9ospwpD4lZHEpifOHW
iBjdPLfqzaRZVyJafl5XofDt2oBJu4241MLPKbD40lgNkcS2uWVdy60ImtstXc1OaFrZuZWUpIYi
E23N4uoiza0gj86xjfmrkPTmCwDTmNCM98jvbiDrrdzbWy6k2Z2b9UIW6vANaOUyUjjDCh3Jg9QM
jGeEQ+j4A0Nc+lbtTROqqNg2DUNHp+NmoPomUmunkHYlrlKOU9S05QQGpeS8gBtQ/QHJliTKZA0D
cev8uHlDT03qPjo2K+zUmW0UXffkOHB4/Zukr3Ra7dmQgjyff9tGEx4mmsPsCAzaGU0faV59mBfy
TPt7YyvlgwLIFnUefnskGME49qp0F483ESDbYtbgc+ykhH2QrIV4ShQxetoMKXsNGa6AHeqUI7Wm
/7nkFzNbIDocUCX9/YZI7eP9Ynxyk3U9G6AxQYSUPBgMTQM1kR3XyaMNIAM45gM/i8aSKzT2YsM3
b6oTEf2Q9GiejCHyg6POCtkGF+zVpPoW9d0Tcx7GfUhT5rqumYbpWzXNIrz06P2G7U89FcYhZ2ow
2Z6l2LEJQOdHbMGl2mtKDXundGQBNaKgphvSicqURfYwvR1ciyOyOgnzO4Oc7HyWAtcCHpEl/arQ
ADDmczh8nnW/BXQEI7CybfeD1SSorVImFCFP37Dcg+rwZqKtjMReFOGCeAYq38/KHKD+YsfR6cK+
BgN4KN3cX4DFWt3Gquz48SprNcFkQKNBRVcIRkTR9ZBtvz6m41qp2XaVKchNC2E5HLh6DxLysRgE
AaEAkdtviAfPXuoMZN+zoW7VWOeMSbDTfLGKqHpDF078vRdam1bdWJ/t81dT1CXeG6nAmTWezhvf
EX1peIPITXBj0W7lrCeInqL8Rb2q7Muq9mDZx8Y2kIR2F/75ZPGm1RflmRTGpTQ8hYLEKMTItrZe
P/pIjs+/Xs0IfLGtteXSGFVFJxu8j0XzdJq6vtpm2bV9+2cDwVxNfVmq07+/jFWguoLBdJK81jKp
TtAeogwITljenwEayyXszmLXdnT3OuanzqCzfRNnseNZBHbcHFYSyKWxKvudEryZiz+t/ZXHN9v1
TzmiBRZdUYRI8C6hT0ebNsG+xkijm5dPhHK0KFHlVWsOYXTU3cry17y7afA4yHpI2vYzkX8V/mwz
5+03MfCtMlW864XOmKaKSooGJIu2jXZQvd4VfOxRSAaq8ar17Gjn6MHeLmbGH3uoStpsW/aZHUot
nIJoOf7v/9PT5gD2SKUFSAXGKkBx8MhKRS7SS76d00VsJWNVYtUubty5h+sxxfYBDnvL+j3cqQDn
C6iYtYLT5DzPwr0QhKzgkxl32HAZY2F2FIOUGEMxVlXXkHpPDs565nGPrHkOXzMs/iyPEQpc1Mdx
UjAU08QqLrjZbTJvqMfrNOZFSJF6DjcIGy04lZI6vvA/ohgkoVK02S4ss6zO+gVe/SQ4t7r8WKHt
FVzqxm7gfgAxWkaWXK+ovx+UkBkvvVvNxLk8AmNoHsqd87ZNmPDgccv02C6l3Ag3aPhsAnOElxn/
GfTwECdZ5qqcrSX0+CdnmMzxjdProX6iSZMFNxP+DdqA4lXbqZ0LV6TMCYuYSyHI/0eGW+Gbpbhh
o7dXgS2e0LqMukJCIGuvWn0F+jj8Kp+5QAzFT/HhEpLgq10I3ToIoTIRGfoiva/akBwM4cLRb035
bj+S8iwTC9/nbvmYYeAzUwrYMpKl9FYeL5dLYa560zANkQ2hwaDyTfLIaGDx+6mMIfMiuR3X5f8I
KypjqVqfSS5edS2EN+G3ay7cdIfV4wHEYDE+ga8mEVMLeAAr8j0HQd93iy+MmfjTZ/2nRWpOj+m6
RvtPr3knfXckZy0q1+w7hXVFHjO7vuLYaKg1OVvXyaZif9VYefe7JgMGZf9hSZ8EC/DJtih6fuA4
ukzRMLbYT7bMpNum13OoB0Hax1V9AxFC+HrJWMPkBdGrV6RNXSfx6Ni02dbiLiXhHv+FA0aFHFm7
KjcWkKWkw3cFXmmMSoMJQY62G6wetQKGMbsLvosQbdJm/l2T6Y3Re6aKLRHazrR4iMHheA1xWhGN
wW+cyttbO9iBWWBfpuPcFeM8eMk4ReMljvCz1KMI7wFAeVog//Vd7E6B/UjoN/Mwuj/PiksnwC6J
FVIxBEg/7MLd9KdpCQuh6T0O776M3kx+jFh0Txji0jnfderBXi6hneQ4s1/wst4UJYmTtQlPm+O2
QUE38pNcvNMCPc4d7g0FlmooWFzNQoccA7753kms4fLu2HzEzV0zJ2dXDTN16pXFUETbOm+W4jqJ
7sFO9dgTEtvdhRk2rlpm0BUP5W7qizIQMuC07LJmBQ8f/4BTMISaknBdI1qwwsqcnya2iygHA000
+/e6DHgXX7ANkqg8bx6p8hB89cV/NjwnhTIHF6rl8YPTdjuADLqQemRgHLbBzEuHCInM9Z6CDLMb
SlzO2gsLyTv5ZbZS2YAkm3cPQc3eDyOrbDNRoW70H2xhCBydv+ILDREKgn7MQuVl/ILZr31gYWfQ
QUfXZIXFNh0bnCN6RInRW2OEmdpLnlljXTL2lnXv8ZUjF0VqhEHNIjJDIFXpP9A5/cHyixCBj1M/
27GrJXoUueWgyH5aDyALZnv3fGXz8VnmYqsJwwPmHZgLb9ngHETREB8yRt+DDecaXxs2WyZMB8N8
L9POUuxu9XdxIZQL/IXSZqE24aYudE/zuhsh63PKBq66dfB1Jyleyt6jWrXKLngS0RuV2csxFUK/
Ta/PHDaQ1231Qjqw43VxxMZIu5DtqhwWI/VvsxGDFQaQTw2HbuRdbXtNFfaVhTRJPMIjTUgUxZiD
ZM/9RHC/Td4CAoMA6+dO7TLWW3kSJ4ZjFnrp4r+Z56u0b6ZSbejEtu+aWpBiR9P9aZJIV6po2+uW
r7pFDgSFkJfG0vWfCDsmLgLiqf7K5tgopOE09ji/opm4DS5N4OPAB9WJeo0+KmLexE0ris511D7p
kjmQxg5pe5n3tYtudoEOXHVKu8WnSHSmlLTdrVLVKkPzpKW95dvmlI33IXFDrOGBwa6VWQOoV9vO
9HcLyPF3QHMLWOXOTD3raXLTATtf/6OZqzsXjs+JyeDRarCPinHjdDYCqBrPslZxkkgTEAtPIYYP
2aHvCmgncvZL6YUdMQZTZKojA1ze8Bqsj4CBUTuHbDs7Aq7WXgigFf1BQWxbE+DXfF5DiMJcDNeG
G9EG2Cm88sLHShjEzH1nsCODNunEr7XYN49CGUuvzvAY/1wRyJQTjYlKECEpbJc+IbP63r5yduRj
gfGJBk5H2716CJ9D1NH9suoW9/06FLmnmsgOSCazfW5MQ6RhWNhObCcKAxA7SkfsBKlBy7C9hcG9
St7UW/IxhHlQi8MZStFyIaW05Asnf5JHCitlK7oqT8jSArEw1wJ+8JUD6We8lhm4wsf/GRlOxsLV
6WEdRuBdFc0i3BvjQcn6zaTRr3F3sidHDFJmaSZSefbYhXpFO7xt2R2b7bqfIrWhLhV6jEfNOXnF
8eVFDViViqvX7FJmLBxcLXtUjzoEif5lJGtzEA6w4ujJXPLlalyHptZHkKtOaT/H1im+S2hIawgj
MG/ZLQ/wL4FfN1ZJFVsFUd4qAHNtnnAevZjiGBQosVKKa/RdjV/whCGEUH0tn0yI8QG25bfrlWeu
L1x0VxBCRKnEvrrBd3o27iXeRiDMHS4xyK+V4lRPzJq3Q4Ze5yKuXmFsZ9WNo0V0icK98e0xUeFG
ytXj5uEFFkRIum/lzKAc3NxBJF1/BzLmduxbNUIp3ZBTy3Kh6BgQNG/sLBmDCMhtOJpdXYNl9g6u
TG033xqa+vqdxfQYGLTiqNNbAlWpHxvS7wpBa0jxs92FS1C7fpzQbnr6WQX8cIzkT2DvOw8Msl7h
NJO6idejl7mTGcwIOFGYZ8lnhrhFwLCLN5LA199DdyvRGLbsgXRkTe1XmflIYuh1pRc6mOjJSdJR
XM69aUHNBgcju60UNHbTkA3w4/fewuC/rVaFFPwq+Y8OvK+asONE5YW13Sct1loFpozIvU/HxeK5
RzgZH24v/xGxftbByJUIzS3ln4zbl4R+Jp/3f4rzTE6wVBxE8Qq8hMw+hCr4+OPDk5zFoHdrN31m
TJrqDOgy5yCGlrn9JvwhFwpGat1IOMsQtpFyEc/OrHAYVo7fO5+depqyfZUX5NjYgec6HVOGuIuj
YciAG8Uv3S9Hg2hLHokvNX4oN4EgyAFb3JD2V17NSNvaKw5lV6UOPMHz19FrJ50TPBwXZ3tLk/Aq
zPAKVxd8b5fJ6VkrAS66uEdhRKay9poReBF2dY2PAv1tycjSM76eT56OFoz/oBSgwqFDEMo4r55j
nfzqMXV6/trh5cm6NrVf1rfLA9tibAyI66SPxAu14p6CHurxMJzMgaetZ2bchijXe34u/lF/AtmA
e23zAg/vG4hRCZyhb998ZiLRWXR6XyW/jVvN7zwlvMcv9fGY1EQJyJ+61r161/ioIAb5UvBDd/gX
49wSDqIUxHPaH+d/5gbNbXPhswfVwxVfq8/r9j39s4Nkl4QZWbYM6sS5yGthxltriqz8r7f2Do80
TJdvJ8/FsHNrT1kqexgHdl+NsPTVWJlNuthAVv8Zr64NeCjT0IOKf6TqgPDbLv58MCYYj3XIfcwQ
7wxtbeVmn6UFfnc4OiD5r9glrWFIUJJn+24bjv35aLUAs/UcKqDxQJ8J1UGlwronGOyEcsG/hEdM
uV96EVcAOpvWcVG9vbkq9XmF0KBsdFHHvCusAVpFHvEUoakN4wV/d+yy+qPqRsE/zyPC35vadNTS
wGObAousPq8YtGq+oDiYOuiarcRm0FvkddPmGe7BwPtaKpTpQcNecKCkVVtak7+g22rzq3LJ0mnu
5GSku5dNroi6orkv8a3xa6GJ1N1enPhBZhvgJt4WpvVgB63VsRtCIO1p7M5qywweFzHEIPVD/gva
Fv6YorxzMjveCXpVFFngHNu03Nl6lFsGSYp1HlMzR9qkFS8KSqPMhMQczESgi2+ufiboq/SSx0I0
Mt0dHFRieNaqdYZwtxdMoG+qoeGpZWdjYYzIFI32EkaqzfeRme0qAGXhpZunYvQpRAJq/WQP2PfK
AxYrFj6uoRtAiHnGGKl84IoPa5nbJ+wcuoPGFnDGF4Wq1MTHw7UVYCfcu4xrJPKH3+pstbw9URlh
FPmBDTdD9sJ+espO7ggAjuJCqP1sr8kmRN4rrlSCYsQV+dLgY0KusokdGNYPj19MjijRSObMm/pN
H1MJ0UAF8qH4ldO0G9u9HxCVt2gdBMltq/p0tDLmoWKoVcjtAPGiDWdl/e3P2txohRbfS6Mj1c5y
l5ZPT3m3K9JnXtctOeDDdpf1S+Pz857SNOFovqyjT3fe7QduL0E6wweTFlQR+/PWR66OfgxsH8K2
vkxY7zsaDCDK4U3PPBIWspAEFOEhrcv9wgukXHKOkwq92kxSLHD/VsE3M8eCqkHQnbEqLnH8xZEM
kmPpdTdnusphSJDqubMzckVRKjZAIBf42bTkS12aTUSBribUMcvg4AAo9juto32ONGhRwh84eEdr
KOJrjEAgVbC9/B/w8aKBe/zg2u/B5Rdo1cL10KiEJbEvIRX3YZnCiibCW2Bp+le/F3hIWU22Fuvm
WJu9VZcBexn1fvCJq8QDPLLakZu8m0fTU858jnFOLhxAHwZPkJ4g/H/bfxgmh4jZus9JjZPDYhM4
NedFtjQc8G6CG3BFon3idPZ+oXqkyJ4mwDj14tD5my7bMwP2JazxqITWrV4za8M8T45BeM5DNGIx
uV/zw4ddPb6VB6m4TpUWixiypsNz38hV8RsbvkytVp+76WG1L5aj+bEsfGB+WtOW8+Onnn2JTi3G
Jan/S14w9KbV2TK8DEo05x2mBGUhvC/C+tmfboZPgUpaX2R++yw1N8/jauxUj8Qg/Xb02T3HtL0l
wJQEbZ3DAoMdrQmnTsRI16w5wjsHrAMzkgLXKZPehCfrE/C5yVKv8cZb8Cr4ak8KNEWEudKYOoLT
Sz0PKN6asZhKANMF8gGCfeF/JQ1+4dpFGaxj/HiGaI10WQ3XeTh/cSSkzMDD/8ZmV4+rVUrQHmce
3ecuRBCUQixI5HLelzOezxj2mIxqeDF9rbZ+Enx7dzWDWqp3lIjlwEzD0dKDKyREJLlSCwJZ0TEt
IXa1Tu52Icl0etY6/eK6vy4LFzM65WOuv/K4xeO3cL1adEA1jsubJyARAycdG96t3QeOvg5RzYxW
PYVGj3Js9DsRMvHpPFdBzJ3KM1+sA2ompWZsi593+IXth+amVFK7qVegQx/1DtrfLghpQPMy616X
kC8yXKXRs5p3CjwlnuNEJPYTQLLWOWPGMx0aavUB1cb13siRqZVpX/krGcRkTF8xkjhDVF7n0x0/
fW4Y8LZAYxm2+HEqR4beRw+4xcrcoHWM/VE0JEsm9I+d/lcJPb/oP1U3TH3fw24DoC4p+ZJmHXox
Wbx7A/m1WSdBSYRBEHOdg+xnEG46Pdd20e71pAscFd/famJfd6YUNZd8XPUUYYxrg5jq1PhfNeQD
FF+E9bLMUrVo4ffrjKu/s6w9Uz257k0N9OVxc88SRpL1NWOQtX3AZZsiRu330KNlo8e96MGUfXWW
WHkZZAee4JP1IgwAQqoqBKCO5UiLBQmGtISAb/HcTpwOq2xJ5Uvel+J1gJYC04gZWdIQwz3zFe7m
3b0r3h5c+Nd1eh+7YrpG36hniZipUh59NwAmOSQvGJ+rneYyrvAmaww2DIXoJ2mMfNujIZx8FSl6
fRbJ7hyinuJdpGD0kYPCojM0lbWNYjBP1Ntdk0an3+eMcMCp6WvAudKsEWo+xsv1J1HeK7NaNs4s
Qi1wiEme9yyKLfAfctE0GNqP1nZMbPYpC84Rvm9xbh6aZRW9d1Eiq20U69xrGuR+/J0op7MsXnBL
BGBxaSDuYhC5nP9B7ExP5N0OecH/uAbgqJW5cQ9pIE59MMFBh1NysiiWYJSXlqShh7kla35Wvi5C
zSjgQWxOjxv07PXbv04BLh7RoK/T1U0OI6X8Mz7xjiUTyVtnam8YopUMhzboKMY6JwFkTyOxmjhi
Kj3390TamS0gPpzK0U1+FGUWNB4uv1s+Pbcd35ddVo06OamoLk3QrS3Gf/K9XQqhEWI8OWaBet0x
xsPLMAC7F5tYz3ouIXDheuGsN++XCzV9PAkK/aTvEX4iirNGk6pexdWFYwnR4i4DaCs0oIvVG+Sx
q07or3Y8q8Tz44F4J9WmrZvs8jFCV+8BIQ8wb/dz/+8X+w8DLgmdViph3ySUtLe9mu1KTovAvpda
yYep06BAUmS0FRetxK0LvxWjpYsqUlg0vpRm3D0K3H2fruNT8KtxzN8Z3LYAGcsuwytEZksRYm8u
74cQOZzLxCAC3Ne+B9uvSFTZTqNxkw6LvLyaZ2wSXOd9u28FNLhdQXfM9hSPm8OIGPgJVTUYJIsd
RxiO3hX5A37kHfs9tkASb63LdZ5uLAPfaF3V5kzHz3NDp63Xm3fbYad37Qd0qJ2hkAl/AQKPkvlK
PBSEgx6o9OyfBk9HH32ry4Hue+PTQEu79r92fmm+2zZxMHqQb3NeTvxdKTxZkrvKCuv6YGPYe/pv
WdnQp+UQVuuZybwSnWyL+U1K0EXr+hreGgHEQYg92ES3HbmKnX+Io4MYpdDoaFS/ucky0At8AX2s
qPk5tD7jKSWh1IrTcaUxe2y+dMZdTlx1Wiq6yqhRawcbaOrtVx+or2JJ1LBvaqIwpTd8ORzONM8V
NfjKbyR7NLK2krFRWmn8+yTB1ZQJ/3x1pH/GedJ7Pfo4QZZoszyAxuizBVHSo1Ou8luHLcs5RuCp
yGdgoAAjHrDwkqKYsVa+xzafeq8rYpozsehZOAhjaMpGBRvns1EW37Cz0m/0bu/Bexm7RgQg2fnu
wB/Rv/Xw+q5eQqLleWYZj/sKCfsghDWZhEXx0N32OS0ZESvX1aWrssLzQxzQjp6jfpyokccuNjXm
dL9qJAYSxCyD3ef0wL6YejNYbp7zSAlKbxxg6eyBqmHAgTqAywNq+LwfzMgegeswEQucdpnL8G0D
zbWXJ/8X+Roti2zVw6HGZW2eMfABT335s9aOh6AIJ8KK5uaNMHEe1uS9USdZuLk2rorY8eUz0PSM
UgTUovAbiRLzcoiSw3v6icOOE/ys6vdBl+HmhorWDGH1Vfvqqmvij3mqBblSX7R5J1pFablBqCMs
eUaUnPVKFqWsph3FFbg6W2T8/Y8njUulpco6+ALT0hP9tYnoi685DTomN6cLvvoXgJnBtVgaE9Mq
031YooR8s7rUE2mDuJLRS6L5lJbRa4SQbAOMNvQe/LvpgEAFPIkKZ5bl92PsXZH73+IbMLemJGbS
Euq2oicX+R/KlEEAkZ4b3ViAB5Wr8+O6uBe5STe+1IHK0cRwGyyV2rl6dVFvZqTWznT2shCkrxbm
tBihZFUOzVjYitYsshw8gULilfgL80Omml9iWPMMnhFk6Rje+r4cxIDfOElQ7e7f6f6ew4RNlsbA
o4hhGc8TnX/FnsPteqm8Xkj7kig34TPk/FCXFa2dM98jTcTgg4s0g7YqA5TfMjJNxlluUG5SGQRP
fwkeqbKiQlC9q0JBHx5vxljrqRbUKbNmwb3J6fptg5XSAVIE/MC+an4pLOx+IYsrs4RKA7CwajTS
k8PyIR7HbT1cm1p5BF3Y3yh/E2iRg/dQKaFWQtCXn1fy6PFJJ3it1vrr+e4yEE0axJRrf1FsHPD8
i+wHYCUlcEtpu2Xjyi54e3XmRiiEkge0hgb/ZFK6csACim5kF35zrsqt4CZ1xJ9DCSps0u3J6k/1
6iwlSxYfqKsZ+4vU5F4oU3LgDJ0iHg82rJqXsUGhjULFrHiI3Tl5XXUBu9PSmHPr96Ey7H1WsBgC
UjlmBHNovbDBJ5jrZwF6R5ZI7d+3vb3PfinXkLtlsPbkMWeYQH55k97fYz+PrHAYBIBBo4MWSNwN
PB1p7qpTVywAQn4LfrhTfoDQXnBKu57LPT0LejRqyAL/0pIOPHSFqgBVguS12gEgny9jxsf3Qcy2
T+R2zq8zjhNvDZdLChXwukfY3ml5IC+ib0Zje5Qudpg27InQxkaoSyyQKvwNPO1ZSOBCaowYMOdL
V8ScLhubJ2Zwst6rRbA7iTwNAVYNibyPacWEHvkrDzik4t3RUNhXU7jrZWHS9caJwxf7KE0shfw7
bkX5CPGQQvBwehOY3HjgyM5DsOr5Et0bdHJOhf6nEn5257hv1uoZZEbtgd5frTCdhKxBWdAmHwyV
C2L7DwhzX+FGcGEcVl539/RIEr1yAksmEkwIjLL8lRaKL+xqd77iAhBIfzkUZxZsxY/POAKwexlV
MzBrEOmpqFkD4CA++BjAWvBmSYNjPNkJNWKhDuMv14uOzsJp6sjeJQbf1LbIcKJqV2DP/VZpGYoT
bOYg7Dxo/bMrAUcnnJe2pz9sHxwJUvfl4U7K8dqqT/Ic5WOqY6qHsw5ZF8JyJKjcJnQIvWqbJCbW
v7eb631m9gKAtzaQyIC1wupzNgUL/HV3Q/UIT77Q/1BWNSbLXjVbPSJ3tG2AOG6hzkMYko773m9X
Es8xPDGR2uYvTPnMlfVtNb4JREqb/ZTet5kyLzk6M/QJ044tlnzmG6qmmgYaw7PGNkfSsH6FCkZ9
TAubZqZUl38eMkFHH5T1/9fYm9Z37Pc89s1PU5S0fNoOnKM370DFr4H31ZGo/tzh2Ae/dxHxQFSK
S//qk1sDsm6Q38EMJqjCqpI4Ksdua1xChVkzBABqPIDHQYm0iMyhJVVtSnlYtjd23U5/UZZdpYWq
erZ4/D6I+NVt37mpj1eZ0gMnF6/2FVM9EJQEIqK5wb2jO474JXTii1Aqsb2i6Q3Z7bG012kVn65h
SpF4j95ezue0GQKaaBbOSjiY/z1ScJ09qevUGYQtHwoqMxPJH6XZihBB6127y4RljQ4CGmpJzpGn
321w0Bx5CzOI/cMKPRwgPE7wHA/dOZHdHAhKlj0MUYJua4SC7PwW1z23G27BVRxxYbRnO4z+QdkX
S1ubjzNsTxR2C6I/m+1/7yVf10GtAiU6KPE5j33BvNr4dC+YFJXWo03lmAZGkKAzdF9eBBFvGN2u
+gn1PnmJC0Rnn7O9EWKpwowynpPfiBuya0BJgONuxbqBe9Jt5GlvvN4Wi8HpF9JKgAlZgtExucgi
F3NHIADsXw8H1vDtD7OI+blemG4n5hDYFGW8H/k/JOaUZX8Co2OrN00Q8MEfhDGk8ymCkrqseIrX
Pi5KakQ6zu0e3P7dYBtYziaDteCPpMwj/o+RSRlSbaiP2fftSH5AkqWkl26czNlQkyhVPyFqtxlJ
5s9BG6LV2Qoo9Tli9SH+Hx5tpa8Zlk7Cp6M1IJYOfXKM6qhn2MldkCwa/fw+m9S/e+xq+IXnQYFx
oFEIQEmJckRKjhKRLZP+QqDTpVn2on537GkGtytS5afpq1KUz3v+knsZgXJpKvBvA8rYB+7nKLvT
KPv2DXSo9fC46gqzqy8B8XY4IvGPgFmBxVKX6YkhVTR6R7Y5bY/qLNE+GbH5KEgiib50yYDmgEYJ
kMLhWKs2266bxKSwwUdsrgKlNImGoknbSNnnCOzsRNK8br1YYtfnaa4Y/V0mLJUC5wNb1SAYqRZz
4iG39PKwhBjyq3U65ZHPnVxu0htr0GDRnOSSj0vZH6lV0jAzWvGeVgYR8sgDIBAYnHfn52j6uGfX
aGCR63Ne5gkA9devNK6Ir1sbbZ/CjvThAzc5TegvSjnL3fX42CxOMuLHvmiyfiHkcUUf2Z+tm3aU
wcHUmXT56TmCJXYe8x9SEs0NQevdVtMIa8UWPRZ/NZkvt3qPM7yF88w3yZWEpPlk9gdJtPlXw44j
ILFbYzR9QGJgfoXAYkKw+Ze91DVdv3A9/LY9rTNQ2iRjLV6VguUd2pqzArci3iNJSAOxnEOaslzq
fIsdWwQKqYrrE1UrvSoZF8ewz2hthvpbzhGzN73Sftq3O+uN7PZLJEORGEPYjykaNWJASjoK2GGT
i42UOvAbqxiwVJUI8IxDMYw8XKmCd3g3cL1aRcX5CwWgYtGbnsZenjXKh+GwWZSoDP/Y46A/iwPP
iUE5Bxb+VKhpxrmix1f1hxAay3JDw+GLEj9d2o+Vhrax86YidflKcxzDcxbX13PTMam0x3wyaj70
AhDk2dN2a3ok1ntVP24krqkege+bakYNRNsH3IKuBg7MO9w3KZQcmtAW7JWEVlegfntW1bY2vDq/
+N32YWa6YSFLXe+9WhO8GwKMDe2ViiA65oTkZOdZD08n96hG8gVC1HBQS8/4v9IFCvWSkge62GCW
p+Up/zHLMk3wNaQeRb5hfSUmK6az3uiSQlPmLFydvY/5QYtndmJ3QA0LqqZbBsSQyMtPk3H7QzkX
nD9aGJnJqp7bHlyhSN78HbjKUqT9EX1GcWVB5CnVEj6M4TZV+2QDlCVEA8Vz9oExLU3dE6kRjenq
DGwpsBL6+b2lAh4HXH5Z8y7q8MznFOAL+ZMJtdaWfx4dJYrNnTuGUnhQeoyyQnUSvdXEiZgUTi+x
MYPIY0iR5XXs30BbhHHsdxzT02+gL77942ck4cLTvlJyWuXXMGQORJMe17LtmX0veCAvofy/xQfq
B6rsAd07aMfbp3A1DJM1O1LG0d7C4ChgJfWyMjxHBeMpkTpqEwZoWVFBj9D5XSG8oTVZCG/Qjx7q
r6eFlq1Mk6v+VdAId6b7Xndo7JUJED8Yic2V3mcKZ4BdWYU3MkJYY5KP6U0uO65uG3qMBxGGqeG3
AsP9GD6oXZyDTczmmxbSrAE1+1irfkOhsZduQM8j5LWr731VjxrUG5z/ca0zJ1+O52q8V86FJ1Jz
wLfn1dX/MknXNnutDtbsXj4o5I2wXrmfFtuMLOGWCaKmOvev539XyksnmXvFXTlw/dRirR9Ps3wm
rvu7DJEabdlwYqbMmPaFd0LnzcdLysctUH4VSecMx4GuwFUyARfseVxicr/yh0NqT9Ysn1KXObxE
VUiUb0q8IyaqnKjjw97fxDYN9rEjGPnQ8mZ4bM07jXVVA98lagwN9lIAXlDtHcVci34OcKRvfW+8
4RQ4FsnhphIbMFkit/TKclaBFYY8Eou/38zmlcUqSqUqWFZ04BZQHo4qNrCAlQxdbE/t7p/SGkmI
A5WHD1umMKlo2paMFfK9zHGR1d71OxgDArMLLoIv8MEkJr0auQYFyOZFIfOia8g3kUIaN0j1775F
Vc1RCQop/73D8OV6LjEZQ6qJXF62quJBP7FDUeGixJHxPEcm1kPOEYRaq1pbKIwb7nRCTWqybc/4
LnQnlAP0G09y2t2DPnu4E4BgVscRPeP4yt1Dc8wFQnIO8PDD6b9BH9f8EKhcAvaWeeePF5ao2vBJ
xX9ERrE+YVJvI7oBxRvOtJb1xaqVlQmIaFE7s63plwfDVnC9MkkvcdLvC1ban0B6gNQbVaJG/G8E
entvarN06fkFJXn03a02xih/sad9WMjn6jGWnCMnqv04YoTKnQEja77whjcSbsrAVlz8zXAU690+
Ezu4uH2Ku3mGPcqpHIwfy4lcaYu5c9bvK3b+ZpjfoUuNOvIr+OYJbT1H/p2z/DQN6eq+qRwGUFzk
ZKczUq8XEIi8c6CC1RlQrCOVB+o5NzDtcSlZWdzZ4eDSYEkZFWjRLskx4GZ2AG+YU8PgKKgsTruS
ruiSHQBi+knxWZ4X564wo387xWO92z8SxWTQHR1DkEvCbDgPK9Y9/3xryFV25NU/ZQ8ubn3grpYq
hMDf0xcvZIEmAq2tYwRPC3wdAfAzbdJYud+8RmncKejCkkOxdlyk3XfjZqrfljnPG4EHhLka9nIK
2t4Hf57CHPypvlsToU/PaY3/xhry9VY7W89kZtEIWsjytZdSjAhjzsTUQOMOMJmvHOz+/YLUtAI5
66vJwkM6JCgwm3+OKJrQvp0nAje48zVroApY59YEgfg/uDa6t3Hqbfoj5HihYlS4JzL2HRYZZCIe
crU2K58OUXSIZlxzmngG+JlFRXpNOH8z62ym6GtWR+yyiWRo33tEZHiteCtYTMu4AXcN8Xpe0DN+
0dYrdzPjiuy+WY8lW8FRE4ikI0p8SOpWEb3S1lrWhHvIQmonwsKDLGe1Eo01pSe9FMIo0+YU5XVK
nlIK9poR9KtwRd6gdiwjzPR0wD3afuFXGlDH5gYO1LBYjXGZvBcntIt27ZvW3WZHBN5uU2k2zisM
mtcAKaWnWQG5qjudlneN77iSjZAI1MtcA6cYt/S4hyeyhMtNKUTwVKy+rW0rcZ3kBbUZH9MIGRqQ
H0Qp8L/GEtZF3IyEXiHRx71aFTYOt6+bz6Hdm3B/ShBqDhVHaya0ZFRGSmW1rU8gscGc4SrmWLS0
i6l8OBfodnmN6kH/B3SE6TQQKc0lItrLQXHBmn0At2+fts/zbUvM5wvcLWZt4q9AJz2YpbL2n9X8
5CzYfRWwdVfE0LnMdE5p33qKPFa2RJinmZwH4ABME7IWqZ90yC5UnEKR5WcvsWDSGPdCClqRWD/+
CM+Qov80oR446tdKhuSqrJjcre9XJDy7bjZKVvYnNu4D/uD+0fq1RIS3mocfOiRn/JqFz5FDCE8F
TNzf3o8eWkIaUZVI4DvKFvEGOIa4pBIM0DITRG3hUsbH3VWpzdAZQtfS6WGS2EJTpqA+scQG5GDz
HORMvqZzm4XHPxURJscXdyN3/WfAnQyeL3Dmp/IC4WOZ7z8J/UFeWud51FaImg0h33Loxk8Zn9t3
yAERvREBKplkpTVCknLGP+QAfbbIV5/UZGnTAu5ztG/1c0KU5F/0s7ogtUZvmAGIuVW9g+qvo0aH
JOnKpydL6rLinFCVe5j7/swii/gTqhP0DHsEW/J1kxJeiPZL1isJYQORd62YCr+Hsng49vDiqVWc
Eyfb1xA7ELUVB5y46vf3dNKfomB2ygB5+XMsRgiXgnwSxZJQio3/43m7Nhg0Uw2lCuANvDKa5xzU
xmoCma6yKECRPp7WD4v/QHCqcDY+AewRSo/5+0YvwCES+34fEpBmnnQMFqQLD1inZei31P9YtNbP
i/LP10ksSlAWHiapMsMwTdM2F0EYgek4BGPW3ofmM5/LlMWdx9isYWzeT6HsWyUYJ0T9ou0wSQJu
l07khX1zdjYAnabfXH6FrdOgpu8e840xVp1F3jSLHT2Jc/o+bd1xa5x7zqg1O9FZUkQQVAhja8yE
7wNl7x895qFkxfUED7DTWoWAKAlD9HjW1EYdKxJ4SZyfTFEIt8722SMYbfVzfP9XCck4uSlE/C42
3diPFGUKAt5XcRwKBKOUnikKQ1hKXVNN3jJf5fL9BjB7K+/ZsxkYn1aApQIerxS2+vfRb9vnDqPw
T3FsvucCRpxzxaITPydxA2G4wd7yOt4/f03ulUFEHQtMnV+iZ4zkVHg43jSMCRqzpekP1FiwoMWC
ZQW4JHuKj9YWdmpP4pQaYm4Uk/+9CWwt+cUFDR02k258QAojjV73rp61Iwpte8+ENZdpWJ2bSNSW
fxxH8iuy04wd4rDpx9l1ljDRvvcYAoQCLunqk1+FI+kH/OT83qRX87DlPncbbzWK4OFpClNFYrNv
jIFNt6d479dChWuJfpxCgIYt0Ku374PGgl4HEE7Hi4a8HIj1Ync4R9eHh6kTxwLrYmLSUg6d1NoL
yN5gXXiB4ZS047owpcw+rrl/f6HfI/0fOqwuzORr2lIYQ+k+cU3MOrQQMBiyywdLrACWEqfyBjE+
ZFqLrcuS74VZ/W2kZofm8ZrBxDgTixAKMp/ENoqrj9cTol9rnLoYgLopvUf2zzJlCtnEkhZL2bVH
bXpo49DkU4W+560djMiSnwHFbtC84DRAddo7pTEcyaAP/gDto399n6+TQCvrCAijn6wdgJE+93uh
TQizvzU/2XLyUtDGZsUiE3hismpp6ECKwkfg7V1qP1r7FBo/WyiFLqEPoTDqqG4ruNYBrRkLdT6y
J+Fg1KtyHfcDsqTtQc+yEIKNL4Oz+F0jjK6qgxSeN4rQpdebamyy74910BARuKVOP/JucXlZ8bHu
0qBhBsRdwIANwQjH5KVL0bTZ7CuavbPUrbJ8vpvhsPRbdyko/WsgXM9K/zb5Ecb/Tf8U9F/vE0m7
Otmy4T8kwB+hEftyUNMYtYGYkDc69e0/sfrLHGYJ3Gblx+GGKk2f0c2ObC8vUn8FNfV/MEcpXC1j
Y398VDWkWImROIyCoLENqdL1rgOf4q+OdlxLty18PuY3Z1s29RUEx4Plbauxa6JxRaLdmNlNC9lK
UKFi9UmxtV3k9AEsTa2VgiVZbIURk6Ib+tGiD9t0dglnUz/tKzkFOlnDS4yvyIa9n5rUH16uQ/VW
kpq8MSNWW844wL7j/287ERbELklWIIwt3Yq9wWwj5xeA+dCq4h/5z9/Am8RBPnxtsk/al+6M+PQh
rsqK4d1gXwhVAM74kgajU+jc5hJdE0vvQwZk/LrczsT0Jf3yJmN7/6Og+hRwCyQ226kO00YQWgMH
gCbmjR25/5N/LqKq34UdvtJ7QNu4cnBzdzK6GHKVMVomI55UYhhOkCntcluXai734ZShZUbdF1wZ
i4NUZkccuD6iBkeVRrw6slnPCYfATJyoFISu0NNp3G3Awd0rNG/Cug8nubfBIXRxmCFLSMqFjDko
dBXrCjVUhwvNVk8pEgZz+e4IklvbfbcxwWb/jphLxFIy5wMXmYlXTKcC4jqb9Gpwsxs5odrtnpz3
0ZVnfz+OYddIrjDpfGubFjpV31r0AqGsreWdDCQpjHgHRIzA93OxUSj+iFcN8cSVCQ4RTcncoKpd
PYniOh2ex1p4jZQvUpDZCz/sE+1TbuqVA2VaeMd3N4UXiUkym6l3sRyZ41g7hJyAt0x8FWau9NZH
JLEJuYOUli2kwGriSfp3b8zqHOdbH6GlOK4v7yI8CQlzp1seJN1QTcfjlozAulOpQV2epbkN0cat
WblvZMiTNkgq5UCWO9HmRX612I8C7l0nmHPsGWIthhMLP4tX4bZa4rEH9ebn5ETYYafjdkpDztQY
TG++UdpFORbfLvEYatECYRULIPoEAK3w83d1ON4sCeIoxva5dBCXwKRGkApFkyR0VuizR7ThheYM
+/xYv2VYheKUN0pGjVi9WeCIkaAIch+P2UA7rF/Tw79RcanMdnzvy4I8cTlk8d2dJy0AEC4ksLue
I2f6aPW4ynaJZWs6e8ERQyNDMK2wjwfymthWqRloTm+VwaW1MGEam5ma4ZcSfdAGHfWu64wCMSSk
HnCMzM5Vq8P7q20qpePJKdE0t9cl034dNFFPuL9KJtbpOOxsBrv7pwUEtL1CCCpj8r0f5U8efihp
cXKkYmSWj01lb/ub3RGni2tdR9RO6k18CLEJOVVPNXPzAgJLgIMUS+xNTGHtuFU1jyaCxxNRw9UU
27Ecx4NUWvx+jfX12tGOKZjK/NKwgDNSdNpqpTiEOTwAm7CxDILCbrp8u9RJYG/urFOxZwB7AlHc
cG6FwaU+zyv2XJax4V01wRyaEeyOlnBOM9gYPyUwEpd/6ZVo4FW4SmwAoc0jDrhkdqNiBQzM477N
vsjL61kLoeojOpJsoF12EtyxKqdla3VxiC52WcmXL3JW41W5euMfTB6WusGWqfSBfeuS2QkSxYf9
QJos68pWYjRhYHSvQ2edbtozKhHmf2Hc5WOH30yO2AS3PbSVx8H0nXYGxYi7j73wova71oSNwPV2
073YCh/lM/Zwd3wFhajrkas1q3mjGsnO6NGTW+PwviS1Dsn3fK/TMOKvpveAsVkfkBIXo4r7bbGA
BMOzwShXyWei8+106TjrDczUI7svmpDVBMQuPdpz3hoCuBotHrSwQe+LohikxX6HRKWzfoWHCkLQ
2YLrT1VpdiPApP4VpxIl0Kai0N9OlOm2s4w5DUrGG34d6YL/2hZwYWG1alB8Ao+d8LkfZdEhxcTp
DSSrxhovAZGerxaO1n6oN83N+n1LqHAVeUGeGfRjPMv5uSEgCDTowVKj8I3bYbo6fKZQSCuJdSVu
PKIJv3KGb1vailaXMFxV0r3N14c5WkGKTBeRoNnIfywA1jimwPSo6fFpI8cmNfpdgLx/cSpC0US6
GURezwnOCyfT7brVu+Gm/EF2S5GpnQQa1rO9tii0HxMx0TSIKXMYF7cIZx09hQrMyQhXBoZVqI8a
99u5AnJSiUNIpXEkP6Hgr5bl7tMFDybCY6bHFcgtrCWurmtk2j/V4SnnpT3PvblGIwZsC/ffNufD
ib0jZuPJAC1e2thgbf5NP0pPxnD+UXSdt3CbHK6fQFvryZbGA0ZzVH/EtiBFYDMB701H1lgaLE0p
9Mz+X4IG3LpgvgCTdgc82gQ1PK5+W0liAI+3oG3aG2Ehdna4L3kIxtnN6iVVLkNiB8t6oQ94LT1q
S0tb0buhgkt7P5Ac6g14bIgdgOD/qBsuD0Kn4tWFtfXdKgNAFpKCIzodIcZ0lJRpwp9nw6lXbhoL
LKY3xWC74gxBrsS08RA3O1h6VUmKp+bP1/hAZv8Q0QTlIoSK/kuuicJcG9gJxsa83LTQHFEqvzmo
dbMdjpzzRhk34toBCW9ezXfO2O4Yp8MSOnh1gLErtfFB0/Gj2uJ4PmpMB4IP5DYlKQd4kaUsNZ1R
KW5d566egq1FQZZMGSvmqqEjpj/hvj4CFt71M2CNuynWKuySDTzWiXENt87/fH++WuIPHmrSwR/0
/n/cPxC+X8ZyXDPJvlMzxFJ4VlAJNRxAyKZ9/4kpCIHx5N5Ogbktdui2COOtYv0C9rBXnaEbj7ZH
+6aapcxmrYvR+hRZAb8E8RHVymQ8U1k0S1Xmu8GV1501FDmV5AsPtendIvOet74pb1oBbKDRsVYu
T9byk2xz+nxK3v9qZeympZAEOdJkCtcRHTixk1o1nfoCZA9s02JhZUNz5b/+gv43VQHmte0maiV0
KsahG+R0meGa4Pe4P7w7l7+pDfIYAuZT7u3PbA+6VuxOZtA4Je/TzHQRiFjns/MbdkqU9v06KF0Z
rbUNNGlElrqlPKT0JqeVqBgK7eE8nds0KyT/oWFm6NUr5ZS1PSj9Kf+UGSFtiNSgNcKMeQD+FkHP
gd+Hwo8+1JJpUrL1lCD366GXUz2WicWgNvk0rnu1uMvHCAKOQWAGi7DO+uoLNm119jiT8aqhpikx
JwbEV/8+HIrPUg+cTSmMxligzBqT8AQE7UgyitHyj3cqk52Jk0c0buX0nm5jtMEUsn8zOybZyu+K
OpSOrER1mm3KXt0GPfWRjPMxXQRe6jUerQqx4FOZO1ZxevUAmrbP3sz0oZKcTsSE7K9WlV+K2noD
OSDR8w8LD4gGcMgdh7fhqzzHzIuksEddptTz5vxR/WaHF8mwxqYe2HGFoD3S//aE9luZltrCPoIP
8+1rZh6gQuNiHtG7D+YkAIZ6BxJ/dAiZBlpRnY+HL1pqP2no/0A1lK6GpU+qi1qt+5ImsWMH8WZK
tWVcT6js4bEgpGDt/yoITYj6LqN0YyD+7ym8cLpGYCzo0iXZM9WyuioYZjvP6KSDpBRWk9JliHkV
YpRQ16DHQMnNC0FUg3W9DpNZfyZww/xmN7Fukq67FiY6+zKaC9e5lBMkf8skyYqBAKMYDXJ2FlYt
djZt6fRQxrOHgsD+nmRtqsa92VeBCSoNc4Gv6xGK7cBl6xW3bRR5foGXztppR5D90v+WsUlmvvu4
r5DDqvQflZGQhiP7GegpbSJSmx98sYo+i1JgUPhDvyQcBf5lqL29Ts1JIgsvlGDeQGcjxIY1B5AQ
xirWOPjcn1vgAUrlO6YJrD9RnjIdi3Msa6eHgA9yF1tC+pkrfwY2XtqFsTcMU+wAF581mBQYLRqU
bK97LE/qu9xFMbXWH7NXvzn0IjilBYeJlYbUPZY6vCogGKSKqOLejvuYMH2uODV4MdPfj3WMhxPz
gJwPC/QomUGbzq44iPqG40RYnGQp1EsBUuRJ33IB7RuXR57JXcP7u/wXTLGrS2wRqdzv0MtTmHlg
Z+XMyqY6WcUs2kklUfMZrEwu6WuSuO07k1b+FoWdzu2vF6nCZo4yu786Fx1rWJLI6mjaEkJHxGGf
9F+jLYEAxtkr+br+tdc3sEObaKXVs/exN+12cjFTxSyp4+DHIehWOzGLATW1mBLQq4ZJe91Nmeci
YlwA9XJ4fAjYTjfHYQEZgMGPHiDWVJNue5HuMjzuxSuymrUnY/dWPBnLhlV2/7p4m/TjkDzki2AI
o1iIYLD5Ei/Gp3aFHeKoIVNUGGGgWmC2s2/APYxMmw7iXWPen2ESKrzV0udNSXnNs7C6phXKXcVT
t5ZpobK7yG64+7ERSdOVVqBvo11dZMZUNQ9sYxkvDeqZKQZP3gXLUtKj8l9bINsVlLq2IUWskhH3
SNrJPdquRyuDNZEIH6nrsLHz0SBeYTmqBh6pWxu//1mfB/iedmb+6HkbuK47KU1zjOmro4gZDOpX
Zgnvl9ShpfSRtnAe2/IxL4NUjGDLPbtv5ufNb4BQ5BF1K1sCFZjQQxsx5Pkbr5FVYAHTbopOX3bp
9Psq3xMZ4BhbnaXG6h/cH+Jc58zNx9tOT9RhFGAc8iuEuAiomh4OCwZDO4v2O6A1+9IChHZRwSlZ
mCyEMtmsPl7mFwVkXOKs3jkigI4QysWSr0aJEREQLj34nAyuiJQ3TcBiMeq7yaiYaZZ1f0JicoYM
lV++eKOM/oaRdNwki2ElVIJU1Ot+CEBmg9hIijcDyKT385XhaN8t5wSTZ/yAtw2PpCgVGWzitGk8
GBx045cAGZszQn4mY/u+lTXp4TbwhpmTrgsBduR/FLi0NF4U/lD/1rX0+/ngqHnUucnKXv8ycaTb
Uo84AgHI3JBc93YooEs1YsRiTs53nHMMG2GJ4nMlfR76yccjnDDmw5vwu7iRqSeADQ23RsrCy1Wk
R+98phJ1qM3vmf/Exy5tZnWrLWA2J5i8xnQQnt/wEY61ctsyoJoKdLO1gtGrnyB6twAFPGwAKp3X
+x+oWdpYwKFZXmj+9nYIUfYzNXloJoVtdQazYepoIMosT6n75jRvsmgpAlMMAGQ3LXiNC1KGp6BF
WGicZT7iQD8Zq2NtDl3mLDjVrAqce2/Mr0QWzatJjlog9q+vOKpQykmzmPE3wIKxSaBAg7aRA7B9
Ctc1a9Q1iNFEg8A7i8wzII3RQIMeYDotlqY9248e3PlFCW2bHl/bueK6kugQ/WHpkXyKXWtwRWLy
bj6bikQYD81dpTkIMmgGaWy0FHfsoaXKcKnjwtcrXCcDNmYWsjICPATqXcG/hvh/JadqW1YaPswn
e1ZNnt1Od94c40bjW0rAkhFNZWVr4zflcourqyK8IcKgGxQovztENNK0qeg9OX2/Mqx9gHgAZJtE
OfHNaOnmwLBWP9y4mTytVa5J2woK8oaIPPAPuo1PXpf28uvaLwIXTVpoqiOUQCesRK2B1rWb2xCF
F5H/75TEoJkoB8ntCnG7eq+NDXe0EctElvMk0WT7blrO0uXv8L+15DxmU7VVXpVB1PRx3efXjZFb
3c+YbqgNm4VZ8IvBym9xnid2uvA/M+jDBq7EkOzT3TE/9gxXTYIYwogZFXjcYm3Eko2fsQdjbzZ7
LtBjLthkM/fOv+9K89tRsEK2RKHnp70gzREaI3YIgRpmNsyacXdalGFd19PIN32j5bX55AEgyegb
ufkSz/eNulBlxeRfJsZ7Yodu0Mz/pT25eidweIwVuihV2B9TtFu5cC2428rXmkh/46WHIYM5Iedy
a5nmupmtc7w6EEq0jpbcUMd4bkTuzwDJtiKTnaWPzZXtTjrSPrej1J958ZCdkiAWXdyNP4PhFV1z
8O1LkjuL6ox3iB2SOJcrzIQUJVDfUTXr4rJalM4HlVQgAtv9/yUZ04u7V9F5qQtz5/bQUaYAFe+i
vIJyD57f6SsHQsHoWjiXpVM2JDU+pTxYqDnZRu9WthbnvxHzGI3JCYsemI+YPITJ1/17YGE0yCoe
s9WXbQlq2Ez42j1QVt0gBuxoIgusdhfoQQbIwlTOI9rpcS1Clozmutjj/MCyeRwdOdjNtFJNbDc9
AZNb3W1TMktKPJGkQ8kg/K5bcJx+1Y1aPU/tcYbTPqKgxmubHA4Jnw7QlW4UP4c23YFq62w77nSa
0H7xMRWsaHg+9UggV1BZLMKpowNILN/Z2dakZWl+lNGtOQvXKqvf+DCV/+xWnh2H9AH3/8+dS+0r
amqjErnlNFPEzJLmkzSuJTJwyE6vU99FxDedwbotB2+W/CtTs3oioC1bcBDdOAfR1bWyFlo9CBvD
5gXz2E0lqppGP2aavwsXUD38/P6jkrX0w/BF5RRnFv35BibcNN7J+j7o6e8DPbZr/QHMIYjfVUY4
M8Bi3s4L+nJcONUVXNDlrd8VgH7zivmdAafv2+Cwqu09uASJomMCxQBIYKyoOAHamBZObxyQduY5
Ol/J+6Cvk41QZA0PDqiwZYO0IAJSEgP0f8nfco3fYpHHuGZxeC0NGsa3uyJrsfD+FcxYPYdZ9XlY
cfuD/i9RzXPEApTtNWyQsrHyPx00hkVZytJiYUlMAEAEdnH50jyeV7lKjb5tmSwSYqKjpIoDfOv/
iA7WKAM7vEMxbUZVUe/KcUq6yxeevTgj1lviNLmHPy9KrufFGp7AI4yuuf4yvhy/zxdOoHc6t650
BklLBBWIp7lzwbxPGycM9X4Vu3cEtIMiSfrBeeBvd8Y0ylClIW4JOXa+sx4a1ItLeZq/7pKwMyvL
6sE5lq5MgqcdrmxjzwF54277pd+M7g4oEgd/pLltKiqDw/i3Sqh7RmPWLCnOOfsYjYGzUSknsj1S
MEkGjCBVv5UwKp1Kvh7ESL74SOx8Ie6LcKyxBrzlFu9YH2gNyQtogXdtUM+mnS/OsRLtUJZ/ahMJ
sz7SKINGM+m/cvk1Ad5c0uQ4YHaAWTPWCPM3fozaWFuR+joug+l1xv6ZKF269sGyOCenWZ5T/h8C
Hatf7tCsRgLCepqxgIOh0z3w8pzaAvWgL6FXJi/nxLgS9mouIPQHDBGYbCOyxSV8ErbJk4sG2/4g
mXk3+E1xsu8XfcimA4sEqj+5pVGWW2nWNWz5TVqGRdFGyRdtTkTJXXe2vuwomI0cEKZQdItq7keS
RoUojwEKnA8xc53vE0omnQUpVDmpiQVHC9TU4GxuzIWkVRZh6afEC3XD2QZMCUA+T9YXwZkUsnwH
tPS5kT3lhJoN4VZFNHCrCDPCyqKOXe8Iqjn0KfUi5MT6Zoi6LpgH68E4QipFzU7BppcH7w8uch5i
HBYY20cmRvS7MYOElTkWjnQFkKpKt5sSfugnwXzybKA9+OSctymqQnYjb+Ag05NaM/5M81iLXbyX
HUAUBQmrRhJrvQAeB+4RWompWxl8v2vNJCdheN6IXeOFtwHpw7HWIbPaQFOVdt1+YxozyrLJtK0H
HeJR+gd/yJK8r6AY2IOwwXNk2HvvxY1BS0s6nzdJ6qtUy+Sm7zSMpJNm6R4QeMpugbEIruww1ADA
F0LoR1BqnxmnQGFmnJk+qbrNYbvmchbbaAKmaINtK7RVHCUbSCKwW60/J1CLMRHaiYtEIljt8cPf
sXdP8+lkri9Yf/HLycNkSYogbjPMsO/rf8lGnHQUso35S6gzd+iVrOSGRxIEPXMHYwZNbOZtqc2y
cLdaowW5vUXRCzUHOyYHfb3EzNqNmE4FS+B0BBXlUObPSSeu2hnRkg1fFq/L5ijSEbgTpMsphDCV
ycm7MyDcxKx9Ssj6tuacQnIer4J8lpjWu58la7SkARvV0mURuoONpZvuDyQeJ5yS68wuEmjRPzrE
alaB8Tu6JV3/hGIAJwaTIoQMnXoA72aumEHaek2tTzkaO/pfujVQGznu1of4LPrZTKb3Gf4WgPFl
CzEjw8JWA5Z1sAxp15sH+BCSrO5Hg4lm8x1nUs4oBXpfDr3mAfvEzRzCTWdNjqCMWGSlshkzvtUc
d2vqISOaakHLjo1NT3tB+Af74z1C2ycleqirCdDLC4lFwuPIYQjtiOuBMB/PXhH8UTGJltTxKeAz
+jSVG0RY3GG7TbhvIP+x2evoXm64H1/FO6Xg2pKtBGU2ePi5vVDKHXI1xw0ErUa2w5U1Qj7PGysI
+3dnBGolzVTlBfy0vXZj7XC3Ne6rFifyGfgbUH/ddNilH1h0Obv+au+kW1KZHZOwz6Z1zBRhUVcp
YUMftsdZ0gTgEzHcBl/Qcufd2zv3FDs4Bc2cjmXXejpA7DVfzHVwmlCwTPFoEjzG3CFUEBWtJseM
RvvX3vPs65/FoI593pl+Fg3bwIgR3LXgt5uy8LDTjLGbbVlpt3FxxYUI2XYGIZx0QS9UkN1oN7xK
bYXPlQFKalcEsULkr+ddgcPM3F4t/6uBa+f75zdpqSApOTARz5zUa4tjmW9rv2UEwycDMYxXJv7j
LXriuswz92KVennGonqSzyVVHuvQG6wOVzXVmUwN6MpvIg5sMDWJFbR9JfGogy/YGhRQnzv1NFV9
DodbfEdX2fzLj9K5/gutLe5czaPdMJr/qx5VPaAlpMY+9HHRVThrBNhM2qQ8OVChFxmTG0J0f6iS
BC2aCC1dyZSgCewI1q1M6lAxldWa9TSWtdFfqfSeyQlAP5GG7n/1C96k5nx19Nb2AjU7lk2j5sGB
8UglcrAtv7S+Dn509mx/MuyI8F+VlRKzUmsU6wU1LXQLCksSE3iukqGzpAz4jxF/IXYhxySYGJTG
pcdHFz3D1BCCmEnfmvanj/zgn8lu/GHOOByE/ypzEPEMTUCXkL02GklqDwZFd4QvE/LzsaWAWAQF
0u1c0ddUPgx6RQ52WNdyyBNYhilKAj0uHU0xTwju4mcwLqcXr7feH+b7Ts0nfTB7RctzHt/WQbvQ
AjCxBFOZwIExL2kq8AhNe3Ax+7hab1qggORLhoQK3no49lVBNhQ1p3g8G0V8y9Y0xVc7H4qjBB0e
ZAMzuRGl3oWiw4VD/gdixbFnl4lEkOFyfCWiKNBBfK23+OrxXdbQxwLrp1V1QU3wm9HFXZlkLY05
rJ3CDC3UQaGQXWaodQ0yWvJsPTzZ6v8WNVWOC0hBrXRNfIUKkclpS7oKSnwtDCut/DQWGnE1R7rs
t5HHoDRz1AJIidEqh0rhM6UvLN+yYzvxxAsOHpAHXOHR/ReQQmQCvv9nVgzOkQN1emB+tPJWqd0R
x6Jr+bX6nwXC8mI1DVHQMVmv56q9RwKUmyKiO6JKotM4TYwn2UxXRSdAZDpEIXDdv65pYJTscmSO
X60GDcSdnglgt1+VwjSbq+73VE7PUQdSUyl9sG1AHx6FTjlY1gr55kl+3WOfWzbwujQ+Z8kfsGbt
DpRRpDVBp4LXLcss0gZssCWRHLHkjbqMGvYPmY0hM5Bt5pY4JorCkg5K1T77AVhJoHmq7eSGeJGs
FvKb1RFxeTC5/v/REJgKQsQj6Ir7p/eo7Qfgu7Wu4TeFiHG8u/6zHg/Hjdic8qjjK/8fv07+OJkH
LtX2M5HdgG7EJpXv2guQXouEdKRUCITEm23f0mytBTy8Jx906OhqmdgNQzfZb88AejK08/MbLP7O
6sxk4m5Og4Axymc8lZZmTz+GzWd1S5NqDpcGizm0lGA1E6tcrKbQ2FRyE3gM4ZePqSstPW6YY64V
mXLFb4w/9oa/UY0hsFJ+TzhsMTdU1m6fUyJSLVhx1pQCcK9kpMBrO3rzQv9JvqIQPkzYeV8RR+TF
GuJ2YYA+aJCxk2SvbPq8gGl8DBp/LcoXR8TjGajmSbP5hI8EG4RQRXKBeJfyFucN4oYREV49IGmx
+Gy7FuzyyiZQaQLAys3UB/nLdv3aTf+fzJwnHHBclRZYt7Z7zc9p49raD19agbDhaAtn5lj3COk/
G7AiqP07z3z+8TnzmVIX8yfVlULEC0O4d6GxAqXV9pJJM5VpLSRn93JhRn1LXyg1P9ltODJtxJ5a
cSkGJgX8lVApyVyl0fIZjMyZBsoi8ZQqDkFboUA3SNfcfkH/O2wV0ih/Q9YOOVm9e9wjP74eIn6U
O7m64rEQDl6CUDXP938h/04j05yMyFwV2gZr3L53PYD5RVGoCpF86kR+093ebpE0IGM7ECE9QiZN
h7j4dyPsa3wn9uAwRlsJcBxD8dNFjNI5plHImShfSfPkX+/FJxkbMvw/J3utwmJUrqo8tngSzqwn
yUdQai5pqTso2TUZv7y6/t3B4UPzuGA7uaA3rSySiMFn8wlKpkO00llNDV2PMxAjmvIAjIwE7Vjb
KpqUCq0nRD6IjPqQyXbgWBcCAvltae6gKNIzUxB2sL7520IGAcQmUcZ9aczovhTaYy7AuRfuj9+C
7+A5O280M9vBzfY+vq/05sxPJG7gikEz/MRdSOItB6IdCtrCH7ppc0HCzP0Nb/0tYLZzcD3ILnOU
5ypHZexmLKWPEZvtf/ev1G7JW2B2btsmeAv0bnowky5auc6qDBsNjOwpB1IRvqCH7d8Hy3cf9/Ld
3sx9ibjXzXhQ8FOvx2uRwJhOebM9D81GNWb3Mn9/IOG4TxdGXYwRkSzpeNXLDlMsOqKOEAffwlAF
oyh2WEHmg+ZpU3l8dfHP/Fy+X2GI1EBx2agPDt8XgtPwfXeKWzLryjmdnIbxZyXhU9btIEZ693Yr
F3onZFVZwQdyCP5X+ZnztE1+j435tmaXxBxX3qeDupzCTG8qvnhpYkZjiczRi2v/DnxVdCKiKEDP
5SUeKQ84f07O7lKYtjdbzIl1Aw1eXotb4QPWqzPO0jy28UszUmmddl5Cyty8P++dU4rbBKdmiUsa
jjnKh+i30p3RGOCQavxLv8KWPHn9VLSrmVyawP4eFlQTskT7OzDIrbC8d1HUgBRTlTkPLImJcqGt
irRcoqUCJ8wsu/R0aT9PefK/CzLGW8Z8CxAa1Z/QBgUVPytgpDgvhHCrNNVtWu0Nf0UqG6l0Z8Qy
D5LR0q4GMh3ZMHZo6OhpdD34a+5wffQQYYGI2dDndvGUFh2FWYu1PbqcG2adg11TMcTubSNSy2NZ
jpad0oqEqwYdr1qvyHYqAvysDQM6NvDxFIV/2u05X0e1WL//IHdXJKFPb/lIE7qBrHbIcVtYBCoS
3OaJo+j2zBGuNUD9JsMEkxLEahQ8K+NOFj8pvEfAlg6LX6FSQd51vuO9wdTsIy0dv/+vTOiHBAqi
/i5zd5R3I1FW+L2dCzX7ml0bdUlyf2XCnDcT0f536ZI1fLlDR7NGq+EvwImQBtEcGmvKPB1R5/dn
lbLXm9wRgTYQWivvEWKy2y356KJuhIXC7k+FV7KinjVwdMisLrccFOxhoR/QBS9fgjmgQrJ9HN9A
yDYD4S0X8UCmxfNf0vZKMobMUYoggRkNjXB5Abu7SuYQ5QeTwtVRthtgH99radzkjeNaCDu7Br0b
hOCBRpIaQPqVF2OVxbqp5Qf13n15vAd72vovDhHprqDYvybZ7seF5UY7loE1zFqpGFoKlu8p5a54
jswl/AtYVQkDcmGE+8i9crTxDlPtEPSkh1PQAZwys9fEGsg1uxNROy31gYhkqYgEUp2DUG6VqKTA
OKH3CD7nNWzknLMNY3GSUWRpznJUzXcxdUeYDw9mTp65NGnG8ag29PbcToWtbKEdzgldcUMeE6nU
jRdAkfCKPkhxHi3WhJT8A9jcHehMpw5/6pEJWN5eJ6K8qvO7yraMN1VNFHftCKHfAJDNW8dMxTgZ
WOA7rrdEr6nVnGlSeaK+oMNE649DJ8GBji38ORSDOGEMW4QSIWhah8nWPUHedbjNjHkw9vFOCNue
cLvs8qWQalji3LrnAsZ3jQoCHgcJE1jnGf7985/yOwMcIF0FfLqEC02lduBBjjIs87eO7iU9rN7w
5lKMCUrizUFnqA9LtjcpwgMQHDcYBDYPHwcmIPkSdExRUkSt85RBgo/fJlf6wlo7aIenjPD2Nbms
O+Z8KHQA5+cc6Ns3rPBUvReGaXJRL0xbuKj6X436TaQIP+unk+8ilc9/wT28tFM2s3I8u3PMBeNS
iRJao07fEPCGc5vnScS/cShJ+JkX5CDkjh35M6qxFyrbnRuS7qj8bRN+ZWICqP4R8Lsft+38aHUn
mizF5L/jxLmlEiy+u/luExDZJdZgWoa14NynXP8TQZ3HYpPAfBANmWaT4LLODmeiDAr10rUuk26B
KHoYG5F4JhPUPbZBLzWTn3tcZhGj07qIRPJpWOz3wldAzwM0u7+fkavmXtIKp+g8O58bTCgTHphC
4Ft+RiJRt4rnuBFbSa9KG0FZcEfZ5jrCsprlDEnkK9yT19o3c+IaJ8TQOqRq29oirAryELEqMhvj
GtDrkpMKBA/DUbFOr1OOvP9tBUk+E2Ls97yGgKvGfdnWqgD1KJ6eGIJjcjrIsRCknPcrwJIshRal
6nJnKoNnpO7MnFlzTMZ52P5cIhv/F0acGnWQkfSZRgql5F3g2jDLLkvywsQjPD4KKe78I1pdjl8k
0dEAgMRw59+UvLbmz5xmV6Esp9jGJt3j8lVtcZc6tNqLw3l8MsW+m0eT1o3ljmEDPty3LkOf6nUG
QqwoBMyFsCqHAxj4VX2e4FuUbJRM4pqB6/enoXtolmtVa99OZ51xmkgnBXPdBBPBM+zOH12aB4ZN
/IO1mFUyT/gXiJdOAGpmtmoNYiatGnJmrbJlvp1CCwiSZTu6Z5/1pVXE6j5ChrJCTAOo14CVfkaf
K8NE3odf08srKUk92nyoIgUFGjm02j+8zsC5voUmO7ov6Oa8QdkxiI4PF9f5vpgpcCt4lgXN/aaZ
xM+tDdckACc2OAQEIbSUxoNV4gw+q5O55YnlNEN/5yJ5a4f3ZlATFXBTQmEzULKvylqcQaa9jMUq
HkVYshtN86BrJJIOuDQabrrOSZ8N3eDvi3dk17FuCPpA6LvpndZI1CJoZxBc5vk1WduoppFpbnrj
iLgUDRvpOFU7b4iD5iLWSHUoUaF1Uv6gg1uc+qpU+eTuC4NQu7gHpfx7oKyzFgTWtSKxmxuZIIfj
ReVRHM9+L96SBp7zOzn8BL0duMqYvcyT1HSzWe36wcCIpYHsDlBsGdSbaeF8mqAVFOp0NlXlnMkn
jLSIcm0eX0Zt7FQHy/ZKGL3A50Ycxq9rnxngI3D6lwOxls8eS6kIhNpA9CA+ztbjIUmBbFlB3JU/
Nqcl2Y46ASUBoswFNbeBdD/cpUvrvOVZadB1WdzJt9GbcUKZ4s1qE1DAGDq1csyfSO8cGxbG9JJa
/8P67MLrNsr78CxzxWjxv2J9/rZXmxs80uTf38v2egV59suruDLmliqqQF71zG7Bo7zmg6aJwrIF
JxbT7WU9m3Y9m1sN/+OI/EFDf4cr0E+5NwiTUgTZ4vgypKSavJ3zPlsuFgUabU/uv0f2DVlSDHzY
wsxLkmZPHm/nEp5G2zbSUboKFy062OSQsiYbWhJVp9pmAz5eROcMI+Fn5CNl9diwH9J99P+BF5iZ
ymqxc6gbGiPEhKpxnHhPOEXGf3t9sCZonvAT1PAiY4o59yHR1S0Nrjwd2nBQZlkXAHELMMoOKjx4
2WlLl8R2eBsxFUc+/X4fM3rNMKqtQ7WxRdrmRLrsG6VnqFi3rEWlsj0K8HhGCXhelnz98JZPUF21
zeOAtQfbf2TX777s/MfBmXxPcO3ZCJaaAiSpqm+GIAGwfDeXaAi+8N1G2T3+mk1Kgq/sJi9gVeys
fA2L/aEnz1KAF7EL4W4xKITxd74ib8Y0CYhxpQ6Cs47uz8SkppOiTDkMhY6aI6Fwmvlmbc3x6NIN
z0iyb9lbUq+y8MvuUg7qnhyiLzZuJ7tq4H19YE/IaiIScPdBgiBwV+vs8jJTnKu9z/hlwlw/Ycwo
vj4IayQs47cjLmdqTUKKaMOwYH9Rn44HzaVJrg2r6n3BIQjZRDeh7smlHWJNMrtF3LHcDqnwrZt2
6M8V33xX5G/xHCqe3tfq/IPwXwYc6SffDR8AuR4+FAiF3/XUeQQ+RBsyL5CsH8jrZAPu7FEkbgo4
6TCeaLoo1bJmf491t/joI7pckN6kMZ/yvhFLVe0q/acQR9IA3LI7ysEbWrM+vr4TbfQdPN0D5exV
+/B0ABDtPaLnjrCUTn/ROIhgO4nk/BFM7NMJtaDyqAdi53cxbzVFqUxRovf4DSlDPK9S0FvFJ25m
F9CJXhpsJkjprN+D7LBIrkfhs8QyKHe41uZKJsPFzNeOfirhft4+/58pSyHZu5GcsYJP3bSXuD4t
N4glPwVvP6IqdlOwuSS+H+SWr5d+1ivDrWrlz9COadIEMCmGX2RNEDEf5Gqt3Mi9dQP+Ru0FS4Bz
w5hScMszP4lu4gYgWfndt6aiUi6IGvH7GJQGajyDWFkY7pIAzzsuYqA5h0knKFnRYAuZ/lnwhVqL
ADlURO+Svf8HlPLveElYIXZZYMFfT6ycT0Hnzwapgh3VAdWezYd0LmUYwpPL4RU7jim20yF8jBT/
MBBkHpofyemjLv3Sl6lSdHVbDNSP790j5vs/ut/LkRQWcB2kya08Ki+texnmK0CGIAhCrXkJ/CLJ
1dL7TONf0TBCW0Z0Cu+MxGp/wclEE7nmFcffHaQKUrcchOtZn97mJknwnhT686G51pKrYnmjZiyQ
rsVXlPrshyQptP9qE7nokC/Fpq2GwPxV9RxN+3pmno3Pj0nJrcmng+lJinDKHSU6fl5NDHZKdmTJ
UBc4pI+SMjE5kS7FTXEE0O7Eu1AiaKv+efJCgIWZ0sc7MpVMThu4Djnb/vZPi+BSj12DgF0Vuu8l
cDUlR3ilq1ac8mRqnPn4V0f+tdaIc6TsVuhAY7eLrPXD/l8Mi2cABS46mHKMRxXxK8EmjYFeHJGl
geeW743NyVSfa1itK825+2lE2X53ZQqsgZ/zibl03qx44LafMYHPig/iMNBaR9uYMTaJLFIfk5Z1
H773TUQTnApx1M7QmrtyJfWto2NN9E5siB0zInrp2jILzWzeV3zuVzfcZ1UYNhjKRFDHM19w7soJ
VWSnp6akOd8fJmoAoYv6/bVr5jgzx/vYlZKlRU0hkVBtqKIzBGbPs8eB5GxN7yCRvHmOb5Fdm76t
KtQtSs9SSrOic2GcvYt0FZRlAjnDFXzGsyiAohYU/Q6wEurtOPUo04zYks5VAyRrW0vXa4fPfHWc
WEFYRuYhQnBeeT8WA1M2r/yfPmB1PSFncZkxoUhIHezSpViD4seQX3ba5Ts4jWUDjHa037Q83KLV
Dwy01EByGt0CNEXt4W2/w4kfdODMJa67KWukrcPeHtVKaQswqkCF5vNbi6UbN43DVAdZnY9VYoN2
sf3udiZN9xZVAb4QZAeJ6+g9Q2VxV+dCdDenwM0w7QUG7x3RF62lv10Mgzu+a60AYbf2lvnHRHbS
X6fwb6TIZR958euuatmZ7jiUE6URExRHXW/o2ZtNAcCl37kW7aTC073S1in41PrXmcXJAgT6dX+p
ullzuokkqOlmALS2TCVHf1RQ1FMBMY9rM+x5detdWsIIJ9MN+c1n/cezgBP2p3CSnkP+MKaBI1Ef
mJOXyadGkFs6QXGQTEN275oRg9dG8WRvwe+72VYa0NebX2eJOAQQvyWbnBf7sLaSn+++Z4puDVts
qf4cQsrz+2taclEQluKyttjYdAcpWpZJLGf+9uA0llTGMnD+ZEbPffDOQAb0iPe315Nv1bDRQFLJ
6cbKSTGCeLBT/6DS3DPxds9D7UWVZdY2GzoQAkDtyeAl+RIYVDeYuWQPz648bi72hwV0/oJUDF+4
HGFv8MMuO7nLyZIikyAqSSZR9Zk9l2mPtmaSKVeDxW5ate18QH0oFuyK9zdmbEk5BIU/UixAlg2/
PeVSVAJdkt3PLJupKBFf7eWXlvdaJX3HYseWHscJVNXd534s5MgYuf6Ff5hGFfafrdLEiIQfR1MT
DwT3hUWvegj4DX6pwIkGc8B5EKfbX9TupRoyuUn7Bblwnfq9xXfSDGvGGLe7ETgK8jJp1xS+F3Tc
2IN5RotbAlIhkIfjidKZoF12kfrbGQJ4nOcGMeSBSgWPNuULQgb81Dowk35wkzbZKKMcr/eKuc23
T60nOyEG1NdESjAnuw2232WLc3/fy1d+ItrKP0UHXlIuH9l/seBIRTVZi3B/QeyYPMZKboTYdmnv
gogvJY8Ez3ZCTNGXgSg5sb+6zPo+1wqbOwt88qURZQOzh6HmfjMyeBprtCdcNj8SSZjcE0k07bSF
XCYDqraLigaqK63ElBuvRsmFLLAh28QvdHBJcVASSQ35vnyDLxTHNSKYNTYV/D8dolXdC6cxNWOv
L842NPXCC84cO+fcM5BtHmHmTL8/ZMZW+dcuYndTW3a0jswjlE8Z0DF+VrD/AP9ekuhoffI9fzOj
RPb+pnpoONkSTrha/TlAtEQEPgGHHXu/Y9j67cemtpweRp++RMsrshw1P5IiAYivKY35sJHcfNwb
SPltSwvlkjQNvtknkTZD/liexNBNL4s3KczvFMvDfAfGJgYy7/D2ofW2aF1RZp2bga4tzxV5W0I3
rxeG3ClkiucijLRWzsFLaJQTNkT98YEvo2lNy/fR9pjcHBcBPhs41nObIuhfpzQb5DX1SNKdB3tE
yH0m8RPvXPX0sZ27Rk3VJoDUVbIXPKJGykL5n5fAcJsxkaGccf54LGYW6IbttFuBa37bWj7rkUkG
R8lx+6T/7hhnynqGFQK/W6BEnvPg+vtFa8AuzRKm1G/oGYtyUz6E8G/JFIqsfKKfE8JHK9Uemy5D
jYi7VL+yFpW1i0mFd0KSQqOJ/cq6R6Tqwh+SdzpRzg4sK9Y0ZPaVn94MvR+4UJ9+wxdAERwZeHiM
DuXyXkC9ERaoixsUyAjSK+ZSNlafdpGmRXUWzyX0ys8RrSMcbBHAO635USiEmu1bVj3mUhgccNZp
UghyHa5wQwunmX9tD3UjBLhOIkNiH390kMl+3AALoG3ftAd5r20eoUo2L4sUmIjm2i3r7LF31qtb
FOKhi0xeUQUv+/Nn0cVOeoixbxvPvmr/u8iAjX2iQYtP/vpotJmFNbWh/SYwgEGPpI1EBPQt0nKG
MdcFxzL9dIH805wzIw/tdz1jOmCRu1lTOJylkseGLeZBdcHRMSPKVifmTq1fRPw/eTPLfmQtB2Zp
fVJj7EfZ1VyiyHLJlMTW33aD6BkmX/+esVRANUkrt7PTD7oprxXrJ/3yHgJuMJ6N4eDsk/tGbxfd
3fq05EcyBWoqR9rUYLQrlGwsif3ATPuFGddkL8HsVcihyo2u8I3D8Y9lTwB1e3Ty35x90rLQSEIK
VMSOh5ES/YfmwC9YxhYfrC641Y5mPBV9HG0qKREyVkwxntbC/9tHdVK3v21Yy4RIryAxh0Mz95s7
Js0mHjE+bmHU3makLHbJYvhW+cPAswtgRuzhFMSKRxYj/FkrkNBOLD0RacLk7Zm47IYa+mOEtbyu
LbqMZ6jNcg/PT1yIJAO9xhsOA42gv9aeQOyD3aQj+v+Ak7Hv7F1Qg4guk/LaM4rvKLpOKkhdzQmS
aUYKPPMswB009YA7F50WdwOGnqZprA4LrElT07Msua1qJnLfKam6NIZIWbfrR6fWu8VxdQl6tcnD
Dz7gu14qql/xioLgt31OBl4onfy1C2KkQ6q52BeCmNN8hWMrb7NdqK2o5QM8KC2zd/lCzpf3KTie
/VX3MsRm/c3p3CaTRJjxE9bgDFWMs+v5wi4EWmwiAl0NBJXkMTvBsTKICRaM26OwO3wDw7aH63jI
SWLsvmKBEjjvtzkitWWQ3zMDLNNhkGBQiTP/7e1Qf01otkVNDGf04E7AsbR5M7KMox/mmX8OJmNQ
Z0pwClB0SWo0BL5sYNhbemwxD1nzWa5eK2vivY2HtMuGcqQ5TZPNOI1qILULEBv/rGX0YPG4Om0B
fJwEVlWo5lb2aSVLZMcB3p8eoTO9BWSVb953LXfV1xhTtD6aN/VW2Hx+Gqo6xetCBk3mtoQtr3xp
d3Q7asusad9eRPA+uzLUqNsTshhPZhWaOdqkR0BaS1BjsndIN9/g1aQoSLKyYQwHF5iWmgkSzrJ9
agchf5te3/+GajKIIhKgyIuoe6rzqi8V1GNFrubrK8h/eLDoQyD62BN9hSA6BLSQ/IeDyhAE8FWA
p9kVtRTaW1NtSyaHtSYlC2PTM9xauwdFfO+n1PKiQsqjeDaHQcBlYpzFrnjSod7tvqS6nJpWG0MX
S5tf1OLTx6zivbyga6R3+2LZQKmN/0OpjiYkeXpcIkdFqd6lNcfmnVx7M7lWRXVIYGXi8MjveSQa
G8z/9x6MZuWcC1ER58JzXj0ZLk/4Lict5islh2P2wC6+9gGNrR3cZMIHguQUHvreGfdME+pcQnkP
6Afdv1k3rQZ3a8WNKjP3Fk2m3hFs/ddlBrDIVnViVhoJXxk56FVVb7idHO/EHU5TZDjrK4crWPJ1
fSV5w7MV7fxzkyTH/NVUtHbLA2HAOaLDD/rpvn26HKBxTTxLrcTr8zhL+PU21PW4fkoh/FIv9l5M
j17w8eN0XiAxNnDc8DyiEcaOJswJE9pC2bSRHu+NusoL4msScrC1567uuYrluXns6p+QiROj4VfF
UVV0Y4n5eau0OgsoX3a7dPBvh21xhar5ZYFhHuzAKa5dUkauHRxwPJAHhYYW7yag/MoLUstWvOkn
u0dTsa5ZwdrPP8qU62f8owmfE5TNBvLThyu0Ol8D7/wz05ZpPXsLJ/B7nfAYShlTwfn98nzROOdT
oPd1McPgehcExLdJBBqbn+2wWc/WlTCn6Xsh0m4YIY9ljc7xuR0gKJrxyU7QqfJ1AZmkdBSqYkgv
5nSH7pXcCRY7Ky9+FdH0iiUERk8e6au8sJY7pv5zRe09klsEKwQ3pMMyfdHyBBrB3haGWLuJMTbA
nus+eS0k1awoc02vAIMS45h5kGzktX7z1I62E7ajTEgrmS/gdWK676tSQ6mqGyPn9EBjlBTg3nSe
z4h5F24B5qfDVoMaK1kXnROKZ2oJU9+eRBxNDUwzOzcUdlL0LESSQ+3quHwb5IqRXKPwO9NtdbUw
JFiXQ9Lqv5xIfjDcJDctMSnmqPsbleqbf9aAAbwLqidQT4LRbD0YvtbwQVE+1hrGZ1C0xpv1aEJc
FQ/e5ZNT8/QDTlH/L6EUt2+FFljJQwiKXL5JEB+qBlD/aX5a8dGSBBkbMxkbyecKzY1vdn/ILadD
4RBo3Zi+/UnWeW9vtNHXqJ6E3Pw7Ow4Ld+CxvLOLJQNPTxwrHu2/FZAjKOJGTTt8a/Ahas7Sq43A
yiBPJOaPmT8Ia6pnA+dTfnqtsAuxTqB0Uu9tSov32qlrx6Y5f5NVoflKKwEpznWH+fqq27N1TGHr
rPCokfO7B1B37caqhel+sNtibpSK5wvH/Wtx4/rAVs6NOCPmu23EJ+9f6qxJdB9th7mxSw4EK5wr
ars1tCYPgweroznX+u0G8QmI3M8uKJv5Iycs4rdxZdo2oZS7IB7/tcvkNWq0AhZp7guSqoIqIdj+
TN8MxaK/qGtNTh/mAhfAj+rPuyTxAbAuY4//ATePrc4onJyJ4OsBqFcvJK9he32dgt1LSLGhNwoN
M8v6z9ZDcCoZ5mIDSfOOsX1ruSD4u0dpxY6kMHpCH+xSiLLBzZ9lshgNy4ZxyePNdzuGFeOIS78b
98IyCpKsWvubod3W9mkHvCJ3+Y406CuTf2mGTwkV9OX+g0E8p2wG74N7PastRhioQw5veKjsWQhg
P2RlBc+mOotxsZ/j+C9PhMIzu0qwEegDc4N48DXSSqcsDCz80OzZYChGxmb+utJMWoFvy+K8fvSN
GBcAjSANhI9MowPzn/T0KJs2aYnHzj+toDCLrveHDu+lMQQiSv1EiaMBvABqndq58uOeZkDfVHq2
8KaDKwdj/idrdPAteOXHCzbTHNylqvhbvexxf5vkhSmLNmL7Ba6drCAhKXkaIwkmbzEGUB6riK0I
YW5ZxsYPTMXmgAyq41X0+Z4n2Ro60zvnq//9Tws1FRGrG9A1BYOm71yJy1cihq3BynSx1B9edmCD
jS3tH/DAaA+CKnlvsINXCLiwkCAefptZu4qX7rB77hqZ+iwENg639ISbSeoyspKa4OzWiDvQ6i28
A/skaLzUFPE7QT5/cvJQBatHH9cK7tMOl38o+iREHXlburArrwuMOFfYqzgtD5ykxW5L7++d3KZp
i2OVDlno6L0efypxVKmF6wa5kTPq6m6Njv6jo3/ynfKXSh4O14+M7Y0m4CcjbgnlomvBiDqwE1DP
JMfMBwvbycuB3LXWgAfycIOw62JRWiVpl54fz9UIjB+hO1EUIAG5c9JJpvFoiq6l9Xm5xBPa4CRV
2jtvaJpPwI0Be4aPUlXdjWX4RgkPjrcaiob56HsWkBC92HigXa2PLYWxVKZxVMEVI/tSmWoJpEJ8
AmEgJ4Bv4tFuHttKrSM8PwSN6ljU63S4z8L21t+OmrXAfTE4hORuANVusCOhb5rqVfLcfKRWAwJ1
4r1/yAbx479BUws1d60iv9REHKDW+1Kb27oDuzyfO16qfifyBqROWMooeVqrdD5lDMo3leGmqJOn
KqYtcR6AZ9Jr/MOZDJHqDaPqiRvI35arf+ZgTP118abu1eBH7PicFaOErBYuJGIkSMCwlq3pmY4u
AJbK0MyuIZgT+EM8HKb9oInBeFvBmxq4iTJkgIGu9K3eEw6T14oANrsgKCXmFPcTTIiD9j0kY+nf
Dult/bOinDtIsEZtOIe2/BPS9wV4GAKQmRSZSG3GIdfXhL2df0KDeTKxvf73zCHNiABTuY1b9Izq
srjY1HoNM8HhHrFJugylrkvLz4Lt+NztF4d97S4zSUK1OcQCe+mwHI70ip22txclyMqkDgD3MbqC
XbQS3KEuEnP1PXdsTewCGqRLzfFcYlRPgTwLBYdmULjHv6/bDCoeLn6RJQKDiT/1bLjThvHBTSGG
6cBFOUu2AMiuxHAhpNuf2pX67zDQw/47ZV6B+eS4XulZ1nMhWJU2eeBIuzriG01LLfzXOY3ceyUz
gqrKtLYlyAnNKlBF+Dyasn9eM8KSWgODU117nNjpaHG5F1l9uitG3VpHqi+PT8hl9r/kg+pLNUen
0+K6fZN2tz78TlQJ5EGV1k7sajB/w7hYbMXtNgT3V0KobCROJQD7wBXjbcOwWq8dlvYI0MQGQPvm
ZtNnQU9BU6e09PS+TjmgApF/9qSZ7pm2ZFVAcCAuCirp+i3YByZvMIc9rHXr6MvH3UskhXWdq4ex
Fy/efOVXBO5Q+Yl8etrp1tTSaG/i6zYTUeWYto8nVB/Lav+7yZOQTCmYg+hq7xHXBVAQ7HVgLWBs
uLBEYFOUtl4rd/GbcwsyKtk0XfF+fC3yU4Y/g5pR4nR2S81HeyjLD3qDc3khzM6griGbcehWuSBb
ezv8k5C2CXlwiD05JdlRX+67MO/6ZGSfgC4+jws+ej8ubDba3RBiw+vN+Ol1Lkfn+Cn5haIY/0n9
hQ4bzEbyUj6NQeGFWqrYFBeFMlujeFuTGINfm4fuYhgNA+yQHKmNLGGi4ZfqWiCu+UyKNuPpyDso
pBcIlIIsX3XHqzS8VcNlvDVHT7kpVPNzdTCdURUXlm6zBzY92lYrY6iMZD90U9sxFrSC16kMkqU2
XwWZWw7wJP9+75nH2s3R4HjT1VNDKhGllR77damib+dsJeTicL2RD54fOlf72YXuTfC58nw0KRhk
9cDPSuPfsNz7wKA/hiTjr1UEbX6xZ6b2iv7tjiKeNXUyGkFXwl7IOO6wi0kMX7r5H5ZHFFdl4MDi
qFX9GpBH/pMAGZC1x2Mel3O+VDrp7DgyXPB80LhLQsH6L0ZJq+vjAjXa3QlzsoPn1tHf1k7aEj/2
uzcQjDL1KIF2PKmmZWsY+DEOSyRfy9BDrKN5k+V5gukJBH4LxiUFXZsePaeE+EaT+AIq/Y41naBT
YEpLMSYSz/eRT4ssx8Y7jmYchODPSwtklU99O+NeAqlJTMMgGhPZN72S/8gVBHiS1Qp3MIo8l3eA
d0qoxWfA4JoUsv5xxIL5V/OkiISGR4DmRSJ7wG/3EV/bTpmXn28UIwZawTA1eW9CNYddZez+t+D2
hXAmpR9RgUi1tzbQwioc3cPLY3R+9o4+slduhU6Z7KpIInLyI9zikHZ3AamBlW+27LY1XvdSmFlh
NAXTlyy5s7Zj1vvUMYFNVB86HBRtVGvz9tCfj//nEgttP3BzVLD42O5KPsxPV43g3pC4hvlyyWcH
HHcMsjYgZWw6/KIGEyapH5WjfK0MAlMiSiYtaACWp+Y/LU8mvae9M1XjLX5Y9l/YKZ6gpXalE1D4
q0VJMVF+Sti/JMHLWnzta46G+UzV50FK6CuJGDmLWC9gHbJZ4yNUYyRSeNkkw6zkTg0d6OTKxbZe
L0fdaPMHi4bsQDwWVSabwcOCmoR+5C0tGm2g1JL02g7+MJJY6GjRDIZVuXYU41xxAH7iIGT9qJSB
+BbW3AmQeBrDVUFVHwvVyNuLM6QIxLeZxk5kHIE00OURWIWlFtbyZV9rJMNI0ta1s94+9FgXApef
Ev6tZICoAzPb83/b9yWRjbyZeYXpo9Ih0kyzG2Jgkh2h7XqC6oQP6j9UeZsqM99lt0EWgcjlWEfm
+Rod8iUDk6xYD8r65X8LoYMZDYqEcTxIhEjMt3JgFEDjK80lq9KnVSsekcerob1rcx0kLyjjAk80
bWRQH6iUd5qTbwfSdxYy4Dd9B0pVh+wXBHk2daAd7xFzBjED6aQ7kBJLGzHcOY7q3vnhSiQziv4M
wZHL8DQ5sHILYRPqryQVkqfVGSXRgL3k0fKcmHllt4Lt5S8CT+aKF88zhtA+Ion26ooBF5TGq598
BLJgxo+TVks3xptH//KuolAv8tNQcBckPXx3U9eBcQ8Pztoc5E1wqgGT2FNNPSBObprbFwMWX6O5
rbdQYX0MXPZl0IT7aTOvxeHFDlZvnokmj1fbtf9Kg4d2XNMN8O4iJrU4PtifiM4o+Hxmq1WefzvK
3gpj9Atbp5dJVRFcChByr3tkUfzpvjP1x/sc+1lae1Drf1bmwPmbYEclaJW2fYKeR+Jlaw8zOhxC
mJyjq0konafZBwh3b46ZYTXl4+GkIH6AcdZnP9JBbjBN4IKm2PnxBUTPlkyAcC3xP0m72jEtaHxG
HorfgOKrmxhv6kaBBm7qBmgoymbAtaxZciZxNQvoZdpLUfvhK3CMElPx7/ZlzzeGKDL+cGLeDbQo
N+j6GE1GQD/XIpiB9pFSeCDt9U4HFlqMWUqHsbOy8mWd3X5Tfzs/t9Mr0xly+RePHUgoAZWLdhHr
ll3nib9f3sGlwEO5oUiJYUKuoAgwpbUIMxToKzn1iyFOPP66ddqGU8BCTzg59JKMz+1RWTAL75sY
zJJEq9UIcgyezJFZ6PLi65n/dW85Hm9mP6IAzn0J5jUOgge6CYqs3H/jtDi9KollrXfP5xALOkpT
NIcR6zbmVZpSFrjo/uuLdmSQTsiQtJ65N3SMixEn5xQO5u+QRPmF9iTFs5bdVlMrhIYywgD/II5A
VFeWo6aSlnh/27tLLuuqikI/4x8RMbDF4GHUio2GzAX3bs09GRHA8kkoUe5NCZyknMpRKag9vKmc
uXXHruQpr+RCumLocMfTRgXmBMDjXLUfbOf7mdjJjRoIw19x3TNsEABURB/3iIScwSm1v8RRriyB
kvDU3mkrPVpL+NlsXXsAz8cMV1sn8nIWND2OiqH0MUzqk0gf5wtxYkXBBXINSUGDtxK07CIrfL9/
tjIdR1HKcvIhKAWrp6o0MpAAmOUhBOg1EIABIq/ddtywtvCFIekb016zJvF93pEY355CwYNoivpM
TQeXpJD0gjTVcLa8EVJDu9kIt39RucNKJTUg0y6PB6gZNxD3HDHvpWMMcJjdawXtFryewQXgw9WW
sPahJIVYRkkC+QeUNEzsl9nRTypSfJ9eeppAP70gzkQAwYKz9df3PGsZLA0sU3GFsdwHa6x6vIlC
8VcbAPOMbHdttJdM/g2ex05/MZEqVV0PI2EyQX8uZ/XECrSEdWIRUqKAb6wfAq3Mo+PUO48LDe9l
D3OKb7d/O93vqwrP/jzoAhRyWMg+ddkwGbzlU016Df+ISwCobuGYaBYDdV0aqfXSbrezSgIA2eYm
Wdrgl0XQkZxA0vQzUApwNI4VkJScYAsXHYk0Xb+UXuEovs8EJQstZvY24iEf9iZEGlZpVPpYGGHH
OTfHDc4ihIpB/+BT7ms5jFE4N6pORQn+fDd5u8mnHWCevOArgR8eU/214rTxcY4vc8QBjsFr/weJ
t5S2LHGKxRqweSatSwxAd4EuigjYHFiViH0Iq3nxLux/xskr6+WVXG4cIOwNbvl50ETpiSbwrYJr
VrWcQyw5oXA0Nl1X0YG6U0XtZZJ7iwPBiRgHHLnVuMNeMSLQF5apK3RqfIlDPf0smf9Y1PZI25NY
k3fKdXLcLDWHfIj9P134+AIoCxk2xUhtd3WLUuwKASXwFD2wTsg7VfrJX3ya0Pb1ULP39rRgpzfI
Ae03/rZLDbJwfFwn6gojH+D0umaRo3lNEmdlPTJGNQ9k8lkTyw4yoMDotCikLwiX95T0FPSKEhNf
aY/pJFtnk5dOISo1qSui+KBpRfVD3wfTMoktru+s9U4uj3oTlcPFmNgj6C80thPV1voHpKX24wiJ
nPlyyFrbHYhIDNyLw6s6Ct699v1V8KTgrI7utol3k90LiKdm1hlvCLjimPhQiguX+wsarWmHbI+D
U2z2LyyMOkkYwNvE+VRTU4eplquuROaPwxJKQa9myWNiQKq94MZWqdsb9Mq0fVGF9R70Z9Ispq6s
H9LxpE2r2FhH5yPkQ6HyBuihIoHWT30aQdQpOPG6xC7JLvuRzLnSXlEc6hX3D+pKqYlP/telcQgp
7mchlkn5YeC1See8z4vXpvIqKgIaWxz6fnWwP21ZLcyOxAqPN8kOVcAHHj919Reh6wIXrJ10dwSp
1EEGaGxtAAZsXqTjLwYgfqH7psXiU+063mPoqT0DJaZkhPhnJszv9j4XT1m9cidM3YFcdl+WEHWb
9+OVXiyFxc9j524ZD2TQmHuJXhxIkviPvurlgf63HJbWOqzrnbAuCQs449NnedxmqsrNVvcBbvh7
XLWKOkxYSGjFth6wRJDuXyOu/LkzyKBO6seqLgFCq6Vk+xFH2DBWOQEXB9qAVz3DMmur2Bd1Wsdh
vT94O0tlzmh3NM9wLj4i9Ef0uZbZkB1XbTPkPLSAZltETeLBGjiLz85eAfjIuvHMoRbZYw3inJMh
dR8R5fqg2ZJQ1lTl40439y9hQt1CwN/k5e9sbLSC6aELzLK/+N9E/VSAQPdxiBa2FiHkA2KmFhAA
3/KHQvtuB59LYlCUoVD9z57IZXS8yYtChJzz4hF8Om09zQlzPFKE/GKctC7nUyaVzVDTOuvdpNit
UtQj62/R+jg6cqbqWvzt1TexHNA4Gud6/3I0v0+rRtCQF3IvPfAlSRBHt6KDmHs4oFpvJuehyFCI
dx1NqeKKeC6aMoJhzsihN5ucrf75bbT213MgucG2/syjV/vZ75dMT4gNLN0iNJvrx++a9ULAoJZo
cpRe1WTe+xdwLNzTmeUeA93mTM4f3iHEYww3nlO9iT5G0HFkC0TFejwYQNAFxXb44WbCOetT+Ug9
MDZIpa9aAtDi2vprPhlm7N+OAyLhGYlBEJhhykCSLc8GNIBrENfX87wrUQyiDDBKmR0fLQZVt0iX
f97ItQSelZVlLG7ynkjc3tsYK8m2RLQ6DYyVZQ2LOL5wMuw78XMtVUe/bdR77mdE99jKpMPWDQ2x
JIZMXrsHorXD0+CebcjP5LUA9RLzeU/1SQCp4DEqYZOmCc/SAMfht3pZpqNffy2Z0s1d+SRhmzmH
cMRJGhDuMuX8vfjVbY2SzsMCEyYgVUnwf0fwJiqPp43v8MfmhNLMsCvENs9EgfWQhDLfTXmN+k8N
6I696vFGh9snbjF6aRWqXLFEzlArdidVD6oF4Aoc67wlmnr6u5PS5gLwcb7a6PiAV6Ir5YQEgj/+
g3Mt0en8TBzyF1/UnrYjplrgP3zOU84izz49B/iYOKXn1fT2mZbn3nMH5JsF7pYG2S+7gudbYolg
2+8Mp+tlev0CGLtOCRaITu/IoiNP/pyBLeinbCOJQOC769aQywPmDxtWHJeFm0UBOlNCT9IWZHZi
jnwfmkpvpnFuuEQZdwRLJ01R2TcgrG5XxympiML87Zc09ThDaLhRb3T8jw/8+QlUCAhq5x/+YBnD
+wT6BXxEwUneInCsEv9hwaN5iTC1RmJ2wU7C752jK9uo7J5ujlifn8tCWgackxcwBvZF03VqqipT
3dOL39A6wCFlxB0yK8hpEV1fgfWu4wPNEhFZzx/r87Dx4qLAnvRXJ/FWAbLT5RlMhKx86od30Et2
mr6ncwjtepDjhEXftOm8+4SM8Ltfkyzvcc8rdL5ANYa6kF7RRQsPN5gHKwqfQnEdZK/AG+B4/25n
qgT9DiwO3phZ1KEISfZiVoOQR5yMfk17KOa1AyUVnTDZRZlUzO0IV4UWJypwwoI7otWis6ckAPBU
Nzwa5C2xMFPET5OtXanxGW8jG2+Tw7YcIqrhnBmh5blMF5ZlWLNUqVOjcmwkJW1IJJhvetJcKsni
uHsDswm9arB+y2RAbWY7xfQjPZM3X0MCA9oBNFIHyxHGjGgoyCX8SGq3JJoJWkEWXOmRf0VbCx2f
yPFjpxV4W36kwPltcQvRpsdB0EVSSR1mgKP9B6jNDF1f1yiFemuKRpDwTuhlRmyjKM7m5lh/0G4w
8cls6ME1gKEeR/8Dpx1JuVYgdG2Z/TEL8ZLo90GoOVvno+JEq6a05ghU/4FIzHC9hQt881QcNBxs
ckjqtPAhtfpNdFEIN8q46Kbz23gAOYlmjhWUK2MV0sWMYWlys13vxYtr1Yy1mAjX+08qGHrkv8f1
SDC7d3GH2fba61PWEBlY+LHOQ0mwqXPwVceErdKclMGpu+3fWCccGwc5TUYAZfLAyBNT77PasWBN
B3X4DHZf+be0Q75fZgFuhL9m37kZmnaLoDe+3bSL8la9uHmoSfGvCQI/xk0+8zgET7seX80DMKgf
6lXIvmjd1Xk/nTkfNi+9VchfDuuYLmwLNWE9oDVFOdqcXbdiv3CG4Jdp2yFfaFuL7BNuAgIakOJq
EhT4r0rkMPG3v1xjyAY12XPGe8O8KxO8FPBJfIQu6cR612R4iUyAEYBJCQ25b3cWv57enJYjf/xk
XhhkZZZZTI/N8z1N7qIeg4kuSGdWzcTpm0qaG9RL+Jn0nJFHQri4Qs38mvvT0YUMwQo6SScf8nrM
Lpf1WgFHE6ktU2JCP96MuNpR8iz6SWeQ4BiQ3w5AzccYAoYTb05p1NtnAP9VBMdEwJXObsfoaztT
0MxfSXdQsfmdBBANjJNuNO67k/hbk3bPLbRvggB62ZKRdamiBv+uaQhPeFhAGo6++ocY54HJd1Ek
YAapRTx16MZvhInF+2xLL2/bS5359HmdforqsIanhI/h4ZyZjiqSDLhuDkJ7jHcQapWS9RHQArpK
MK+6Sv6CJz8+kE5CzHHc0aq34MqcsHFhzmaIVow9P+T65/DCUqhLByDvw2c4mGqjC0pUXdmYWugk
BeYb0jed2dNjBN/6HRWzWr+LwIjMjN701+eKJ3wTzrJV8GrLMZblMdeeqZfcOsKhO7TyYRrEfvQW
jk9QKj4IMDpjcED3pxN4z7kWW51MYIjgU1uVct2EikweVzAadOhqvQEjjom2geLQZQ7NgJL/Mcq1
w1JomVwdqM41pxUeV6tQQetklurSxhrWH8odAlI9b52eMI2tCNkQYDCtpzgeJQRgG70LuHXlLvI7
z7ntTkHWC2Q+oVtHGtr4OaJTTSw2Jel/fgggFskYEzHvpFNrAmOMx1UlgWj9XBvFCzUx716bngid
bDn/upgey/1oWgPvH4OgG0Pxt2IMihPKsJjpWBudKKQApZMtEOZfLOC9j6FibB0PCjuSMHri+bBT
2po6A1tave7oMmXV4xWrRxCWNEdIU0fwPzGrONVulo5Zg2PXSGIk8QYDwAdJwcGJelEJDu58tM+5
gPz17gaubHgdNSuANLSO+05aFHmqukgCYyTYyC8qVnMWLzQllNUu//WX/9wz3ImJg94+cxsBVfol
qoBxlnYD7Qht5Wao9EVxflWqR5h3LR/FOdNU1+DKODvVHObTt2n2ljxNE9P0KlXHUL6+ud3ohNPj
YaF1eQYDjHxRaPFec65lnwh/2uvGRXXIc8HauOeMx4G6IKo4ww/KTByXoThzZnRwPOiV6FO8imWG
NqTYVP0iJ6bWpAEfEkvoVqsUGgg/2A3pUNknfHI12BVmg4PqFoEhTXnDUEUPQ+o7dIrN1aisUuCg
fhv3+DzaOp+5eKifQI0HFiMbbjFoxcuu5Y5JZxtVlz8ytAXi6ao0WfmfQvIgo7STiqRWRIWcK1Bv
7Rrxbm3l6D/OvzJVerdwAGLfJGSgOA6uUFhYG/+YxTatjar/bzGbvzla7Vmix1xZa4MuNOCxHPlh
DcyDgRwIozC+yXr5nJuccZDrI2a4MbsfW75XNLSSMFF5UXHJ71ivCzw40HSlqw/MRE4P74F506hi
1QY6S5/d/oWpY25qHFcfZaTiSbK1zY1KpAdAzAjQ3f1BRmThFrBCAmcvHnJx4uuU2xkNRsIdYt9+
Ehd9VCmvZLpd4Py6OF981+EGQQAzO5j7P7tLhP36Jef7u5xGF8KEUQmtvRKKWH1UDFhCBFvA+2zp
CleRHo3QjnahZv+7wRElBTrA30+ufUFQQ+Ofwr7hWLvdOUOiAULeagx+/n65YKVoSe/PVTDcidgR
uKHjOh5t+ZP7BMfTwvDFTy6RQY7XvwqskmbV13dHr0CMAQ+HVWmiVaNZEmp8dH+mwl2ro/vrUM2H
rlldPTTJz5TN1qc847DzMN8bv3k1cbEUIQiL3lmo5/3VGNDqVRouCjySII4eQRdgU26o6SjEuW9d
DT/suvQZ9oCSJ66lpDjo2SbcZ3s4wt456DDYw5m8ZMYmG0H9VirZaNjfawVBPNKjCbwE5VOc+zyy
trcWicsoLwj7Kzk/msDAbCd3ne8fJsnw0Qo3JMUJtMOPIliuoefxGZRGFgIldQuw3X1qYlBE/AxT
7NwWl+BwncSYVRWke8XF/9F9JJvLb8e0Yyt+l0jJu0vqV6uaeOVHR7QglIr47+mHIVpYJSOolgGT
7l0jJHKf+l0ihmTXTJAEytem/HkpvofqB+IEoIwoeWvegcyJfFi5FVyO/gkKxcPKxgVoFVvsmv70
rlH/52kQbdfbzZMDXICBJw/B+pE3T/wY5HhbPY1AQMK5w7kdAsM47XcbqvOXZROFbbU5Ur+uVkxu
JeGYWkO0pQP0bC09qoH1PkA3RLrC7hjJzzPf++WB08JHkRfangYEdVo333HNUPlTgyi7vVsAc4ii
iVcZ8lr+89vxiPaY4WSYdo588Z2asB7x91H9qpycVzdfIWeLOlUtejqbLPiMFPJy+Tjfl+xrnROY
YRQOiHYKAS2jE2GNlySkxMIhSIkusjjFGq3Xj4GYg8DnF2nXYvMsVn56Pkr7eqNAKt/ZFzysHPv7
JsrWFMkyLiWekUExbBZ8C6TPZL2vdaHnmQM+bqlFdhIjqkqapZ1GdJzWVqeqk/D9rSKqoe2zgXTH
ajfUo4Z/Y4aDqnTBlMScwqhSoYiznRlwGSXnT3Rjw3OPhfYzDyFBszMZk1Nx/zHphjvh7ZaTgx4v
4yO43NpjaXEq79AkM83+cv56cefmESKzlUiundKZrrQc/oiWjIWrA8QLKNtyRbfMPVZGtH20d89Z
gdV4Wn8lwnOVEFOJ0VPVWmuZR9bniBM+ae4GDAQSNL3W/eq9f91CW/5jnCkBCFagCM6n54emT/p3
dmXUgek7/iFu5IcUzqd211wQHjeB5sDhqQ9RPsb4RjA26UuE0lYZepGCNF8zWOVEAXViZNwqO7tx
ekgzAzsVF7uT0e9JfRallfODlxgjv/YWcsxf/j5JvMgSHFxC6gqiTWb4zw+L9aTpH9a4ONhsc+uR
XyEbttTwru7oX5ypecuXgFtF1oe1/W+jBNUPgs9CydMdHDcSmMNZL2JTU5JBQPTJuAlGzIFE9lrF
s7BH8zL1AZzTFR95SgtUZXGMFkDXV04HvGsH2JdkoyFxNr0hSwNjpfst/sMPmiiN6EQkL+VcY9eu
hpuVMeFKKxuaas9i9PV/isUzJYmtr/lSqdiNjo9go/eRivKNjUPQ2oPIBQ1RQ85ZEg8NGiiyma2W
7lUC1NemrMgC4cczjAINOOoKyAfGk35BIe8/xN1UXqqzNgJNHxXxdKVpDLUbyYtnlpO/jKprwQY6
Cbz6NqNTI7O+Wr5TUsHxrwGr+8rWaE5uqtZkjOHmoBZAsl6xxaCCR4AGQPmrsa7U4GKnfmBb7VOj
XNF6w84eBK5UXaq5T1wuMshw6PmeWMxVdhrmIYQ9pknd0uJOX6b030jx2FWtfmQr5WbygJM/z8rb
qGqkySA1k3ZcNbFQS9lQsGwD6m7x37G+EUhEOTg8sQme0t/vG1gEW7TCHiHxG1G4VN1tjnYH+N1u
ATCTIUJHVHrzS1P8fh6ZI3b5e86PQLLhQs2ctkL/k5ohXz9ngj1FI0cOCVL5nORJUWgzUwZqmMpP
gNCKMt10atNRtDACc7ZG3JsMXyrv43Abhf0vJyQa1GycFPTJMtYYe69SjZnLSDKdt09S7NMq4uCg
f3f9wbKJ7f3814JtjIO0nlC9TjKsgaGrb5Mdmwu0QJ1G5CwMyF0mPa543S2g+aMTctj8siIBmYdd
u/eCKWQrx2BvIhT/9KRGT3egVbyb0bpRp4xsJCozB//GOUFgIXsOum3BxZAtLZvu6Spoqg3Y0XGM
2edcDfyKSTc9Dl3FP0B7tjpA+KrZAIAiUMIBTKS9dlXEBi6pzLI1URmw2GY5C0HUIdeHJ/gCBpIQ
m+aj1hslNAxHd5blK2bpiqLswwvfqP4q2V6py3jT+ivQ0NpxX3Nqmd+k3k8t0oIstb40U7eUAz2t
WZdyZzKNb1hkpWrKQo/sfD9IKyZTYlXLpQS66FlVLGS+EZPzp67Z/C9jf4pXkTaynr5y914B0ukX
a8KIaHaLhv7xorF5Ah1Yl1PHL8EVpOuBLuMi/iz4gRbt8i6099wKfSb534ZxUpLntDzCwcLT54Lj
6XWvuYbjtKe1s4gKtiMNqvwhskhq6ybLZT/8Mym2shypXcXr629JAW6/sAUvOhAlZ0KZWNAZUVlG
hbGZC6hKG1z4bCki8p7O0eLGmEH0mAghRJG1A+1bAp6368X1otGqMiD8al38CW5FHy9E/gt4Mz7V
S+hv7EprLI/Ip59kMuAKbkv1wvVg1gDW6p7KqKmJtVRQQqE3iT0FGDet8gyj60okY7g6YI19s7y5
E1FdvwKJIGskliY20zzll9VNcsVHhvSU4gc0OZykOepQPKYl983nGDeRwstvS+j18tkE1ORQnM6j
On6JqtHBKPbtl61S7ts6p3OJtZZz+SV2yliNVZelSARSfoHoIh5oOxU8fk/t619axzD/Qa3U1DnG
7zyQOcxgNNkJ9PtgiiZejWq/WCaBR9Ov9X+EjRl5OjRnuy4nQslVgm5N//m3oPj5EHJt6b0WsF7O
CdMrpzI1NZMPMJdipELrtQsVRQyP47zSWxsJb7hkZuvV4To2Fv6BTbi2xQ77LNZgyJ+UzDb8Ec2s
DKFRbskMzwaYLWufZzaGCjC6yeXTf3nW1kX+rTHiBjPZ80IZNuXBw8Hz+SW3IRwuVjkbIgua7acX
YJ0GJY0KsEY8WDeEd2J+cObORn3Y6kDoWlO3SWk/EXrKyLd6QGPSZrIYLlWsOR8IxnPsq1vgEoGJ
Eg2AaqX3LLDv4yQ52xi2Zy2+AFZj/tAaZWZVjNLulPoVHPG5eKiSjflSQU+LtVz6F0bCiQQHhEKf
u1V3iFlVtAKN6Uyp832N/1A8S9uaGyl/bdkdPHfBwEaNqzTw/3dzaCcM5p3wPk31hBkksRhEJUIx
SW/ZFVe/alr7uxLR2gmqNr/OJjHLoO30NVe+TIkxi0W6q2A2itsCWveW6CkXmO9s8/W2bmwhovHG
ZuSVyhaOp+g4lHGaIbJTOC9G8eDMC/hKln9KeDw8pz6E6QLtIHCtRBWOBe8zq5rNawDjwkXWyTMb
VJnFnfZL3CF8Sx+XIEeYsuzAUX/ncrHNDQBowcMNULSVr7zLc2W00RQdi2RglxXXLBzS+hIQEO+n
DRzA6aBjcxx0ZS12uA7qB7Uhi5u6LzYIXLGWXc6dNg+rggq17kds8zlreAd2PZD6uRAs0kMfSW6B
Zf6xk1IhI+dubCNq3pkKo3FJkzi0pZqDcL4ACjM6XgxoMhBC5JivdXI/ghWs5XmDZwbilxyD7oog
2q7iwaIG1be2g4xUoqvl8nPnLq1800EbSbSCilVKr3ADtAtvVRTKla2bNSNacUStLt5h2jPkDd5y
wsVUw8QjdIJxF4PxGB0k0dngppArke3RjM2Dh/W0wLFsPqzvoExGb6NNl4WlYkVnFhJvqr1wb83I
v5yDfCYy4RYyIAXDFMEYSJej8NebrNcBZdl3/ok7qEMomIPgnTLFYNGYIvFesoqFi0eKZ75DPHf4
r8Po1ZFz7Ag/JieamhiXKx4Uqvb9mGRzv+ohc72dK/3KUzUBkNYhQTCTLP9f313GlLHaLHz1N7WY
U1cc+gFHet8NH/+uGI1bTf+rLuJ/bOBvmCpZg1CAAXBt3uZXHGwX/Lo5MkbhIWqZMDCJBbLzpqxz
hxVCSca1gCISXVkSDnupOpKAVYnxQqysA9RM9ovbMhpYZmBapATbKoFQ0YioPE0+JX2zMLHud5fh
FutsMOggtWefs+fibsAOWvgSWJdamOPKf8LOkzjugjuGdMTVoV+HX05JzbxZ3VPowDssEgjn8liD
eUxSmhwe726A8CBUeLnAJzw2l6CgTFRKH740Y0Dx9eIVLMS2yWgP2aRSg+JNHe9uV2LWGduTLXre
QZqpy0obc6xuJ7QITP61mCv8MQTZ4fXwamREPkkjSIYNxemS0riVO/REB6zoUGlOFj9OT4dmja2n
bxQfzybHUyG6A1CGrEo8tqj10FebiK+FeHPiwMw9f87jeP8vJ4eBVurlO3/ALR0aq4tqdThw4DFS
c6m9LePHLSxcg9fuK/GJuzdoR5+hIGydqm2MwYXPfSQVbqsSPlP+xSOOLYIMZWXBtFEg0jGOvUln
IFu3AHP2k/YQpa/nCBr8+M24+DNCm6eucU+8M2WQXXkb5SWwNqFWsDtDxcjuLqJjYfHh2Bk3CNLj
xbCcA4VGMqs0nTwxjYMOU6EpOQR9tsxiUCIScdd/Dfd0XHvzx49XtvSKksCOEv6DTBl+m8CpH5U9
yfWG9N2T5DLBnn1BomM8DNfCF/4BRV4x1FvbujUhK2Vm5I77ky62vHNv/iXhXvKVWL9k/SkDTZWx
ZxJYk8NXG0gxCZe+CSvKtP2kpUpxzRaPBCO495Z59flVHvZV3xjlOjoNotWoRtZBH8Z7iFrqpOme
3/BEMfubynk8X8QUksbgZv2eKo2yVSMYSSmwxjhzA7G/nggetDRdnPn6WrPzhO6owpULpe0/1BAK
/bagTCy8GCLj2vqZ92RpMaXeTROVKeIhSuZ9sfKWjku6iLAnxA4BqjmV14P9BxSUCthdF8/aYPfz
AbVZSSjsdsOdF32ebIotlLngaC2H0DxLGigXB/4deI3zrC0FJXS+5tkL0Xz2RVZ/IhAjqpVWjpNw
WgKegLbfz57JY7ulWWdZhUru8qHon5Ds8DHSvBVED2MC/axsvoZHcAoiC6dAf/xphDjl0IiBIUkU
lz2Wuc//8ueFWP95b04279kx903lxsB1bgOIWWKkRdB78ID3qIZe/6gyZEIg3PaqxeYMgORD6S69
M2hUKS6Pj0Yh7R3XnF0DDjmW1ddK9PtvPFl6Xm8518tIg1LQuMtq7ZlEn5UFEAOFW8jiKpAmh82+
eV2AqvJ8XDxFstxRlAhoOJbm9EBMhWOniLIZD5o9R8VDPkbcZKb93vRHWs5sAJuHCEWl87CoGDBd
NCJqJGVJ8as95OiX17C9URTETQPg9t3Lb5D99poqemZgMY7lNT++B17hSPStJJKDEmOqLFTOt3mR
PgjgoWl/teGlL2yshDcexQTMyW1fhI9kxnibKE9ycQkyvuOgCM2HWZJJASgI56Up4Jlm8d9GCvbb
LAEGT4MfmoCt5ISkMYc58XGqoOYxyiKCG4LdVyVM6Ql4ElFekzZIqOZI4dowgh0K65OGkswabSOl
/3AafZx1RakkNdyalMX6Md9WECAt7Cl06E4BjemkaoDhfTlWKJC6fyoDkuGKANOs2gLFHfD0HORq
JLRqRFrDr4d/5exg6DUKa2Kt2BiEjGtSrlL3gvRGj18fCA48Wsuv+II+ZRzG0UBTI0zZqYYwce/M
/E/AbZkyNcpVTISvOY6XaYCaQq6djxQpxiLeJdyvlc+JtAgu6vi9CIiY2NoDe6crQPrFOR80DuKS
nxGeDeiOogh+A0nUYLq7ryxo3ciPaPWu/MasKUFP1OpBFOay7alx9/vEjruxvR6Z6jU1WDAcB3T8
cfz+nl5kYt+aaqe+WiN33cX0CKzW24KHGafaqT3pS3TncQwHsw/N8dJAxad5B092Eca3OFOX6ocY
3krHRzJq6JDGvAHpvQYSmqatF2SUM0JAKQ15deGQ5SFYYhXugPmLWpEnslysvPFDmTgoqrpM/FDO
3NDivozspzJFvdPpKA2N5i7mDa1pKZhM+KIOdRTMPckr36O+ExjSwY9Y8CrdSojPmaFa4nwESlIU
CnV8VMy7QpjdEJnD77QskiIqJ8jIpx2Uv1IPWLjBNoklC0Fbc7fspyqzc/s0Xe5397804ykr6iuc
gHdEGjO2A1ElpQOHgvdiV+G7y47xIDcCiPKMtMm5HeIgUpCYKPqKb5AjyyYFhtbauK9Nqanzpj8D
4CPNvW3xrieYEO/aFWrwsd5Op+VDlDQVIVgGRhcS9ikKUTIpfvt/B+vISz/++CSNf3WtoMGsaIwb
qjTf7Vx4MuvyQccvTRM0AAs3zxKKkKKpT5YVVOhomdhEKUlaf2pbeXfIst/g8SFCfp/6+8h3JKhS
zk0q5qm6hVAm+DO3FTRpa4/7ZbL0Z6bYpbVc+tniT3Q7bgvk14QtTnQ8ghDz5M/lrAxNmGNHrF0F
lJzjul4Scfqc/B/3Vx8V4GHjuyGI9g69iUiO4DQaAO7+Pp7tpuM3FGyarUTPL1nUaCivR1fPc4ss
+F9RuQZDhlBRwheIi7sw3ZosByOYleuuPWMPWD7lfJLcPhagdQe7NVS+XhxDOnaS1RTTLGGZwh2t
rxUBcfdcpA+G7LVFlhfbClfRdCrLXJ1ovWbTmakGQmD6eNxgO4xlutW5iREt/sK2lTMTS9ZQnedu
pP3IEImDEQRHb7HnnyuGnw9xDxEBY4EKvxh94DdA9BdH6g7ZiOuGQWCpC23BoveCRu0IavJjd7FK
AWNVzWgz851mNldhlCb5/UD0t5qk2LbF5XAp4szJfOsDlgrWINNBbWdB3NJsdYNZS+yNjb/aLuRr
42VHRBmRRZrwY/Ld8MlZtO8NNt1r6q4fWkNh9VSjKYKgqcLQ1aPJb3Cchxr+8Dh2PREKv4bMO/vs
Fya1dWA+bG3skI3j8AewxN5V/WXM2SYHzi7WQDwT0gyVNWtGeZrQfeW1fiux+fRUfYQicwgYGxn7
IA08Z8yH2vlTwJ/IqTTmYkL0zPJoXQ2I9BMtqkdA+Aw4xEXB7B3jheMJ+l+Hdr0pktANukDP2BC5
bX004thhaOFDTX9sIgt1wIJ7xNnj6x3sV27Hl1Xz0+JhIXLHEfiUaWDjaKJ9qpEoLLK24fTyxVmU
L3FOqCMn4dbmm7hxJ5T+ItB+2EPtOD2rMV2lep95XXAh+l3OfJWVFcYmV4Llg1uDzdQ1G6yvixXW
T3o9cpp0mDFAGQ2GM9uxs82jrkLpcBD9pwxb9C+wvWtQGox4sa2Zwtj6xC9J8r+0M9aalnQggOky
nhGaJRfLzZrHHGY0E06b1D69kFrqQ/q8ppG86AHlViv6QrNFwrxyyLxO0bPBptt81YAn5rFcuruB
CVaX0AhR8uanrvWnO2AF6kgzw9Cb+WSOoXmGQopJu2gl5DGVSAgTgDNrLw/PiJRULm00/A6l91m5
Sx9UzPFzk9zUafKOY3fIFjE54oywPoz3VZpnf94kBQ5wQ4ebGwyRGfBj9ckJ52A98jjdOIjC/g5J
LpqPR8U3hGzhtfXQrGdHcaMW098O7G9vaA1R6vOKwUUiQOTV1YZIV3zPZ8oMh04qZh8W7njcC1BV
FLgI2HJGhacTHpN0yfeFVDDosxyZiXaf5dXxs5E2ktLGmR2fj7iIBF84oJNOEzCvqwGpZSsg23eJ
Bk7SSks5me5qxDzF0V6aMq1BmYzvrWGywcHkyPGVO7mMfx7jLMCoHn2YpJY4oUBTHsZxETXwrEuE
Rhe9xemH9lvLpJ2/sfWAUhEPgX1ljdOuf7xEiXbfm9IjlbKa11pXGlwsRNddybUBaJZeozhHJqev
2j07cW7g0UewPEfRr4NtbkgkrNybxjLk75EacAwmrggKlD0qvRa5F8QNbgZlxg+xmdI2oKgWBbiX
UPKUXFLxRe/kUN4RqiiHufAMZf9n255HBDbLGM12Id2WDi1ji3pLcd5vYalDCqcBU7bKKgByt/8V
Njkd+NYbbAU/kh14sm/ZXI5DIwnUlJRHhOkp7pffZ/JhTt7qP66NWe4jj3hz6e19vzdynj/rfhwi
7sefACIqoUz91x2n6w/I4h86o4Y3vgxiab3jVjl7jJmbFCwFLq6CYMfx7LQRO1h4U9IqyVX4qz3d
8iegTj41Ou+R6Rn8nqT1Z6wmanR3jHJae3YwT/A5qOGknNWSxSrHkQmGdSllPNJow4SPuK1lTynW
TKPw7weD3KxV1tHBc0hHqwauS5jGvvTx7x41vJEsnfTAYuecZR4lmjsQUcH8YvKzZ+1f37DesrSF
y/Egjfl+9eyvgIaDsxNrvMTxUZol0PynoJNEVtA//u/ouEpzCJqgLsjW0dtpZPhn2e7hzwg+//3J
yfaED4/SQEznY4XX1HZQuLM+yGZ+jcZqLINCUgg7LFS6lqU6ZSgcg/C+udye/n7ZA0tx4gJNURgN
ODXL7zaGwPp9YK/2e6m4n7w+ufAJZjrYW+pcx69DH221Y1Hg/DSuZVK3550yIuNkutIxmSDKgji8
1FPybk5T4ax3bQ2ZBM0JGf2osq4axFVRJYDSkr+X+Ag/oMyXkovkq7O92AWl7K6lIfumtMky47Ip
ihvtjh2rjCi2PDiuNTA76cXqJzTU+uInAHvS6UCWNNeLuz93uM+g9RHqKEKdZymOB8WJ6ovrI/aX
PndHeyPwvnDRPrftGhEw0RYLUx4OhpJZxTdTErDOEi31lPtiVAdxuFK711tbIahh44uZRBQ3xmMf
pobGVHZBQgoab3ssH6mN0uKLS3qosuOYTtE/eFpNqf5zAh0gQ2Yk+XDJEBBeIrc0EhJ0yK2dN6Bm
K0lOsFeenZl388oAaJQZRnoMMsiq6rScbAGMkLGFq4nG9GrvPEdlJqzR/DS2qEG8Lb11daEIvFA4
7tLPhe33fxgmk71SMKNb6wsLQuOIaxXEFi6j/vEOPcVgtv8Ub4r1vzC1fFfsuV92G8BDkEDAb5xu
qmBu+JNOnvSMcP/qOfPZOfA1AC7rJ1QCOH35PLO0E1hpHeW+tAPciBN+qY2Vw+9nt9MS+gYdPOmP
8sjNkirjEtydvC5+rZKeRhu3Sy3/uCX0341KWZHbW5Nd3MWc3S61oFLmrWpLwLQeQ86M6nL/fTcg
0nrp/3F5NGpQ7QgmLcd4ie5FSFQ6CB+DqH8mxMzRIry5l74XgiLggqKjc5OJpTtcHy0bYAuBMyQY
xXvOn7tpfa0xFEWWBrtnS1ME6hTm+GQ8cvORHbke36NaYzoD5vXrXjhlQW8/Os1GwwiTrtvndxO+
Kic58FVZ8/hERkHXUzKdnn7o0h6rNgbC9j35mWSipF/aaW1jF3a7EbX4lNxbMj2nH9OMDSYKtzod
c6nHRjYg6yEkke+Lmor58KspKMeXq964OIvtgkcWzDGlWLHObkhBUWpkS7rV0U/neGo1sSVG+s4b
WB3pZtyr/EzNfUE5QZVSAsHcOO0cCQnASeamvdf0jlpN3TkMmT1nir2wHY4BHz4mVW0JpUX3JHw7
qYFekaK0o/XcxH0Y+Ae2R+CYugqeAeZzNPSi72xGX8T8K/86qyvoJJtfEEgqZdU1R3qlKpHjfVYC
EKtxIN3ziJk+iXgnz13gBgx6B4EAlwEpOCQeKyrT7TjrwkLEyxNAqHocDIgFxVz7NOY6Rm6egK/R
Ypx6vBEtXxr6LDUzTqX1UVoMb/21k4GRIs5Wuf87NBu31b/oAlTgs51Wx+LywHftvIXshje6zj8w
93OYNrc6mJ2Zcxc/dsUEwZr62uVca+AdAN8w7Lo06IXpYnBtun3AA9m/yDmZV0KuVPnDqr3CN6YA
vml/gd4cH0cbD/4Mc5q1yD8O4vALPujTBs2MBoGsG593riXemPs35FTfI+abUwKLRbkEWyLx++LY
dLieH7MdWq3XjutoxpjHCe6fwt5XS1/fKtv874GjS1YRXgvA7PC8+6OE042Z8sSnD9Z4CB4NOPe/
U0ewjalqDjSej3v/BVdgBBSgd76/RmLADWT2sWTJq7henkFq6EIJqN+C5mlXUwfM0rYoI/mNa7tZ
XZouX2EUA8zctDA8z9mzczTE3+1WLSOsnbSebJ+m0c2X5qBxenFyiXUVH4SMcFc7Vu1Xjv++XxAG
b0MeFQ2olBYaN4E6hhnnS0uYu+mUWYutKXDVgsQYZGce4w7HMz8B4pl5ez05zWQOqHM4MRbrS0lm
XyPso/qz51wEMa1vqKo7jaPM6bMAlQiWXyjXS+OT5U4OSTMb9XBC96GRE2FtM6mVIm96w81dNk7G
mlEP0QqNqO29umi1YNq30IzmLibEprD1lqQnbmNCMRXXQGMbcUKc4BLQ7Rpto40G2O6zkU6TGRf1
kCy/f02Dvw45LDg34+jvPjc7FcC9c2HmyGuCHdAxtTJzoeaCH7tqF89Zet6uOJIUJt6GmQ4+3NOC
tvOaG/RKqMMtQ/DQiR6CIL6XBHSqBwwvUpHmeW+rxOU99YXWqjRBwbzQBFYaTkI9rK1FFoq/E5xI
pj7p0uympLGT4VrJjX/bUeh/gKtkipTohO54wwWWnvLUhPsCZmHnzVnQjTCM51m8UdiWAlotWmpY
h1t2AdHa2I/xk19jkhU7sfB6N9gHP/nUe41LlrxsKtLjx3kCElPyQ1lGY1EiYLRTHnjdrgoU+8VL
sm/T4KX/qOburflSHFQ2uwPORrg4G9UBVxB5V0rACPTj73sl4FhoFz9gmxSkrWQpP7tPl3Z6y0KS
DV8haFWrUk6YK3d7rlju+1Vv1cKLmhx46/BpXxCldHjMZ/ds8s9Q4ZVbSbL0Q3PrTrj1qlUgkP1U
8k0MpRKpIVDT2j84CeXxx1z2D5Cw3wsDvDGbzJ6FvRl1j5aapUVmsXd6B8VOlcc6PN76voeLOkih
mRNn1lXoKqZHRGWpm/8IFE6NMtRzLb4mxWYlunDSiuUdCqDOl0wNcPCfdnPMj//R5DQQZxcX5isO
qGC35N3tyHIgqZH4Ni29RpIN96NTSBSKKR9u/yg7PAMNxO36sLTrTGk7SscbifQGFJoqW+yMYJt+
fiVeH1NsheemEnZlkjqH9ttPJ4ffI8wisEzirPwzqKUIWEssIJw4FKJnPFFgSWrVJ0nxf1shlrMQ
Fm4V+CoalP/pxmmmKTdiALeozOT88kqNT+atwnEQDN72rWmV6FJLE/Ejc+jwOzr+BMHalHJMHsUV
MAHi1UvWkCZiYdMJMFpUbPuNWsoGfNEXIeyl7Tm9esCpejXdIQQ3mF3171/AkP1c74vXUoocWxw1
w70DZbmJuLegJpILSQlzroP1RT7qZKhlpVLWtxqNr48BU1b7Zy5lA6iNcm0rW3rx4/abGdx6+RnO
AwcDBXZb22jE34+t+cpjmgBj4h4SlW9hi+auK7nPu4qN2Tcuk+nErFCYy1GzBaBp8HgJctHF3hAE
tM8inAVnz71zYJd+QDbck1dnHizAD1XKbmfZ34m4E1TqCV5tORMrLKYhDFus1EuwvxL6RWaVhZIp
D8epadcCNuzYRZZj9wBS7U4Fp7h4B3hh1wCsICuTVXYU2Td8OR+AvHfVoqG/T+KR8ASRHeIQ/9oI
/eBzS6e1mp9+y75xEckbY8hLD50wfDY91UM+PEtsinfEfWppkyou1rsbI8slWaSQmQ0GpF2sHzjZ
PaRk70P6gvd+iIi3XyhJoy8TNYmiL0zTHVUF7lbtlBKULkqXh5arp5zcEbe3HFrZcSLGmLj2Gh+V
wqCGRRlfVu+nxKmAqdV+MCujZaj//m3GnhGzETWDn1PwC1B+J6dVMoKxYXkL/ZjLdq5XuhqQI+zt
tEAuMRpXlkEpnWaEpsz53ZaFBOw6MmOdbR+ss7HmZ35qSLtShrjC1xvRTgWZobkJW/VwY0HKb1E8
yJdKw80lozaayiHEeqdTRTUsnxVcWHexB5EzbTHqJlG+mqDX76w5u8t5g4bM9v2N43/pu5mJmihZ
Hemnle0wsgTPqIyKxky/tgp/CGEGkeWa+yXyrovERXtRFy5646KoWF9Tfl0MOSbmYoaafX+zEiq4
SiJiY4x4Sf5LUerXO85Gmolvny63EfkZ0W+CWfELYENemEgeeif78vRQsx4Ckq8osnB616Cho94v
JWlYSLkfZ9Lga8zGGDJ6/LxTyQtv7hazHSMzsQuUMvgRuOYWgRXSaABojWw8IvB5xZCTIIHZsoUy
qg3iXqHQk8uK5iOvl2FMOS7BNjGgPF9dVaPy+ehfE72X4RC4HSy6L6TesOLat1Hq9niHoAPPNM1h
Ga6reFmDPLwdSdQzL5SEXHD3EGR/UiHaF1uKArNSIudIjY6l/vNT3P13mbn4hqoh26DFUg77c8aT
9T9NG9Vajr/f4OlrQCbQ+lxb3KuSFPNVm6HSEkTSq60HuQTs0zBDDG4fimuCK5rQMsj9Cb7wPe9w
wvz80zAbyBW8zPJFeuYggsil/n9fB77Y5IiTm8AX1poopYB7aVUf5JGWptgx+k+1L/7RQ4EmRuZk
uFZK0N/yjXuuJr8JDf+1cVTuC6cbPGPeTyusS9cbrKuGeB4+mwsfrg2TNtyOrRpP8FmU6cPWokEO
V3eAcQq1Fl8I4lFtH8eY4pU4vXdwJazuaPCNrjwxW5+Osm0poMM0rBqCYvvCnZIhxTxJYkAQoVrr
LW7CyEWjSp/SSGbXuCxuHZ6Og3Qn1S46FrwOv/TLd7FYWy9oybX+IoXSdWhyb8T2E+PK/Eb+S31B
VBAsqhChr5hl55B+dSvbRJj8/IzZTJ8grWl+edINWB9UKy/JNavFfhYVo9RdC9Op1xoRjK4tTSaZ
jot+sjk2DHiVvArguoFx+s9fPktrN88vd8k7b5QTUZUoc5YHXHE/qWswIjifcm1912W/f2NgzmNh
Tiu6lebNzLtFjYLnQKkDH6uX9rqr+YMWKqQ+M6z/ht4HY7llZANqmhs17X0Gi+0bVYys161AY1Yc
Mv0aBZ9BEPtYdwv9ERbrkFlneu75CNdhaz8oBMCYySnrt62c/Bz3xdRtqh2180fLvOrl7HueGtig
5u0zGaZqUk4Y8FLFslsuMK1+43bAv1U9EuAqRfAIjMly1/+OHpIsgT9dE2oeDKPrlLM8/+52UIuP
64ZFSznFTSOEV9ut8Hx0j+a8D9AdBftUt/HjyoWunRrxQLb2wwJeL48b5abCpXXyR4X0OFJOKSf8
j8aT/jb656kxFhm/u0kNyXyr7WqMMpW4yvwbqg3PVQ3pDadesqk6/J0NGjuczi2gl6Cyn1byPACk
w152Lvm+ykoGPxAPXvE4e7ZUKcqpd/tGXFxUFWYfmknVHkbaODTf/FBjxWdoda757seJiB+Id69t
B16Htn+rFQgO0egJUHkLLijZjK73mgfsui+CxXpVzxKbCotWCfdK1hHoOw+kOvDBzo/RFei27eNV
+tOe6k55HApmwLxvVgXABuyR3gfdIrOU5+10xI6eqGNDd6gzKgzbgS3/uP4xNVlGk1cJqNQ1uf2S
3+vbohok6ITjPltzmpZ7lnozXlrglSg14+/0/iR7oWVZtkbANQVZc8hCu2jQnWkyfX7EsOtqpc4Y
sCjTNDMIYCrOE1nXbyxOKc8bmDKXZ6hMnRhKJmhOFMe37zwI560wT03Zxb7kQgAEM1M3hz98cASh
KH724CFdBoma4UZUqru+bWTls9ahYYNDSUxgwNS4ZGY1ooz3s0muZ3VNq33r24DU6wULWq0rwnbS
duLsrIw3tJwEKs04T0o1ClTAsL+idOwPFkQHpmV8HB43NGEyzWwWKP/UhmgyYVD6oSTIVYYf/Hom
XsiHXjX/uoO8pdraC0/8yGcM5N8qFis7m2w2gVxjYzxQDjw65pxQ2x35avMbqQcQ7fEj9QV8s2YF
8A3ulEEF3KI37bH82vMJzjEv7K+VxDiJefyo3YruUE2ks2XjCt7Mbd133cK31JK6uREGtvbD0SZV
9JToBh4nwO9ePZxQ+y4lRlfYg3K4qCbGmxhu4+rqFnUnjojnXTjz2cokr5b2wqozFgdEbZHhudo3
EotHdYFZOfkkK8z0SJ4UMwdu2erxtz6OPkYAeu4izllcYOlwA6B41ukAmqxZpr9CkfTGLdqBbMJu
n3AERH4V+059dgl3Yo2dk2tDCKU1kg1HqxvFqD96+OjBK9hSjv0++XhGTo3uG/7pw2SUxt8szy7M
RcIvYudqt84++El6zM+Cuwc8BXi4szAtx7fSOxuGzPDUI17Jq4KQNjXYB9n7uNhyK+HNv3kD3Bhk
A7AghA/GcoejYVN3SSvo8AYuTRNUmRLFrprWT2PxKZJ/o997WeubDv9KhzBw5QZSKSWlarJgdmP5
1llcSWyv02x7jVo+wi2uyjdlFj4cUBUqwQaf4+G6hNBRV26wvYvTkGlgZTQ7ZtlFKexng1nnERtm
Ifem2zcIwm0KxA1NAw7VEtk5zklVNHGS5mW/xwVCVKCs5zIx2Ik9JpfWq4eEJrBI7OHFfUihxMZj
coL4y74+zQrgyGb/mXmJWOeZ1vqTXJ3WZOEYZ3HNu++5VXqaPBcosiIawfcVejVZFoZRpC9Yk5v2
wXXuTvhB0sBo13OmGGSusDRUiTLYLvidnytG1v69a0oZIWK7bunhWpCBVeQGVj2jryZ+K/HUN1Zp
+D5EUyIlyrFyD7KPwMtY8ttErGAzYKKj6NmXpP+t1AGsxBL6pDF6J7+DyKoxyvDbh5NJQ++q8Jbr
DYAGrKbWcmd0ty1Kx4hqIhJ624IRywlLGjvlXhTN1tV1i/rznXZ+XCSqIbfpVNDwZYz90cbHlD4u
b6NoZDtiWLqwQc7PEyj4lhCdCTbf1j6HvpbqFTgofBSffbxZo07sYo3ZpCOrd9m4yf3C2IRB8dJ/
VodGyj2Qblk579Fr5nanvvCXcUMJIxkyO8fISv16uobBAOMXLsJg+Nor6MbXBwZUKsatZ3H1ngbM
XttcJJzcLGAU+TOZmPWazP9WExZxIs8j18JWQ/2byPaqbb15u/2oVO2ABgnvhvfk5PIo0ricf4Qb
0xjHuJ7lzQtStCh12zSeQHtqXvnkysaIgRzTOTIytysfTdWKa+eaFJdjEs9PIejtiZ34+PVyXDkG
PVW6rprQ3wVrFR/gQWjAqY0/46EpxKNB27qtUhwwfe6UFXRcIh9xVaRNGV4rKYHzCx85k031KDQI
ScQlhAKjZHRuUjEQlz6RRBoRSFfeDJSXzo0zh5+/OJfO6Ogkl3Gpe5IZdh8uE6wNHZONsOpZvgoI
GWBV4fgmY+uFcrR8xfiGMw6W3aEpoCdiC18vRyCw59CU/UHGbFe78rgk7BX7BjoDXQysHspsFqtW
XWql+RX3RsaLow4FnJX6QCtd8M89zr4UDUKjSvhNa0GHL/oqlHF0t7EZ1UPyLVTjuNny7Wm/a9dG
RjLRODkDo30A+ZhRsroTdbvwySHIFh1Ag7Es/RpJ4ddSWK2afubzXMaXHfOn8hxp5iMd+/Jq0eEd
3bD0CyY36d2Ia0Xd0FO4CBgw6lifdtjTK+hiCTn10TV+3cWfrGGF5wLQKY8WqpO6a5bsW//qB1L3
kBGxlzB7DjWhssxwbAK0Zt8cJA0k7nnCyGqmztRU5kyuRdDZcRdr4ynDj0FbhZ2/i/Cc6foqdgeK
gx8vjjkO9W2eT6O8LQ+pGDE2kn4VUsYIiypu8s1OU8WnfI4vnJcg02Q+uyoEeN/YqoxHzEJRfRD1
gM96mIBRMCwfBE6UgqYvws/ZKSoy2lGfmyt/6NZnzExJ0J0Q58Mv5gNB8c/xE/XalYvnvYc6ljGJ
EBuMdKBvfs4IZ3Te9vIUwL/PU76UfztMg6GlfmZQDt/qDHMfcu+Lc6YhajspVuqX20946eTsYAG9
DpeAP8NXlwVvtwQs2g++BQz/VSYatmZ+BLpoHmFfMJdU+LewKFtvXgX9nhpNKRa+pOU4Ytk4Na/k
CkLKAuhsaRrbd8Pp75hletu6M3geelhlMQKxoDwBvRhXAHKIOjjNHAJ/qd82pyuqLFpny4uP1QZ5
ekrkVrLzoUaHKO4xlCodLUmx1DEvd0KMLI6QL0sSoG6ZrABlX44O8I4wYhrEn8+McqU2KGFMtYJC
u6IZ2htHvDfNlRjGn2s1qJ/JzOEiDllWrT8VWYMLwbrzA51ENeCXOEuabk2lu7MOH2hwzhlAgPdk
/QEbrbpw768IhQhxJPgY19Zn20bPAB8tX5j0WXNp99m7d3VHEivUWOwUYkMZRxwQ74mamLrQd7tT
DhIDQXqPKCvqFVigTAH2Gmn70qoJjSmh0bfN5WhXf8tPC93zDjPs1z0HNmyo63jnhto5vz4w0rRa
FrKclrkzMD7yiDPn0wBEvU3ZY6/TwKvs2Z4D8vzfHOY2OEqHxsulLNEY21Uw0bhI1OwbKIJ9P7O6
z9bWj0s9AFSMxn9Ncxuow8wIyH3BxNNBqPeQwp3emAo6xjFMYpHmUdCyFjLrP32DeRvWcyYYHnOV
mcoUWoPfm9W78+OphrI4raf+m1xSQ4MqFP1aUEnO39q/plTQ6FkvYC1m2FGMkZVvS7ZpmuYZ/EqR
DAH9Arpxs+Mw2Gg77mXat8UrYlMNVqWax3Vz+afrCY6aJcS9attWpjhkKpnZvsLYZ9HIwjA/KgyN
uvrumMSNB8+8S8bsBB4hGc+2DWcnP+EqgsDFwH/VHkIoLn4E5UNR+oPhgwVMJpN+Rj+tlmS/lqUZ
OqKWvxcA4lt+k5agQDH5cwtSRKkwEz9XgJcNCDRd/nRjUm0h7lqoZRwAFhY1msHFrqMsa7GnxWqP
oKKUlfpx8DoPsVLiBzdJPlsKT6gTMFldlqvGLlITjnIuQ/KelQd2esZRHhvpLw8xC/C9Xk9gx8Ha
n0TL99agShhfHAt0niz/hrfRnqblf8klBU0x246lRSnw+vGhnPtgE6XDspZgjZ4TKRVTYX0OCSXa
ddD/sBSXLl+6XqZ/NvFwvOcF0eoPazMOCmRWB3C6yxOeuWV8T6qJlN0muiu/fSCOCuUKYxBVXQHp
ncIxcHdfCfYpoJ8XraVDjfdYoEjls8Fu5huowUhjM3n40/M9TENMBcaEFYv7h6lTB4/3UIPiGheZ
uF6KCMVfLw0GInib0p9oui2nI/MVPf7ShZinnusWkArIKYQkP7VH32TbRYha30wpDhH42g9u6wDo
malKvXuOYRoNTicqAWeaA8WdQcRVJ2n5vEBnH6oVZAIARZ5GrzTXIB4FMrqArKEQNRlN12sCr6pb
VOdcG8oBl4gtm0Q1jfm5ZigSN7NcMPhBXgR3jFYce2KL9D4Wxya1QtyFFkBqZy4cmG0cwYU3FG1x
WswNWSyS/X08eXihTGN7oAupyk9jXAlWgwCThMeWsW3dB2pqojGt48QWyQuZvJGuojwuhfWqXrWJ
xcUX2MwzIKqk5fMvw9Ps5lNtJHJvJA+qw6dlFNXwNmPRVfAlcEgkB1/C+vqUmQc5kOdFKcOtAN0q
WdjSLVHt6IlrZArqjf112K7e86SOX5RxyQJRdE4C7NkqYhUAm+RlI6z/NElQ4tSxxgh8P4m8Docx
wAhXVgNpVEgBFEhbEyQMwZKYMuewWeHuhpOtPoAnGKVDEbfejErUoBIQ2onWUOD4FaBqrEQG9I/q
m4uV1xjk/B+iBR9/k7ImDmroaxIMTG9wS6Vi11nsDSMNM9VwnruKeGdGYfATenbCOvvl0HDa8Q68
d/PRGQwFOSTHdD6cz0/fTfBZpbQIAL+m2qGtG4v/dRJeul8Ernoboy/qbhZlHKiFYlRi3lrS1XBP
l5FiFjAxfGrlmkwN7r3l7CXzvSlTkqmlZGynW0xVluTlG6tSZeU1iKNutfPIDpSa/5iz1AkGnjtK
9sgyvKoVub56a10ICNnD6eIYXBfzZh3yetPFH0SSI7EwkNl/f/RqOvh7TVZlamvJG+OUfdknJiBH
xUBvBC7vwsjhhLRGgnv6Vp1BZ+ZOzhGQ3OaFmHwfNb2eA1jJflA46QXs8D2SPOy3zCMl15VX0RwI
pUk4jYEd1v7fW/3Xr7KOY4aNgjFxkSqjVlBfKwsop9jn/9LbjYzizxt0PQxxMg42JDFvhROBmjAC
1QdC2aEuEqw10JfuGJ0ddfHNG38kWPKkVnp1vSODaWeZkvc1Wv50nGJDmWF7ctSVJSv3D55kID6B
pdeqNj+MfvZED4CtAmtNZOmukLrqa5XYn7F6MXTfuqAjJVx1ajCvXQ19RTn2G0FGAL/V0grmtfRn
aqoF4hn8zoMyOs5YN3MZFzFBr7UGN1jvekZjNwxENIzaT4weg7OjznFhamX5lY2d88MOOLuZooOV
dHM1jOLNBaUK0BtyTZCOmkHPkC4o0mdNWaRqSUC1YGGU2BIsZWLSzgoqvVX2fmA4bXxSC7XuJX8J
J7rOZLP70AGM3xe/NrQxjUJaE6J/r18jHBGvZg6yKnGsGk+T9wKZHXLkJbPOWnCJmGmzL1pYAUyQ
jE4g0K8VtKllcBzn3/CImZt3KfRMfcy+epGwJazWBDWxsPTDHfe/xY+zTOzRjqMpkbA3/yuPvCE0
U5KIHqRSu7jhvy407nFcgdqgHJUPkN91NbqLv9rdPx/1842bep8urdEzm4oWVKw3+HeSkQIv6Eve
QJ++O9+qt4YQnbZGIQ15rl60RcnvkDCw89M++iLLEOpYvHY1vbNuAEUpG0raWYpH81S1IXw+5lQf
8ghqnuomF+2L1a3+OxuBI8X8bQLM/tm0WH1h3m6Iwz+DPLB1xOWkshdUnUr7dBsyzbNZkEvEV1wZ
sUqz+4vccAflPwQqA7/MjsaXkwJpmJfv5cuSYqh6XfCsNW6hAvTmFgMr4oN8RyvtK2NiJ/VgLJ+X
s1kEFzRdxOLSelGtPGRoEyJAgoRrkDZ2jQvdCmB47ZqdGqCAAqc4k6Xc4tLNpCGRrxfdQn8y2Nm+
mQnfhIVsrBxldvpkKhTHl91vAWfTQHTrebis/mampjR3JYmh9B44r1CiQAe2+JAc2WNyuoLYAYwm
vr7Snmg8yJwbTM9lNyOYTjq2B8cNiEbX2+fb61dNkO39Pk9sKhkdOTKNVELqo5Szopu0h5QnQ59y
5u94pxdAAIdzgbyW/swKTsJS9/tCa3Ul5LcD3Pn1RlXCo9gTHA4QQKYmTxRxTj6y2JhN8oliuPOc
h9z7NrKX8wLCSStFDVqfI0LNJ3Flj5vhAODpWhVMH2dUoBzyP96ACzoK8zs0lAqVa5S8Crlcn2nA
k/yWWvdBQucMfxJMsN2slrEuTc9mjJuWezzRPRftCD+DGk+zuxy1ACiJmqS6vgXf3FWWJRBTnD6U
oElVeaXsjdI+y7RtWGGM0M3kE+ueOxxRm0VgurKy0ba1Fv4MmDgLEubmOBgW1VUMIRujiFsWe7Vw
+XhvF7EcMYk5/uM/r0dB87+8FeySSlMYifQn0TNH5vw9HKRh5czEG6jVhuhubE0SyLKnylndJnw8
K/ARm37HZ5tECSMgzPJGg1Te98fJeAz46uFJN9w/006nlFBKPxVv84dANSvK5eO01TRfg/mzoD2s
Wypwj0kQ2cvMf4ZTy3zS4GsnEmuicXT4zk0iLDf3ODQsFRBEzh/V5JHGzbUI7q9l/WTiHBrKE97m
0Hcqeg456six7epvPppw4fDUItDxUsKp5VFraIOHUNvkW7WuyUDptLD3VQcmnDyWUqsQPUHZUxwA
KLZTAIk/ntHRyMPhFWZOluivSYcS5BCsmsCC0pvwjpmhkVAUUTdJ3OBJvbDeyaJngEPNE2NTG/1y
BEOAhp5dM0B2DXfHpBtbJN5YqUWRwT54fJNjUNS7lSC70uSS/6ioDlwueZMJGOXS0kdjqNtIurjO
wIWqiG8IDs+Vk5w/0dG58RV2f8i+k28nLYqB79X5qEx0KI7RMclmDI/sfNuv7MNsPQIfOt8JTe/y
k336xGQ4FHXwPEbtocvGsQn2W4u3P+sfFd5yz7GnAvf09Pru+0fxDtTeOzhQQVYFp/JvSAxDnnqC
dbm9rI/9kWgj6Th4itGLdNMhEXMKYjI1BldsfoRsO6mn9RGYcbY0BmzaJfrpWOfaIEunCD6Q7VS4
dpaomeO1eLaWEC9bDseTGTG2zcxm812fASk4aNycFSqtZL7oErG84BsCF7A/IfcCjmQhg2lFhlxA
lY6hXfn/OR+guzlUS0v5lqPUhGIJ3RsThCPXYV3d3jB1jiQjNKW/sFx/DZGAbIQ4eQCC0+wNIKAj
YpT3aDtm7L7swbQprNWDZwoo7SJKuhua2/NOlITqNRIMzAqz2alaAlg/IqC2pVHPTB/LCyGHPWYK
xEsmcevCckbLCs03v+c1d6CM0VvNwRDnAuu3xUBaN+G/GsdhPQUzjmK7EORdd+6lNh4ViNvP94Bl
7rzc+YJ/hKFK+qQ6MGWHJjQrFN3/aYYfhJk2CqEpJPrNJe8DEp+HJW/7F4aPtz3SxnP2KGlYRF3f
b0a1+QtawdPDciZpXepoScLzODJiclhyyAwTkZ6v/K2BW+WHX3LWZLI3Gaa8OT5qUkX7IvPqootU
HbYoK3erc/LXc9BErfyjZe7uHcg/mwlB6LWLSFir670w68pWWSuMxLw3oMNDG3HCWHY+QI2kUjz6
uQFfc9LUZ6lbM5C+CS5B1zraW0ArE1EiyExrrnmXEQkyPBQ5EmY+XOIXFZwPxhzznh/P5UeA3n4e
tiL01xm+X7KhtbkEY+G7lIhynA3ejSE+34gVlsnpYE6HJEUPFXehmtUw6zeWBuqQJy7Sicr2phXR
o3D51Dp5hkjuVlPLpeVAqNnAFtBLnjf6hCiDca8+i+wDnVfVLZ55ck0tDoxQY+NW06r1AD+82+5v
Af4rh815RXr+/62jFs8UjoQiVAGSjy3fa0a0GsNPgFN7t2VOLbjphPdpAFl7gwrOg6rSceyZ2do0
gsSohonm05avfmReDlVm1K8jgs94GavNJ9TwpfxRaZ7k5C987bAtCCoJTSUzFLXYF+G6osC7rqJ5
dGO681WMu/IhAMvVo5nLiLVOWZWDxDOVVXiyIo7rLrBVeZ/r5d4FivQw9APCzZKJmAdCnJfsPsAR
fUR3sYYRRMwq0AnerZcK7AkiAPmMNDo8I9OYZXcjG867jcCXgkFp+ngYxgD5+8hcrjwwP/Xprhm6
MOaT08H5KX9ql6yTG/h88iG0MYDI7DkRm7LxJ7b8wogw21tQQ5/XdwBzmtadUZTFx/6zB5OcjKDa
PNCHgBDk3uTxD7x8wEUHBiGfCZz2j2GYnuprYzbv0PTv9YkbNYdSh1NPaz9r3LrAIr3qaNBEDtgz
xyQvsyzY7BL606s09qjo7awj0gRn7TD2XKFUIc6ZYqX5aPSdzDfnNCKx68PwX0WzRR1Iynsd1QY5
GHRtJ8EE05tDFDau31gIWWpAAHuIAz6j5gLurxlWuJKkH33e8oFGjX/SuXddeYe/D0jnzia/6ZqA
TEDlGeQ35B5aTRpB+SiTvGHQL38ihJqVSK7mZ0FNUPbJ13j1nRtnVulGHA3AtIo8on74OaICP3uZ
tBglxMGdu22J163L59vh7Wo/MPHF+hEnvb3g+WXbs4j9KcbRRouE4DI25R29uisZlOnvjso2Za/t
Z9y5ZRIS5+FjTHThJFqevxrMERNqZSUk+EtHXlo610JNXFybhAYm8lcWBzMwYwsBFVei4GzrSYoV
Amlv32XLu/TBwyr32GD8BIEU/hMBlLQEUz57xW2ZHvWsiRinJkKTu9Hl0kOONGCxdtYYj0JxeBXS
ldLnXLe5IKBRT8uhsgoeyLQOQiyUdlFQjFWZ3782LfhSGgb19samgSMS77VlG3cEXJ4uGZZvLDVT
l5A07Nbui4MUiSNqPOncUJ+0RoXem2cv0kw5iN7cJ4Dy/pPyVTfpPpKWHIUyR2YGxkWYHg65MxEZ
KDdW4SdwY6G7O0mF4/QpKheylskrL3g9VzftQX0+EmyURUUAruKChwXdo5vsqUhBSQ/j5bvYidCo
UbAl/iBKGHRYzx+koKS6xr1k24Z5MAi6z6rqEfi3QTgqFaGiA9vc7sHCxcNGACPeYWjhnHKHrhR+
TIkYdbGwBuKzaQQSXo3qih6po2iP5ymaj5B82rWKl9zg4GetcYOZ+7WlOuWkLjp2MChlnBwl9CWE
dA4+k04N67ngWuIEtP1okVODbnH4xb1SUZhsXLKImvv1l470erffH/GO1DH80DNoQOnuLb0UUtJf
awvV7xRht/tuLbpFM6sUOQMyr59CUoAhHw32vbJ8z6QbdjHZWEcY6l0mWmEdQVIkVcJk+9cHMMaj
CqSdRJiohHXnvFbhYV++FCBWnUfZki+Zr+hIGLG+U2Llkr3tF3Q+hKda9OB5sHLotTsF/mjtYv43
SpqDBwpTaiq4wIvfEjJ8Bn3k5XgGYedUfFXmT6MFY4wgKTrfScYKCtmCdlM1+zEvKduZDOvcSMXN
0Cb6nbb821qzpURLyoc5bHp0tl3ipvbjnXx5jSDoGk76EWr5GN5Rf6WEF9Z5szf7F8SG84Y7f7Qo
fTZptoHIGQ37ZxcGMjhPmKUrXeBtJ8UDi+PARVjT5VQgEwr7eaS8lXOal+IX4sr9ziJhz7u9vbxw
sIiXGC5um2ZT273ZA3jA7ZgTQslffADH8rehDjy/QL8si0Oef16GKv0zC/ZKWLnBIOCfBd9hVyD9
0D6N8rAHK/Dlv/lzETRPjxAlPNQQwTBYABUFGPrr/an9gjZR3/0haQyo+OA9ErRhzCO501oAOZJN
HOra7rkIO6ejd8/uYJe7zLWwHkA9BdrkE4vGjFjBReVEYvIMVe7DOJfxN7eWKLb1LRwSsUbU0Gmt
iTqEY4mj/HCOzg+dVEhQK8OBHGg+5GZ1wpdU2Yr9gZ6ZHnuNOZVQEhHPmWHvnlvPDY8c2n80VYl5
uXM7k4sk9lXPCGrz1HqPw4jMEgRqKKlzBZXs1x66cuJWLgwPW/ORD/M8DPLCwhwjYb531sjpl9EU
xNumjR8iC6bQ5ic5S+5NqupT7PYcrFZuFiOQ666YtdouNBZfyXtDVYcRXrV9ALGQZA33tbXrMpV9
U/dsZritUw0dfAT0+YS7i599JqPXYd5SkX4Wg9vaZW/vGRMjrn8RBxnOk4NKSMO3xA39ZmnDEFH0
vFCoe8Fmuo3LneY0KJ+XHQEun9Z7PTEDPDeXJymtZSSKCNrX5RvY7+fKLNofIcajXCMJRzA2RmVp
d8QCfFrEXlidoscwiEk2eXqP9nPVccwdJoqPaovsLr4AacGprBSOcjZm3yrV3PQGEYyFxUhCpVv9
NL3XDqMiWlo27y1HFvqU2BNsl1aR0HR+jEN/Y5wdetXDhGOuXd6xs5HfJcH92vnd6ak6BHOksBEp
S8D+F+7StB4OUVy6WrC2yifpG+zGtnGX7dHc/c4PdRVpcMq4IXWyCL/EbkeUgTJcmuSngaKcngd8
xJCngdznUqZkcJwA1bLGdKlbrQpI9urfWxYvgKlS4NLvZ4OVJ97sfql97r2Duv9kyUWyr6PELN0c
Bhxw1ACEp6vr3eur6k++Z/UzO55Y3KOseHOGYK508+8kChHP9pCzB82Hox6rMLLRHJZQKNikEPfS
miWbe2a8ZCbrVgjahK1Ojw4iEy9YJOjS/AUq6HU0pZYpbf3mWx7y/soDjqN0t5N+3Z7HkXHm/HgN
ONX29fJ830oIqSGa+uD1PDu3EJhZzZjrvmp2HNX40E2e+r4qeE+NlLrmN+X8KewuCv3RQ3Q2iePF
yiGihHsUEN87HjbdiUd/8UqTAj9nYHnz1iIHhS+YphAZRnXUG4XexR41xGKPugyWvuy7B6efNaaQ
S4l+3d3VJPTzLJiqAnLtF9E/jyhgGYXE1pDmsqbUyDBFVFxREbSE+d9Da1rRu3croLqabfiGe0sy
oV6B8HB3/jPybGZXhHpt069FJr0xbB/zkUcVfGGTJTPxiWDnMbwZIzt3e7gMK4btDOJFUMrp7025
/4f2pn6UQiSazKd/8NRk4lHSu83nqrGeklmm1v0Dx2XjIJhHl/piEhplokEvr0TBymO99j6su0dJ
IYAgUzpuQNjdQw6QHPZuNfnl4q6cIYqv0tv2hZplmKfcKYy+Ht+kILxB+RJsSu7NlCMpgckPkpwA
PEolZyo+/NjPt4ApxMTq+AjK+5Y6HDaAtaBW4UXqPQiX4TQ+8u5vnqF+76m4KPOPW7B+2xbWopeC
unnZCAAkwX6/9rtcBv5oIrUXByXTX6uP8fOz1cOJUv9MggmqDqdpTZeJi1wniQ8SqRGJEARk4Y1b
Ulck5kTxtrEH38P0Yh9LXjHI4i+3QqP5+bLs2dikCJAkZxLLaNXRNE0MXs1sbP9pBUo7hqaAbN35
kcD1Kjr/rQ7wqxD7h46usavcO47d+6CV81RM01FatmsQ4+VU1mTZ5h06E9C37kwrOpHTFhD9ddP4
R60Gw4wtxFbc3lfPQ31+agHgNXjwDU/OW19IOS8RGIaxxvog5G6OOx1ug2pPnEr6xrCLbbd0a2vp
aQ0GrudT4BLoTco8F3vL6GWDVkIpXTzZSw446wXSldimk/qMIh3IbpxrKIXGFdChvhln8eSwfA0D
1J63xPK9fAPxHaDLsuZDPMz7sLU3PU/s+C4m9wOOi7HwsMsbI+UJ7HJJQK43+gxbLoOzjcLtqVya
P9jxZsJrfYQfXRfrQhXQwtXhaJtG6jkt5Zcj5pgzsaPZJVEpIR5nuyJbug2B3zgc4pMIL6nblMvl
DBYQAsDxPQ5OTbsnQESQlA2KefZmXNCCJbn4SX+ifbBIjde27cIop3LCbUp9XHi+Q1Dn7+Poeb4P
9H7looraptjeC89uJ1IR0pFoixQTFYR7wbMB2Q+6zNHf3Feq5b8JKY26p+6P6xaAJ2Gf2OyrAMtP
eE1vV6HBaEPshp/TWxOQONwh6XGsVbpLneadXQ33pV04yzy8YcJ+NQElM+PK3qfonOwZehwhuMp0
/STMrqsBDMsA7R27Jl96iPHm4CMcrlaZRgfDf9lbGAAc0aUozDdP0nUqcWCQos34feS8qYPdpk/z
bctlsICWiYDSWw0PQCMpXGdczQ4Lr/mmZ3k9j6lfKgiZ9dDX7+sUXXlHbp3keHy50nJg6rYKQgKR
2t+pp1JYp/p+mt07BueEnH6wPGoQHRfIkt2zDJj5CUbJMqzH8TsFTRjBCoRDmUcRHa0IUIQcwpX+
4H+zE+yO1eKv4OTj6SNZ70j/qL7tO3/XA5/Jg9VFYXW136PPNwO5LOJP6L4sYUNq+/OrhicCquSr
KimV2ca1USW9RvKXFfyE5Y5TvgRVl27hTq1joxSpgxsxct6lD+vIFKmCoDm8xbejL2447oz8h6Ib
jnZADafEDMTXhS/6ctPI7KKT6M8iIE1Wqwvp0V6o+kjNqGGc5CPckNflCFt2HuHUQa7TAGoDK73L
KT6FYxMT2JuWj6qSSMBmcAM96rvP2KhUpmHzdqHoEcsem8d8GG/XcTKYG5LGQtNm4LXqjPjIvVZ1
ozLE6pnNwSpXkK2kw47IWdrxrIwmZv5AL8Iy8TZsn9EafleegQvEjlBCwvEAAy91k+Y1T1sarw4a
Wwu4jMS8RucApmbJ0g63hai8/0cBjOHAPLQREvqT0SNx7HLNrKaDfESWkjQyMzt/VzOndbXSSAg6
RUitYiZ5NPtZQ+VOqSMH+xm4BAC/mt5i11bM1Km6DxxI+WyeuQ1CEy+cBgikhpnDUjq/qxzyZEHd
FMYN4CIkdmytHfoEQHiCM7+tdpryyjEZhSsIw+LAfp1y8BV3NHd7UhRS+2mSt0bs8T4W7ymp+Itj
g10VApoRH99D+Xa81HB+DOClkhdF8ExkhRUq+v9FuTTXzasQ7BPA7Z+66kuMrHQn8UudHlKf1CdO
xL6QeWoh7WOMkEuTqfkmGvucNW/wBBK7zcn5CRQ3KSAKHw/J6MK7zRA659o0jCFCOBP9zTOjrCdV
UDqu3DvkJdUeGabBhWe6GKbWgTz7DpQH81D17T+PG8/BsmrjOxI2usQYOUtEj8AKXyXU/TI83nvD
iCj5py7PtsdPMLwP2y+zMFMWNaNxC9IdJBlGuGoII5jp3QBg090IhB8v1g5aJnIrasYLhAEfgkka
xZfqY2mwHIgPF/1Recjo/u7EDWIn/7XN6RPYF1uAA/vVUkIbOozMpN0r8YPqcZBdWDoMpkW3Blta
0S1c3UocIa14TRaTAkZBc7vPwbsr3G/CAUHymuBpEGKgs1quG64uG0hHeeGtl+2+/WOa8H+MLXG0
6IdLHqReFxWAO02rZNkXOe/ZKklRIyv8mAAB7FnUaUfKLCoegbR4gLAtJ22qSDLD0m8NNv+djbXC
6k8BFuGiV3FjYMJk527sog+m51umQhzIPQMBu77KJdvIdFyoOj5bbhdL5/jaV6PzN9kIp1FCnjR6
WDGeJmH3JkWQaCTmlg/zCkFPTrRbJBWPuIXP8gxRWU5uXLJx5/zlYk0l8dv5epXhkxcQeTtQmOjX
oscKdWYX981JsqEAQ6CczPxPxBtQQL09EdSX/Os1QFF0V9enp4T5QSkoZMAGKf3gBow77idk8RK/
Ylh2z69VZwZ506OblGSjY2qwkI3Cw0sxK+WDmBft3z/G6dLs9r88clUVU18+/AUSY0383NdWXg26
1W/zGVqUVYnWzCOTzmdcWADrI1zXufYL0ekFTlTTg0Gx2kgy9Bu6R0lOO20pnkIXzRitnKpILxp9
d5v+1z7IVqB90lK54mwa8HhozqP5a7fhAefMjd5sQFoCEFXakuTBoLMGYM/3H+5atS7vzWO5cztF
wu1wRTrAFU3grM+yRkGNfPHAHVzLcI3Em7oH2G2VwEGkkvJquP/RFH4aMot2SxHzVDUW7FG/3dA2
xi+ISsfks++mDxoxeps+fqUOaaByMMLBBLBK+eNsdL8hedUXSUcAOyVpav2udXpBN8l8ZhfvQoFm
B1EXm/Rnq3zrV7CNzLD0UlKtvw0DvVaB+ds1xmOY3yv3CvVYrZZatHU694m2YV9JPrwILJKQuxfE
4zXyfLdyRFVTS/wkjl9dCSu+AT3Ckavt8lI4j3YL043zNPF/h8O6rlrxiA1Jr5jr4VgeQTdE2fN9
haNS06XgeMbLR3xBIElUZzTcIcc0xe0F+rPHcsQfvwgWbMGuog1rLOV23/Hb/mT5q/Ej0NGhFoiX
kMJjxAzDeG5pGeyPLI7Jkdn8vP+EiyYalNYXioCDIABXsEvd0gUJ4n5rhTd2cWDeLFiuv84VbslC
BWvUn3i2FrtJCgB6wrccN/2Vy+42d2N3uvKlMNDdm8xtwoFKnvSpUaQKOOH9Wnilm7yUuB+JEEKq
G69Sl8K5QD0EG4bQT6HUchp6xuqs8FOFEPIQKzMozwlr7Area9MSToBSurmO4IyPHwKEpEvQ3TbL
faG7JLRpH2V/GV5IhJ7KutGxWOYdPV9kFdCMu0vhb0PEjv0pb89OM+kdq3jWMtU69VztATl2jwr+
8RJenuXb7BR6PfAtr1Yb74R1VqLb7vpc+7UId6noXQ82v1pHmevsJf7BqCmAQFXyCoGqiEdrGHrn
pj1SjWh8WPGTa3xNIqSD3cPu97atvIBLwa23z6pqMOWgBeFOIcp5MV1UqCN+TDWZb70UBaqLVRIe
jnTRISqu310MOHK1ctDhhh4njxdI0hMbD4yreH4C7C9PTJ0bi9jQulf/Ia54NEbzjwijRRNrSpQH
DDrycay3yZFsSxuptfvozPiCqVGSM43zeN+YYo1O5DlYSszc0CCH08933lydwma0U1TGH3kE9hAk
lgTgElGl56aUqcfkcJh7/E4i6yFdxk0X+mngx9YdCK0GtpYIJt41XZFrFEGO287xOcdU40XXwlwU
hS6T556Wv/QZq1cOzB6Wfet61klUL7O6nBeL7ollfeOZLdmCTsOtGXxvjIXg6tkMP/tC6smj2CYj
PGkOeY8j8OmuWEJR6LWaKzF+4h89rLr8VwOSa1mNHVnb9v8TrNYBLOpDKablt0gOnXG8N0qh0VW2
uJr5DHGUL1VbF0UE37tsRJ10x+TklBps7bHWKb9b475TTpy77miXzC6fmj8iy7nUfmMGrSgEeXsj
UNJK8sYYpNQpKkZNQh5dhiMUauXpJEUmRrYhxx/l0nO5SPtyqoAD7WnXFbfSeXZUfOCLM4YBpAUJ
6PdFP9Bu1wRAfEs6f73eSjOmTnRvfuV2C20Nd5cs0C0lGN4ZCmuvbDNmN36AVwy0FP+fvKt4NAA1
SQFlNpsMEMAPwGyaHRHrz4jff0G0LfprM8Kh3HyAEFkMwIUl6P35BFFoCWeKfkZuWTU8xZ7nhyOO
2tAAuesUV/IX3Ji5yXrSnvr7SQWjxjGd8bewkQw5Mu84q9xqLs9OBOmEYOua7VoTMD1L5Q7WMEG7
vPA42fjXVPzD3SD01YNGYgQWdkNr2Nx7arewKocRDvIL199FcszNCKpBb+6d/BBWVhPf2csaPAeN
M6cbJ+mZmWvs4fvaO/i5by1YORPiHJE1gzv9Yri5x/jt0TmLbwM/M4HqvtOZH6YZo+wLXvnIC7vL
iGtw/8q1TRPCvOtZU8wCieWTQg/stx+F+e4nGandy8bSf60kc9/eyChpVOL+W0Z/fm+Ir2UH4if8
EqPl2yXa7PZJH6RBN9/XAopKCVRDjV6PDkWhAhTLncroiCtwgVG7qVYlfXCvg7/JRvnSRJdKDe9D
VRqDiJ3mdZWmEcXn99nVI0jjYNkuzDk9lOECkraQO/IoNSGu9TEHv47QCRWymJMkf4V90+gN+tF1
mSEysc574DFhfoeRpBvkBr3iJA7/3kiXOBRFpjTNQFnU+CgE4b1EHOLGhW1O+7MH8lEtliiiVmC9
WKo4n1yAEwYkzU3J50k1CuzhJLYlORsUv9pvwXgbVipVGBkE/GATtClcKEhz4FO1UsVKaG7s2kz5
LEx7vq3tNTRs/V3y+hVrEDwPlbjKhJHbnCP2OpsxQ1eEFMATNNQEFtC35QVB40PfVeCWNLK0wNe/
gF/ZPKF9mKNv484lrZfsGaYvvOepY2DxjpBxmzKgfNlaYeS8zgsoVTnekN4kwK2pUFsYYoGCkNfO
HCX2qMvy3joNDQD/Pf4UmeWSoxk8r9Hewlv/EPFtec1rhfNtGR7dMpaPfNsKOt5DSLg8gqa7gJ+f
6nFgth0ywvC6jNFvfNlX5YJApAyaH+ViM3+Uiah19zrWYXicwjbcZLhjWzNKgZe/lF3xHY6sUcpk
ur6N9GAvoJg3V8WUI7ie9HmCY2Xljtl4Faa3euGutJxDQt+AnQLlur1Dd7yMzSFM1/d8nmi53RUw
HJOJ0nG19v8OMOVIYlshJ7edcGlXory/rI6dMzNlRYK/0nXWYovbM72h3ue4jUOK3CE9uzsPo04O
adBvDFKd3Ls4IU3OXoX+3rvr6AO8XW98MBmAk2uUrsjs8KvkHSZR3CQAqVctjI+AA7zAj6hCnqjQ
YNCQfYKBLA76uC0XU2RjWap0wF1VMEgTVaE0jv4j0ZNoaoMx2b7DGq6CevU+AM5noVpsk3BflsOe
jkKwpOMTPijtkcb04maG6yQ7X0Xc9ph9X9WkrN69kG2H7QNuQzC7BDzBaAMVxDS7Xm+Md2fGBwMH
1aWKNNMkJiGXOjikKtCcMm94wKLu5G9SQNp0gOX2OXjQ/bymWiTZrN0561RdSxZFdB9LVRvEeC/q
0BiJ+k+BqJLR/mHdP5AQix2PLHWtxPltmd0BhRyY1S4FoZZM26nHWOoJ5Ndnbr1MsVp1G8BWpm09
739hm77pOnFFPq6q9ecjZeMRruaNYMfzmE+sJiHOyUe/DmkJe7HS5saLqT4qmpPXihqUixZwZ0wk
jj0xZj0P27tUVEvTBx5EIce8nNczcK4H1fBPzp+sGMKmlwS4V7cfTd0LO448QlzCoPtWEXNKnZtC
0+jY+BBZw9wegkq6f+V6pNMliMul1Spy/VfBdNveCWP7gSz7UXNbcePqWmVPuZn8rSivwBDY3CR5
HsLsFY4V/TS7xehKrGVoJAfD7vSMtu2vUMGc30Gyhq/WbdlyDOAH8/dPuTz3PKXC24NO8eDsRstI
A7r+/5ARXOIX5vpR10Fe9qtLogeBbtEjVLmOxvcqTf/OYEX3GDUZLLwguhpSYagC6x77NCkyEURL
/8tKLIGJERkb6T3JNiHBZoiJGZtMMnkOu5GUuRezhdE3FQRMZywOdJE88DxzmC+gUqC+ke21whiT
qCmn7MsFV9qLZUsAZrKLbd+RvQkaZeDZSTdNzwSn0bQE5lFtLxzYwslUUyGGPLPnOWdv/z+aP0Wx
APnDNTcTeC4ZMrXqdWNzBtDIiE4HjspGaWOznwZPTOzJlzx9Z4uX0SbGsv2GsS8kQKHPSaZXMjuS
5/xZ1FX8UhnF+UOEd1So7YQbXXlKN6iELV9AMyAGoTv9CWp39MV1bvqF171BtT1lPIcWVlWKLIAa
a54UbrJcrAuChZauNZjCdYlT4a2AVk788dIvjjISK4ylP3nPhH32XMStfrQ/szr4ya6vX4H0UC78
iJatof6oqZrtJ33orkfPvqgnK3YO4SLL9IjrZxx8/6nl+Iy1U5YsMbR8GNL60WLbSmr/D0Wzv60l
NTIbbwtkU0FtPvZQZgA0gV8OK5GwH9AEhEEyGy57hpshgg6u1QT/Rx70W9d5lq7RLfEOgX1BjxJ1
XuakigmycNE0nFHJ06ZKnbhN2kM5CLbSBqi4eM1ARR67aoxlhABmnv7vwaj0fkkL5mC3WZ+jklJN
hxA5ynoeOjjj51wGkdLY0+We0UtZbHyPpJ3NhmHNBLXo9UgTy/gRLDbxWLdPhlCH4oIG2/hZnXRs
sTOK9yD5dMlZGUkTzXy0wbRvNvFbJUOIXilkyS1Q+cj3loyB4h3iqrU1Mfgv1M0/hBoV9Q01Y+LX
FyzgtTvKW9tu2r5WOEYinKY2NOMfnqbU4Qgp71AQyZfXQASLaQDKKen5hxjhoF1270Ta4FHz+fuu
zi0KBUJFVhahasbeNST+htlAjXzPa7oDZ9fFycOR4uPTuUdpdR0+wKHoFpnIlgMAs+tp1bxyn4+H
tVxLVz4PDje6whx5xrJg2tqfby59dqTfdvv9auWDz9H0z648L/RrUCVpz08yVSlNW56U0vI7ekRe
jPRUTAeukICB2fLVD+vcLSHVErIwRlskHiuH092GzsR5WjIh3qTSUK2I0JJHsn2XAc6YSL3X2T6M
muEwTDXdZABrA+dgtcUXxD9M4JQIWbcmY6CAXYsVdWTngR4LGl7+ccTqhBdeNuoqfxCyPhQElt+F
0rCpm6l7DOgM0syoYeNNJk5wEmesKZo7YbDoW+GCbhIKd7ICZDaRvBE+GC+o++fw50pBcMbKjMp5
rnhIdWKFVOrRuYf0M6/XmIsGGX4XemvFEGqzeNRXGQz5GaSm9buGzsaK2HVxprLwJM9VIdAA1ky7
lJcfImWnHR4rzLPvAIqL3qtlK8/8RZt5g57NC4zDKvxOdaqAZutz12NuCsuAtnYEbUwnkLg0+/Vt
PF9VGEZmKm/cJLP8tbPtLINLXh3zjKFKV6k4+HbPEVunH9P63KlnfFZ+/bUXtpjYV31kbAmAr4aY
KJM4eK9bkP1ytt0B2tgz+8RU8z30KOsyQGqqd29GUBYIFQ/Vqj1S198UHJi+q5np/X65mO0/6GlN
mvkDWjcRzjS7BDFVCM7GvMGT1iy3SiPsAtwsCT2tYDbNoAcrhI1+xF4FsELMC5y0ZuhAuyJj+MG6
o3dRCElcssEelUo1pK9o4cpM1DuY+CgQtqbxywzpdVZSbVujPeHQcWBJUfzAh31JZDBgrbZGjEfj
gc7eyx7jGPuUpwOVj5EuFr4qO8wtdUiio4nBCAmZ5vJ3YGmKGfKSL1nXXSfLALBnfymIKyJXa6hU
ptepoyDM43egRX+b0f2MRIsqUK0d5irOeRTPkFeOt+mri1gVpS0d8C+biGDQJdJFK+n8R2d7nNsN
ETO05Q311wqaSIA03TVSX5P7MUNgfTpVflmn/gnB/ebDuwdAY5Vng+Q10T5vOIZsjLbwYb2xZ0n5
U07sSl8SiOg+5kaTHT5HbGbXOkMbKu9vmbN/dmlbLUHDtEZraYdhKSZLLX8pNUx87U32ICULjaez
h0vSnZnK3GKgHHswBv/xYsD8tNXASqRK5dgg1j0YgMy0Q0zp2saFR+hCeQG4jEqnxcPJcptfn1b1
E64Dp7cm/hE+tIp9n6+TDPRyUc01JoQP61WV6P6HFk3wEMjH3I9ZB7XdZQthubkVxkIBHSBvo5qv
55WJvyAXcbhSuCa309Ked2xEnmDJ7pFkDn1UURGLPad8kif41fJLH5v1AnmyMQbsJ02Y+7xV0aWC
FrtKebERAD+d0aOluAsXsBBYKSChUsVBbpjiyCXWapZizn66V0KZU0+6bJkxcVFjkgiM4sS5f3DL
z/WfGt7II+Ut/vwPGYuV9ahVFiRQTR0wS0InBcxTcK+9AcB3FXMyoman3TXjLLD0tJG+y510BpKS
u1OnkSzzjS/b6JhxWSY8amGXUVbXVw5Dfrj2wfk/Wj9Jq9c+KASpMVYxp/CkpGUCZ2h4ledK0NV8
puZUagLVOCodBk5+lyHgEzFS9eyv8Im2Aglb0f1aHa2AG7opRWvAXLM5ansHsRCjM/KoHPO8BqY0
twg6WW2jQqZ/ofcGVVl1GUz4u0XvhJmn4rVxdrKQBPkZKpZI6ndOsgeXBkh3kpcCbmpAjdVn+KTa
9z82yDk2jP88Ssh00d3d2O5SLPRrMHJsYkUoUbRrTTbbY2FR5mBCRppolH9hgulFrWpldJH+a57x
PdT5nd1vvPaXLOj8n+ihCL1/qnf87f5h9kvNygFVtyJd9/6vSCqvWlKEi1sQl2KDFOViy5T88pyA
w4YtXRVJUtXRnxW7wSmd41jUA+zQRXFQwqFyw8MtaugMz1UL7bG9flrRigR4AEXEx+qUVeuAJbCm
Dw2D4NqyjmGCvP3T+YGlMAQW9UA1S3OuN8tX0pcEx0qErGyDmKvRalqPS9VLC1soHkwPVrSAqIrO
owb9mIPx3HCVUZjcVYDDmNuPVV+Ilp5YSXtivChWv5MD36E2ASxqINPNtfrVpK2z2YYDnWyqGor6
1+bFyW70SmfI/H9f9YxA0UIXpC4iXhPmCyLWE0hZvSBrUMQeE9d88YLwnvW7nwj7QabFiGsDV7q5
1+m2eDFBxbp5ZxdsSD3XJOwDM34fO+yHSmbXjoEPeFPxwg95esALkBQnprcWg0riG6cHRPCbkKWA
P0kfYmZ9odtds/yePSCjtRZ3tDJqwmWKKRxe+PRoJ6UyFIjiOnH78sfPFtdEBPyD9GjOb6bVlIkV
nidlhFpnGEv53yC+6XFk5SQOI3ueciF9uXYJnrBLdQ8n0pzOX/+qme915ezLp+OQPQSJI5LD+lNt
1q800OouPUZR+jUkeu+6/M63gZj3BiZYCPY1E1mMz/4zlMn5O05JYuV+9F7Lszx0KAK5RWcZvuq6
dP0p4sKt+VWdYjvZN9k0s1zEVVgqDROzRU8Q7yEpT0/6xJNzVBcsGxujEf7pzGa9SU83cMaQJDeI
nBage8i3xzSlF0trdaTaQHtJF0T2azTZvVlsyvHM0i1ASCVlIl1+Rf3RJW1xb47Hi21/ADSlXEux
JmO0iCCv+W9dPH7oTdUh6pbcQZEUiObcKfLk/dJW5InQikfg3GT9jpAOzz0ZxwlUQr27sfpl2KmZ
WBdShgnkl1lEell+JlhtFtcFX7taqBB1O5h+XfuuykfexEmzUtzeuR8S6LKH1Lf9A+Vrz9LBXueS
sowUKtT6xD1nKKdhlzhbIRD0KeXRz71lWoa4pu3s81921IqQv0i0Vttbe7p1FFe93NYrb0UxNCMb
iwr/RxeUG9EW9V4c69XAsZEPYgk6Z1i2PNTR3tOQwY277x7s1iYfal6INznLCb4Cq/EQjjdx11Rs
0t4fkZE1RGKNT44/SDftBMzxM/SBSvZKN7KZDWqZ+gyFpUR2vRrE1vYpXb8NOvsmvmkEkD8XqC1V
oYBh48WZcLa5s1IFw0h/vlNYNig5tD/fKlAswHTf/+Yv+uAT4KV98YnwWWDl7q1Kvk2YiOY1eb2H
LoIQdBP99ekXdvBdO1FWooI9zwaRnodGTUvjhKbvxamFVh271ssrdvnaIwtaIcuYYy9/YTfoaQwJ
JkQC0yQVPu8/urkBoB5JrbWJhRSiOGm5H+CUuf8EjNcQAuWka0/xOOPToSd7DmkOZkELVDCFdF77
eUOk0C/yUTczwaCUHgu/hCMvtiiUJE2eDwgzwS7GeG27A+Co1vq8L+sXbf5mJU/rNaSgEn7YoxAY
GsQgkomnbWGN6fmlRFQ1uk9m6TzzGd+w2IRPelVxqBHLQqaqfT3SZ61GO45GC3/kcF4NUWpSFeWm
mwOdJOMTLcXlGzgpUiD17fAuq8pMCEYptzlnRe9De986s4JjIJxY/1k86bxEv/j1kKWM2zupSven
Tb43RwoBPEtw4Mu7jd2xKaHJXYyVtdZAeaxnIUC7N3eSQpHjDsEGuSqRTSzgn4UNXqbBQbe3B5sv
+0tCYTX26mTOlzEK8DhDLqEr3jv0h+gUf7/GrPSqs8psYXvBd5pLw/Iv0qiFqX8ZJOQN+iq3zgPo
WFIiAh8zP1QveoD7YSsdtED7x18OHZxwdmTO7aLNWyexFEtJG97a2UJmC+7EnpnQ8KIpeUfWj4IQ
sxOELGB0m5+fJBEa+jSOhXb/ya8IhIi7d5ZiYMAlJIMgJXBPQyZ76cBCIpR5BPUKjJ0DGgkbprZk
vseOZ+RLb5p7RKaiQQcpBIkzS6ll4AK70JnVvsF8D3wrNLyLCVcXv0P8QgNLjTL/TbdDjqoRAbLU
K2qwwxjqozho+rbiInIvcxtmgvs0d79ZSkkxRp0yi6tDmnpMXfGeSL9uPm66lFqO9KLO8aSNSwFs
iJTPFW+9I727+eJ0NF7CnIh3r09oXJ4Ad4tgVd/CTYmiQL71Uh2rMFiLNYBHZuyA9YXCBnNG/mHT
NT4zlrNhHcrEJDqunclcjdrrQeuZPQppu74OS8hTWG6i410XceCrE9LgqBhHRx3+Q1NNaTPGvGlI
R8vRdA4H8RWCChWpwDCvlTohEpxxONFQC1KIqQ/SdSHqEySbmsn4WhCHqb3mKlbmKfVf8qUCBMZY
zU7HMxSRfKZUGff+FoyuuXwt2vkmrm5mHiKaHEWOybDCiXkJqtF/kNQ3HePvwp3eTZajEyMCIXED
Ax89gUMMjq9MQTbbxvx47iWan/a6l0VS/Grfd2nsL8ufVj2AvBCuO87hC4tzdiHyQ63wWYQIh6V1
Kve5mT5pLX5FPGPuWw/2p8G/+X+jiC4pjkbBsR/C5Z8ABu+OxXLvWROqzsAzvAUFcmMKsLM0qYSr
xQKUD+rYDz7cDR70tJ8Dct5mOR1WHjxbiqK5cwhFb4yGMuIbUOEhyI3tQH3UBB6SDCWnadmf+UUX
Y6VyMqUcvPr1w5m+d/d4GuemuPvDj3y1+u/9aNut8f/g7z5c0hvBBM9qzkif44Hz1MQttrvRmdtj
6y0MdpeyB6jUxGPpMse+6aOavB0w0LGTlzfV7/n4uXA/hIi2KVMJX9cPtxOcTyO3beQyNHbfC8lj
apdMCpCo58CBgCJzOIQejxn22MbBpAuDkUPHpp8y7vKpQ98J7kGNwROC/qYGGeR5GzbApUUmplRf
D9Efmss8xQ6SDHM4hzTW+wJ6BsnOfvoTHyIug1aDUjemtdGLWuDnyDBduPCB20j8BJHL6UEtKDjt
YXXF8ekGidarEjYrOkpRYtrXEpkXUtEtPwEey/OBs9NxoW9vT3d/Bl8TXM2QzAaMfbS7u3KrKuAI
9Qw/Xajg9N0Q464L6O5bPuF0RpeupUXr/Zmw2H7J/MvdcKpCaE8nagrtrK4+5LrMZzNQelK8Rruu
U3/a24go3v0P4b7ieitt0h5BY+/sxjgVK7SkJ4EaqGyfDuNPAssX9P4C4Ray9C6mCp6P6NZqbOSd
KWK1dujoqj5Guw9FXcwsaVQw8xIrSsrhOalPFf9MhR1FMFIdepTSas4FCg/gS4TJ2i9qY0QKQlQf
UvkBSm8zEdeoNNBRBQpfqF+n0JxzHMXP7ck/F58clGnYI8f+PqZ4MhYeMtCu6ew6k3UokApSW1Od
sCnwm/UKRB96HHgMRy2Mb8CoJ9wM2wDZpn2/D7MoWgxsS19PRgFiR2x4rh016r0r/Nmx3egbuULS
zBCJUMQiijhr0eYt59mrP5iF91RL5UvBeb8o0eA2gH6lc2zMByQLX+j6C+LE78GP85z4IHxt6h/y
eyI1025bxMjGtpXk6/YMog8XWCRboaXGH/2SJQZJNMka/BU11SRComH/rmQe878ymCEOjxMJ9hFL
CKVHtbWRRmBe0Ws/QLAH0ccX0tO80C1235Wv24qJTeWyN+lulQe8iiu3o5yk+uVKfBT9/YEJI/nG
jFxgtQQaWKp1BFLO29V1UQH7aPk750Q9U3GrCFLaukPUE+k7XcqM8tFccb8uDj5nOlLw0fI621PU
9dKrUQbwaPBge+tv+aAShkYHRpYkjb89p3BnbK312CSfO0BPMj6GcWCUbAWk74qE5uQc0q3E7rCP
gxXpY9TIk+CMH1yQne1/zNmPKDuvOvBhxBmLBYfpHc1QUpyAnYv4upjfL1bLnkqYzxwJ5DipJnKC
NcRwY23ZYODnCfhFu/jbpsVnzVZW2FtbS/1jlMDNoDcOqvnGUEoy0lxe9mjnj8FJJQcXkIsxqpBZ
chb9sSjjOuqqZ8um2Cm8Uj4+/edFcJPD/mVkSIog7kHmREg6y+JkYN8n2wHsSJia6zjjlh6gufG7
NiVD7XE2MhxHVA9EFVoeu8tOtTn/iW3vC2RMYUTAvuvnNiPVqzNbG/TaoKS7uxWCh5cnhFzFQPOu
4e6o6d4F0TmiukbdwYtNmyL51i5yK6H4fnkeuLuEr235tW6WlvleFKbN/6xlKwasDM287F2pTFq2
etKsaB1D/qUDgF+orHNvWmgPjOXelAQJtsz2VVwCd6HjbonL/FpLx/nFUfKcQwfATrbZ6F8rkdbA
djgsfsDzwIN24YGZSUKgkYlQwmj1x69/6MDGsqWQ9eYb9tozo2k/iOtRyWH+b+UHotJE6tGwVF8o
xT4NSxkzFrfGOkKPdPHjPRNeXnknWj7aLoXlt5NX8HoV9nXxFmTOezOiWg2rARX4ea45I1oeFQrj
Wnu4vMQyMNXJT01T5+3AtVePeJT+XgsiaKAOQdDgFDgSndSplRDRKfErKXOeM3inhy1otLmZB9TM
NgcwP5D4PTKyolrxv0+enIfQyjsS3N82NFTJ36IH1ZjjPCWUZhm/c4wxz/bhjgU6fGFaFkZrxOCx
a1k+XGSgKA1zsEosIQig4Ou5+vE9nC+2Y35U8/NucttUN2+4Ub7oQz4Sl8eRFNsWXS6GrMf/Zs6r
q2iRmcpT0GOxuL93nfYeLCSnSz5fIEHhZ4+Nq/cdnkhnP74tt3CZFdQd7h9FFWTkFxCPSEly/ghV
YRqFLjpYN25L4XX10y1ifIQ6MUoQ7n/R+P5rJcALFqI8YkwcSHtYNG+SHK7orSCRVYvtPgj0Rodo
e+aoWN4qBxNIPEl9NFBSNVv/SjomIZgvZgeGpwhbs5p8pZKrHMRgJe2zuMQbQsXWjR4KBSWiHrBi
TunfJl6gGGVTS7ivUC8sYq6lgufH71T4aY6+323MXbK2ok6//wnhv4veZrKirSDOtD3kLQGUpojE
IcHBdk2HwSl0i/QWV67ACRZcPHBy5YoPH89Vr9G0gAaHfIi/A7vZOQRnRZRgCbdIHh6GpslAj+nt
QDFrYPpHqFVPd09u7tUuelqOJ3AKoKCfeT9vMIxRfzhuFsX4010GvR9QInKv/5gK8wL6vT1+Zuhu
7JXS2KeuL6cez9S9SnD5R/o1Xt4h9Gy0tInQPdAiSx7n+y462E4dULA9LqQgmua+ba9I7S7qglpu
IMsk4An3a98o+HuvdXFprW5GJck6+JN+Kjtb0B4XT/lcl6gmdbMyHAHtfaondqPpVwtFlPSAYsqL
J/3Z4rxEWQ/pMVz49dwhAx/lO7iErZN6FQad9ad2JydU6XpNe2GjI/PKk27m3HgeJaMcbBFGCMa7
ZOkPXOO/en+b4K1foporRKDP3ZWDDySLa3692wZe2VZRlhZz9LxkFSFdjymWkyrhED6qhaf3o71l
rqLRNSTiwqXPuOOgbtXwLD2qj+xeBUZ8PdzzQqlk9T73nQ2VdvdPTk1QesPW0WZnN5SWiW2fvX8a
oO70+CEnih0Gj+4yZzpu2S5G+fyPhMxsIjqQHtztSSBSqnzQ5BE3P5BB+8z/yfh56e/U7Sps05kz
XaQdAhs5JE5mim2ald1ImYFHW9szKlS72bXfVsnGZseik5aIsBntCH0OXHKLQ4SbiEWMEfOF9w1K
frT+BkeGudImacgiEkKJ2wv+CkeOb4B9gsLvWB9vNPVag7UPs/mdXhikJ5EjIZ9ZO7AOfjeOOtxV
ij/JZxvVN1giT7XRlfWXrszGICaR/nOZ1CduDHu7oN9Cva97jqPpacQ9iS54ah7cj7k/qh7A4W89
4B3LbqitIREG8PZoNgX1HXQz3+HNoiZ22UdHMoc3PXpAwW08nAuoCSL7CX1lMJMROzNgmIDu5Kn4
DIPHurJygc48qbSas5TTttWRI49mjIEL8dBDs/It+570qJq4TsJUE5G76Qksbtch92PoP274gMDO
3cxEJXqv1K9qFYWBMQylxNEqdXDHiC2EzELHxgSGBtdzxxcRqzNx/b0i1PbZ3H+anRyxp2KV31HP
pHZVZ838tpNS33friaizdaolnGhqsJzhLx0drmIyITcr/kDaaxP9O5atJGDFsaAou3XeIeDGbrmH
W1dru5ou9jtUi85QUNN5CdWEc+q1RSlJdT//78aCBlH830LA7JI+9J5sMvR3UuZcfpvOQrCP3/ll
u13SssHOaLiN/S+Q6hMt7LP0Vr4fkwXGmrzX5eKnHcT/sFKDhp3EDeYH7NmGyqMRJcWATW87cpfv
if37gBCiyE7fcgV3VRnXYkuiHYTN5ml2HCTzaGT8O8NcDjIGsp8CjXUiFKVJPgQgCB0MQPW7aX73
sZWuMRr8SgXnlSBzCK+gSrNU4A7gyFNqvmUyamY0FDk8IXOvdhTtPoLAgzGn/JF6F/O7fsyZ55SM
5t1AZQKvQP1S16+zypc/w5k4rgimw1CNkoVi0KubPOqk6XBdcO+/aFVSuDU+vbRghv2423V0A5Hz
M9P9ob+zAxdhlMe6Upoe6/1IEFKZNjR8wmgrkI6v/5N2hRytrf181VwGnkf9it/C3zF6NYYMGM3O
OfJWUjQh2bIYRkMbfTZxL2Q+59cB5AI3Jp5NQ9/J1ptzH7LeG+3wcQmu2Kr2a77ix7Ot2pOWBGsk
WcWugcE4MB9IBTWadUN2tCjfmU8GxJp1/VBhLfcnsjpnuLNKVytWoRPZ7jvH+g/RiuRDwbVBh4ih
rV29jOnfs6FAZHYkZmENvnNmoZ976mrIUpgKzz35cAOpq4/TJWQqtqhzbVdtLDw56ixzMz84Rupv
2s/1qlx9iQ11KWRnBRUky9Fe+EIHIjh7OCOm2ZAEbxpmDEJPNxT4rS4IWyVjzWHdhiN5n0Ivfm8U
xpR/YegQKm9i7yxX3ERA616dR5S9B6FeRBzH1ogbyqXEAc8G2n9SES7q3n2yZlgGYlkwxbPO+e7q
RVSd6wi7IFoLug5LDssE7wx8z7IBFDPKV5lsPkZ3Tp//n7/G/2GmIWCEE7ljOO0Ns6s/3rzU/n5S
3O0XxErQpDQTj9kgM3XQPMJHVZR4+xTS8zaQnUWMF9JBtVZxH+6hGmhc28gCJDwNnJAdnXuaNEG6
tgRkazSQ2LiFUh6wnRkaCX7fIVYYd33ZKDhygLJxPNyXirEZVmFZBDhN2fY8Of3g8HVwAjoaL/Le
8g3mHvm1pMmhFS6pKWFnS0GcPDZEt7EW9L2G15hWJWbBVjo3hZ0iuEVuvOgBaccT9+hAxrOXHbmn
k5cLG+HyTXdI7pdZ4bkSvb9TZCzPeL6L8xJStulUSL5rQXEI2hTFucZoPWH8JL6uIl1NEO8S6q6B
WHd8lr77znlpu+iqk8F/irNrEy0NOqVT8tG5UKTq9p/3dJaHbSb3YOAfYkM5wEMILXEe5LprBZVB
tiKOSBsjmJwMwSCV3tPb95y0wvlHc2G15AvsEMBwZ8TfvrlhO/JjvHo9a+zCaTLtjAjkGOSmJplo
mCpUYp10nzDX3AN9W5aCCjV15ksz0PY8AdHv+llFMSAFR/53Dkz+6ZGTcst4hMq91+EGhzlhzOcA
uFzW7M3t/y8BtIF9OuystxVqxrc3QZ9So4K5teOJsdqMq24Zhubqg+Jz1WGyUiPd2j0uyHWU5FnK
NyWYRy98ypKKMboM9Fdw+D4LtsrqXWLVX69sIMjHBY6YQyQb0EIT+pmxFJgQwHh1JanZqglL3PVp
4QwIna9ZbfQC4hOKZh5b+F+A1Gwuhju+3I+MDy7sW6Q6Rns7FQ3AghgQZ/ALHDKMCGwAjI5XXbnJ
nF4gFbMdSmRZEHXfKxHGimvw5UFSmC8nYCwCytF2fT1je/zzEQTUVhOUwXOo0BEaFJO4M9hyZXBJ
SCaIvk0OQDgnZlEE2A0r9IgEUtsed6YBk7vxE4U8iO8nDVmqTdfBTjr/JaWKnuLQAWmUqmHbqo81
j6KqO2j+OjjgWS6EueyIcgHMplVX+uB8tFA72/qEP2bKBBPavbskKwg7EJ9bezxl8ATo0V49ofnu
ZUUWQp9i4PpZb1LxjeHZAwslIDDGEMVt/M86NZUWC32caPF6VUV9OJpVwYZQtYDugW+TGwzu6uD5
GK+NaPPIiOzNe8hQKMaPys88ywf0stFLGDuDGZWbws+48D3j7a+d9zS7XibjRDqqtnrYXRec143Q
mBKdX74fQSKhWUC7q4mB4Zw+ZlkY/v9OCrd5zk0IIBpsPKT/gENCGGKDT+l4wYUpYZmfoLWd5dXB
bXzzCz5/zSDMzPJGfqWUiDNcuro8jd80zSgn9mAdnqBRMIjrm27nQUbQZEnu/RNJUJpfdJ2LWQEY
Qu4APydi2mYLbQ97WHY8F235mupm21TgcMW9OHropMAoVWS4jw1EVQNBl9hHvdbkgeVjehEYbOK0
LZ9R6C4Uov/vBGws8bA3w2uqMHN27PzCeg4x2uqdYD4LEuJza298dPF94IVujEeoezUTMnliHWvs
REnaG3XYIeWJsYc3pojpkUdUTiDbGn494SeS6dW3hbNeVdh0Q9XcXmIW3dUR1U8sRHxGrv+KXUZL
/HWKmHvwxVaRVEe8VM+EPsqoam96pxaQZRGh1BDO21EEax3HywFCLrWAmVtMMAe/ERuLfinwGK8y
ocKUmCFS7wuAHJxJ3M3GJtFF4UwoouoTvziE/hcjK6vFY4aSTst4sgcRKYd3rYc5bc70cRE1D5UI
ytUMiIy8atpEgZfRFJ4KpxwpVVdvbfNDAO4it2yurpArMds3cQne82B7Nbk2uknYPsgUSiAFEtil
trFiqUj8+1mC7cUvku9IfOCaV/nG03WhcVADCI29ouPTteHcbPog9Q7nsn8P49gQU+nbdMfMo+ge
sZF0nyaDNjvWw+E2FkXJl7QLtvQm87BjbYM/VLR8oRF0Er1iOVX8dvWZLSWLJei2MZhUOHClL2bi
JDk+Z5MqyvjNTguExm+AkZSPJDkfp5fZ5u6YAB/2/CbxgBfiM9yDyRYw4GIhiwtHcDH0jVMjEtld
NtJGO2ya83K6i100da0cW4VisyazTPCWkMw+9jZiTwg465jukSMjmt4DlerZm7piRWUkPrs1pesV
iEt4sUP/LdwNDAZbxNNOOkN5g+9jxurU6y79HMvwFcGnxjaWdD6Wri4C9inJPdKRmtk1KNiy4CAs
j9/GnU+UwtTSRgBOeU+YZ/r9FOkxt/gclT+ChXxwyXtXmgqN2kTrPkTGUHuXp0XOwn2FIcOgyBi5
95czBTY0llxV85BOhf5TDLcsZSmZAAN3TfreUhJiSIW2TzzNR5NURKk2vZtWtS2IgpVAmVI6alO5
NTPxpD8NGYh+SxS2pJVq1lZHQQS50w0XyXaB4dKZIAEBV9Rv9LclW+ycfKJdfYXJE4cPAzMXn8X4
hxMJdWZncncZxI92uaF7ZJHxF9Lsu7KK0O6lBKHLUbHnj5mrjJBgnneTRP1eueBy6gbvMB1P3EUU
QBYVfs3gmGn9oZuYlKTIdMLjBieqvZD0ses0KDLkJ93LMYnGeHEj1ArMYPL2Oe7rKW1MxhP2ztBd
itf5HMzbLeAV2w/JbAQ4Zh1pKQCSJ09pkcWcmcnUhriux0AQbaGKH9eYkNCsHr11VxawxCfNYHoC
yE7+NXyjQ4SoHPLVkMRr6e6xWPMigQ5J+ZhlHTRGO9qp2gmDvNfy00YzrzOuiv65djcJSc4KNaH7
rLLsvzfoKCZOwFryXj+/X3AbSXGC45toV1FRtN9h5E4tg3JlonGBPg1XEgSsO/aB042GBz51NVgY
EEZ5QRSy1vRzjel677uLOhd4CiQeeH11uJUoHT/ysFy7OIRr++nK94WFt5qk3WlxVr45gHA37z4h
WqIyhazkOx4T+V5PG9ONW9xhBLe17I4rkW1WwEVVoivTIuxUYq43lOc7HoV5Q2Zs4LlGG6tmUIqR
1xKPKq9ukUIdbW/jIFr3+bmOO+RvSD6E7DrNNOWzYvIvzJyiJy3oBJnRAxHOU8CBoY/ahGBQ92wi
qF7WcerVfqX0+RKADlBr0HluaMDNslJQb94+bGcUDlO66I1iDPc+yV61xtwdGJQcC4UOOiGDqJ4R
7pDFiijYbGe8/rM9fK6N0fkQfsRh3vhJpcqKRmCAHtoSBEcAUrwhi3qThw1VMzhFb3gx1hlS+Kln
0ST/gKOE41vucyzEsN/1xJZZDCAm1TgU3Ix2T4OrDctpgHPrYsZJyWjM2GNfNqEsG6e/Bmk8ho//
PTvKbrW15JnCvoDqsfIv9KH+hvxjM1QnG3Ua5zHrfyAxxyDfZ5tnNieQwRm20iterSkUc1XyM5jj
dtXKqc5OQHvSIA3VIE+7Ive0aLXogdeWUzNOY/uey6eZvtxxa0ilc4MUi66+zxojC5sbjU/szOHu
pZhRf9Y5eoT15yy3+DdWiKGpWPemuERq553cYY8QxsyBteb0RbEQZhLU80gif6qOwBYFC8e4vlLc
eFaPhB5V+OTehWs1P3HgWkEyMOylFrrptTDlOntzBPlWg5WrSWZqUDjHfIKae5JldTNBNO+VfaKv
1u45A+c62PDZ1QZKFA9I3/tyDr9Vy3k4hC4le1qVK2LrPbQSZmH250iWOsLigU0vcIMCyhy+clnd
G1BXSAtcU1AbEWCSSWiYMbL8wVFyxFphnLTuqddslSaHT509LiVNPFWlUcw7SyIwkbcKZgTqIvrx
B9TZ1nZyFaH/sKT7h6B5TXj4JuVVqPSPY21FQSvaUEBn1/TEPSSzckJSVJQJpqUwRe5HWO287azu
BqauPhDb8Ikc9Ybd413wCbw0ezk3qRjBOXuUSsA1fbnMO6sb5sVHnz03NUb8lhIhCkyq4Qkyrmp1
xmg4k3s0A/MCnj9E10/5Wcl8rfK4MbHRkBaxHFnJ22voPb4GhlIDz3oropyKZ51ps1ruvrnhXDqp
LZYwsx+alIo6J132Wso8izjYJNCaYGmZ+qNpMVK2dzBfMh7ahpWU9aINbe7MHxhjmdvxKAyVjZ2q
ocC83JJpLiAG5jgLIiaUHPiX4R5NLc6V+qSSF5GOixdg+7yXxNmOAQPMTNmU4r4sY/BCw2TcVluz
m6IH9zgJQcjOUfpNnijmjFa0+E8N303pV70fMh95wmVokXt4e+wgu3TWVINuexI2FphpDwSvf/iw
Kwg7aD5mkP6gVEf9/uct9VQ7IIUOUxPdDlECZ3DrbC25+VvTfMBNdCRf/2b7l/fkjA2wKADDI7DN
g/u5bxOgnjCcAMxVlKhb7sedQLi6xnVM33YnpW+K1IrrOQfoAabpU/sxozgZ3iYiLJGzqcB+r9VJ
brvgesRQ3R4quh8G+edYiuGvHo8DhB7FR1ki9nG8rQAR5t6SVV/sQAAjMjT3KVvBLkV4N6b6dQw8
cIUQZgxQ8ksbnCNJkzgXNbmBsMO/RTxZBupV8sYad6PHUVNwBGQ3zo9JEDNPDCzt5NduxqV66vpw
RN5i9rtyPBwY4ZR3LfI3i/aKMLFquZoVrxleV0lopsrFlznERWCFej3MrnzfbNf3zYv8hF3/Sg3I
h6cL9je+/KWTPp2U3PMgoFCtFeE2W40dIWiFwxKuKKP8XBSa4bsUUwhLSYnuMw26LB0nif/RiTmo
wRIPSx2epHGXivoDevnnEiSgvnScW+opBMPMOIWHDMcUA43mMTCshNSUdOgyhfqUGFKnJorDqceS
Z2Yftt5XcsrsTMaArRFh8WZWLFZ+Qe/+qxsqFCGz81Kz+BDlaovZrej9IaqHHOFw9a7MLJpw/sX8
dpx1kRR2LMZk2R75aJuAO6S1/K68170FoQnGib/N5JS4rK1avpMXXXfv6zbfgWVgZglqxR66hi9E
0ku/r6McLL1U5zQuBhLONmosK09CGYWo0747nwRINQmXOsJ7tQmAFripQ72zlGRn0IUKy4fnoVdJ
PAK2Qv82gvK10KAOB/UsIFIBdqkHcYIwoyo9nuQazX7Sb+2YJXxLKrsw/MuncT7eX+srsQ07e1MZ
aaEnGBk81WGBre+AIvU0UoxwyJwGSqBpvX8OY4y6uj+BWY24uWZyio1gXUHrtrenetRBHpXeH+Wd
s4KiHqe58Bzh+W7Xlpy2aICjzBF+F/UDBCyBI8FXZTVr2KbNEJ9HVp13NRlCL23xUxq2BJwjejGM
nOipuqQ//SuGRDyNaAJtUR6F4pU1etH/Htmo5vhQCbyzkjDcLDO/KeZcY8zSVX+BpBKpqcWkjgFr
Y/3rO9fTN1Eq+z5iWSV6iM5pMC2+6Y2u6tzcJJwmVtKXyCOpfS3pfxCnQSerBai0ZUWDZytxihrF
gAnS5MsL7Pq+ZnCOMxWBHvuD2gL7nIe7YlmWeXnDJMgxKWl7lWmZNKrCO5e9tuxYoNP0mumAcs4O
AHh8BiC2reeyn0DH6QTiZAWiBACRRIWJgyuaQLdXF1ulvQhlzgcMrGvrUopFBwD6NfIK6Nq0C928
GQdt8wB20gV34JQnX/E9N2g4sK6B5rn2VQ4b+Z+l9nXxBVsFsx9uu9ld67kj4d1VaOzEnLmw2VdT
UQzxleXJnOtqhwP8F8bTT+foB2G+iffZwA3p/3QZcaYup6NI1NPzfbJ1PAVKnk68osKsSsUUs6aZ
IFlKbpejYJ0oq++ViNodJdYMtYu1ttSf+cNuaCdpT5yy+zhy61uk00JsCL42jZHQTrAqO/XZlrz8
w9cwxxnmauGumdBnMDYBSrAoGbQMDIE6IP35S28T9kVhi4HTusQsRXPsrrzbHtHebtg/aAZM3uwK
H+bt391sXaKxCyQWf7Gz6H/bU1fZXAF6C2vWvZcZdzPir3ByC6csD/foQCefZPNSODmYaXNYw2Gb
VMxOrP2XMyfvUSpTaYeAmZA56ZKgbqDYysdO2vOvmTjIu/J97w9aukmxZAjPGPQpdHWCSyxp4dwL
vwmLF/+/sAce/jr/PLtEB6mtQRQwYlrZoVOGj1pmqVp3zS6aCO0rhqFB22y4kqx/scEGknAUTJS9
UyCY4l2KT4FiOde1sGPo79P/V5sUO6LuRIhOixIlsG9/4yYuxTInQ5AT4GWUngZm4Mso7LdNLFbq
DqGi1TDEGCQa6HE4GdzivPJ2qjH0Grt4gODhW+pUP1Rqin5vYTo+0/CIsmwqjKDWnWFjDJf3MnWh
QhAT0Jk4DFCrjkuCi5LKugVfWw87HVsS/9Y4DlYIvRiagB0blE3lF5FJhwJDYofRz3d0jtrSRAac
DPmJkxvK0A/d6nfReuc0wZUsx2/e5J2MtcirL990HydsAoA9JJG8XtbAudnz6zjMgeiiUAFrCfIm
iOfcwQlSdZ7XComwY20zueg1QQyKUd6gyaAP0tj2S0Iua5a/zhaWS/T0YxFn3WI1+UYMmzqRiQz1
nkr4HO14xGi2qHKXLfsLbBXshjM0cKt9BT1280+Hq4T3w1NaWXnoUaJdzXiIOpgzVRQIyXaQrkPZ
/a37MfDKR3ZQTevqAW2t0sOR3NnfXdubnJbrcKUkVhxUG/28itAgHxXzhvxzqqnVQvXBPaA3iLSv
YceJQDaILOYGJwfpneyUOCdW3kP7sk1AQDOgENd8PR8wLvcu7+OnF33Opa+1A2+8o9U+0IPcj0fA
KTRGEPCLho59j6ki2DEabMLairo9MBUug1ip9GqPOK7+T6bowUj20a3qt/W3VhBlprjDIKaHPdWu
IsCtNOiI0hTSL69iJa6f3hbtMwmYsdfCWMHsmUiw0uAdsBC2GICZRmnHm7OfRQ1dK0IkJF4qDjHw
uLfil6yAYUiZ8v0SlaEYLvXXmcEFdxYxU4yl0Lhufjvchy9lSRiI6vLSxvPxIxl3TUBvwASs2LUQ
ueeovu4nqpnIEed6ng14l/v9X3qRjilP3mUNnONkkoaB0VHxMKmgSK1dwzYZ/JBFNPkVHwBOELIn
LNd2nWrpJx6KxA9I/vUT3tpAiLWtjO0HZa0bdLvJWIjxv5jPTRHGt0Iz/36Q46VOuHd53XcECXjZ
5ydE6VR69WDeHQ011QJvjeMEWmosvdX5fHyyDTcemSn/s9a9MM/4hcx5P/vbyjSqKVmD/tJSxbGW
dXSop860MQqZMcG7Obvr0d53IdG87Yc+OdijHaQjUW3wCTMNYJecR9x6+3lTxPoGx002HV9Zpj1d
piO34KD5+xFKDST/jPQiQVIZ+KCKXPqko+seHgQ5dl+e1zInYTvCwRfUbHhjPo/3voAsK/NUREkm
64diKYptXSPlsjDartKiZd5+RFojuwdYJjPDSWkvmedadqtXJ6blFV3YnJsPDyVkwRVW8EPlufal
bdgyz0G4IJ1mmwI9+qr1alwMrvTQa6xFAZ0UOUntnefpHB0PvQ1kvKOiZWDqNSfwW2zg05b3wR8e
AnUfljWKVrACx9pA3J23xvtCu2gRNv2Ov6gd0/5Ci8AVqmew4zpcb2wq+EArpNis6GinPB9HgBuR
KlyeyuZLL9rlW0zASmlpcxlSxoDDTZ7II/BSI8bX5LyUCpkxgIw+3xvWgGbGkHzDcrRuVLWgQujw
K8loyxDUCsx9Ggn+4qjd1RVRf59nXqFye7BRPmZjbqRBu65atQ4Eu8xs+m6gxq+LsbpUcdR8Jffl
Axs+U8sur7VyKwB3VtG0cRI9j0VTtsNS0RTrVFbcrUDacb/5lfgRcAxMOcnyTngHfFVQJc6/mLYB
l1BKisrB15ZqQ09ILCjqi7nWlvjWgziMgFbCQ5fpghrHELlKuW55M/I9A/5CoMccIpkb696W7nCB
tpw7EodY3V9hWhnbh6mSliD6MkgrVn6Yxa9tKAQ3vA1BbZhNncDGc07S61vSeA6bM9Y6iBaSI3Jt
E2OZq8FPvGYFtlF886p1tpTW0bRF9r4+S4G9sFs5xCYPJMosW+7uFm03DUJSdz8pegeHOhEHEZ/X
Huuat0IG9BdZf+8njk3af6F+hUO3yT+pmcbm2jT6drlDd+Nq6lPRHj5V31OLo9ATwlFSwCqfkrqR
UPAbgOp1BDdfAaNL9yl3QyY9FT4I4bHCrQTIFzn1rpOY/rrRr3JA+Bze/oKXgA3b8oMCpr0ITaN+
kDWLVBa52nmSBM7MkoGMsfhp1Gx8zDU5yy7r2AhpFtESF98uplPsipHmidaU85gXZaTlEWQUro9S
dq6ud1j0HBbkjp8Nb2yAdAmqLFS1mqhrJD/h7J5BpCRPhmIqdKzuP4wH0vi+maSNM6eJG5LksJXA
CJlKe6oz15GSbOCd/hZQhpV+UQ/KGHRkCyasu5uG7JisN52PtSeE0P/Nj+SRvuShCeoqNV8V2lSf
NAEJQtJthN8gZkXDD2TsqpNMAjcMkBwj1mTYabW9+VPnnEeB7dc2igwedA/8vOuM5MQmnM73x3/l
jVIGkRL+0Abm9qti52Xrm11+tS/aVtpxofEn+8iO5c5VhaRcqjxa0HrqgRnUuNPUnBWFFdAkdAtb
lPF7zyvJFdCeDJ0ZAx0ELtqQNk7vCNSzGQFXci/5RoY+BStQ+sr4tPAjFkdma0EdG3IZmAkVAlwB
C+1axPhFQtBDoumGNcrJG1Z6oMzV5TukNYesrKY+TLQyyT9ELoXEP6AEblfBPmsxnQxoSnmzJ8bc
P0TPtUKgfK0wusYVvgbtfpE9oD1nwc/MCc10vt2KVQxJMKm56S69OEs6goTpARJ6PbVDP74UikcR
+kCJCOtJbNEeMJV/scTwKwzCi+qU3LM/oPJFf6bZIYJ2QoqTFnX6bN4UVcHrcb5oG/0jNip9EjBz
m75w6/A2CeAXRuKxTQDbWoNgy5JonzRjPfoZ1uroS1VM9rE5kJ9vNCPOhIO7ynQfXrELsEYWiCRi
ENtlJhkhFhU8YCZB0EbClQpwjsgJeg6jBxMzTskIorP7w5ux36slol8SwX8PMOvbZ/Q23gS4iYZZ
6Jp2cIQzi2hHIYw+H90q+txTo0EFdk0Lzhj6/Ul4iUodwzV+EGxsSALqQL/0AdBs1+GGUJzqmz+/
fi7QLKuJ6JKNwr19Zzuev/cy2/fny3uMuoa+vYBCVnmA/zju8w2lIfF5GF6l1uw/KjiThWjwesCf
F6D+RNjAKrGSdJmWOGR7AiRBTMM0oCP4Dbi7DOz0ghCW9fLR36fvpjqmi8tOS0zbRJ3mdhpfVk82
cvww4Y5xOzvNaMeQrj8D2I+8tOJrWTyIaiLjZ0Mz47lMcMjkzHPQ0E1fab7mCVLV3wrcLXuFVmKk
dBURlf/onh4Gbb5suE+iJtIGo56GLQzp5jdL/yU/ixX4EPuhMwop8OLTKGMlP3QrLZPppfwlszJR
fP4QSpFTJsJSExKh/OazQTSQsgTniMb+2LNESXLKuUJL3sJgICmB5HIS0FymuL2HnoDQFIr31prt
PqMceROGlhahpCYw7lFvt1nhY8iYK27T5mH5RS162Kuw2G1K0033SKlJRGFYsILYxQV99hPqATse
4R83pOBba+3vBECPqZunI/TWESGSVgpFQeblNI3eizb37uLc4dgYH9ZIgkPQvKn4WL1A3hNk2k30
/PvIRgINOtb/3gwqd6foowqtsHG//vqQaJI9Xr33qReyMeMFq9GglUqVOu6xZT9S6eQURr4BfFtx
Ii0QjnJUWKqNWvfkyOmohCuVcgrT98iDroXwILtLKLxjA/7QPeRgLIomItfe8HMpENnQiHJl8Hdq
7DxM1lxpYSrizwNlzp/Q34/r9/sdSb6zA2qNUabLZeGJrsI1LDvDsE7J3HDjJdeO0ffqakJE9kdr
3uyCF4Ym6fFWluMg3S+XujgoiqQHqXFJSUVVkMJRQGYrBPcnXqK+clTFa+Yu99uQzmsbQY+ehj6R
Rl+f9Tl0JOTxCaJZzrmDuFAe/ZTv85n2K93xZ38o8vw+hZoqwUcwwy8sKyyLDs0AH+ENBtLjuiW0
WjGYYpEfu2qG0UX7/BaYvAH6OMVy2sQElJXQCN6rZtADz9R87XZ9CdcrwehVk/5w4+z+zQFZeGGx
CzZv33/Z8KkRpgm6qQ3lFlcD9Hw7t2U1iv2/CPGvkx/B1mz9cFBRa1Zp4WkhDRtxuqCODMyOOhSb
DREmYOGGrnGVFq9FLv2K1UzQyhKYWL70JoYGiw6Y7gqQqp3djd/dJqwIiQ2Bq5cx7JUw8OrGJb1E
349YE6QXx6e58ku0EnTUUVIp8ZTDuYhDX230o1Ta7FHbY45KzHj3J4wV2sGOWVA1wLoc+vBSSByT
IMeG4/Xeb7o4hW6UEETrTryl5jNJ5zI7M96Eu4UpSGip0eUaJ1iC5B8+5bwiApkVzdLRz0L6sQeF
O2BcD0eczFAPSEryrul3TgD1ZZ3fgFG+Vj+yst5YYG1PwAQgDVdnMu8NEmvtR8lL7mzH2MdRCb44
F1fdUvS6xnQGvvjteQDnRtlVaWmZ+GawtJ9EX//VHTEOHjeNOVyzbhbSBYAga+2xWwKo5Y1lkbYW
XCfNirOaR0/OTQiEU6q5/17KliuWPQQbpxv9do122VQch7i6aRtZ49ECPrXZxFgXIIe5b5PTqeT7
8B6Mh7VvvN33RVqwuFpZyZ07fTodmdCamsLXZ0Bs4xKwVzBge0fx5XBa423rwzcuVmre6AfLAWAS
FQs9/UfSJqJr+DSVTcj5gabLUAfeMgYmWm7Ts90sxhMTE5vC73oipsN1IbEE5nxEVlDeerdcyYQ/
jIGzhTqpNy7YfkHyBkO+Qq+KXncp7+46uAJSLhUfkWQYmCgtVJzmhkjGbxwUJcgakvXM8oN0G3xd
oZ2hIojsCA8UHLiAp2lsoEeT8W38Y0Vd7AI6rrbNH7/D1xwylqYIU68K8Rb+WuK6H10JUWPprGSv
OTRcVrEgWklqrhejEQxKQ9DU/XgpzBhj5Pk+PBYP/2cwATtZRtVKZsyDLbDp5l7dO7Gq1tD7B4lw
TH1BiTB6x0L/SUbxcYPS+/khhTeHwizyzQlhGRkpJPCGr6+wXE4BOFhxsJsf+bftmwW74d4cTeqJ
vRngvjmWRSRcYB+64z+dGNAiFDuIdHsz2vm5oCd+LaEks1DKW+y52ng51uuNuevtJm3oB7Qj8RT7
0S9EBeUB1vtxg1ePNKvn5Irb30TttVc5zEqaq5bQdL27mRoL7MUVFczBXLfy3JU4RvjnFHKt5aZh
6RNjgSglZYQJTMItw9uI5pDRScSgF91Gy0KWtdzcEuR3uwwh398Btk79KROZ+a3qVTCXK2EHVoYI
Au2UpqGeBezpzq3SoSU8vxdh+7JotGf5hqmElCBRa+dDanxvDL0j0tfuW4V+G1JeBqCTT/KLjHAm
KNiRgRIFUKPWL9Ud3I3UqnuA/OJU76WoH1XrfEHs3Iw2KfDD2sW7Qdl/O3/qRMAE8FKcQqG/3xER
9drxQp1+pCYSJkyK0cfj+SHuNAgHPpPHz/1m7u/9w5nkBGbfAl9JoIB9HvzE9aZuHptiNGbdB3iI
oPTe2JKEeJpL15i4Hg7BFjlfmJCOWPMrYOfEy6YPSr/u/mlJBqjOb0Y2rd+pHc+4zyhyg+F+0J4j
i17Hr2qqJXMkC4QXoTjaMofNBDuBrXz/7zPRz6FUzncDGu/iD+mcM6WvzMLDMk2gLpHk9mOtWkuU
uYoVEp8gq2VZdaSN4vKilDDIrjO2QsmyvRFvl4zq//RVqgjfTMeSNxTIQZDLyaC/lLFUTY8XTXFd
ANgXu+K9aMvjKbQdOVl6qeVkI+NkqWacM+YnYCSkXHYLoRWgR+fxxSl4amm/xGr49SXmUPShGcxe
5pTixBmwqth+ycQaqHcG+x4dVMJYKZDJIVVIkp9iH0I09kKuy0QqkdEB1lVRKLJ81We9Ce7m3xj3
WvyIcO4rruipwRVn2IdQermjr7gEjEwnTthlAvIY8D2BoFqJN5ijvd27SYLq6hf+Vb84WpZ+3eBr
lfC+9rabJURb/MKLqwmnOi3G+oq1okOy5AapHAqjJ7nDYZfkhfyOmZTjZU5jDqbjGivNWJ8ZXl+T
JbsqHSA7vGd6DLeVkP9drf0IyOglxcfA9hDDZDyK0pLPUfIFq5OQWpkQLTW0iwpbNx65mXxOcgmv
PY6b/FDLuO7R1NBAuQut82E3MKsRF+JhPkP2fHi4YGDtZtsztthNssJPjX6tXTnxJDqSbgzxDh9I
5G4ao+OfCEMrg89yZ8epFojfWlnFxyDvK4KGOiZzTk1oFToPxti1/6Z7nAiFVNk16+fXQNj+aySw
TY1Gmb3sqpkgF9AtwubGqLocKR5A4PFsMLbHpwu+7O8ZMybPq8DN07htFe4gfOQkcF9v0hWc19V8
QR2cGaJmSp0cGvrgJXLgOsFHrTB839hvFa9RIvnfn5pgTD+iPF7kqgw+FrVetU3Vq+RclRTBKE9L
YbLUzCxPwGRQbNIXSgS5ai8Siz+aGvz9VJ+nXUNwj70t3HGT+E1OMvqr8dth4F2IyzF6YlcbYp5Y
cvNdwMbcRLIC9ovv17MQbSM+JXM/asC+8G51c4gE+VP5yPaZ8fEFT8hvXUsmj6gekaNZhnQ/jtgW
Gox0OE7VEtyp+O1sWUxVPQt6cgo+p+1ftASs2dSb9SwCikAgFGRF4GpkWmxg7aplxL3MMhPlQ0ES
5eZxZAP6S9lzedifMAsNnO1GrIcE7BoON3ixbIYtInWyqPbEy5bbp04q1YRlOR3PH1jkVmb3NQ/u
W3INqOiklasgl4lwyldG2dj2lDO4+OTWa9Ud784Ae64/Dq8A/Gix751N0hrgWukXe3dQX8p2pliM
Vst+TxRPiw9Cs+hXBS8jsESWEqv2GuNqTXQu0iLVQPopH24vBCqcmfsZgoWeIq7R7acvEdBHSAB6
4fl99mbdg9W3mv/XXSVF/mfLKMGz1HlY1iCjAru6cd2ykTmZu/iNMSinCgRE0SLv0ubbTa+2RTqw
uosx5zZlNUITipY9CK/8hnc1kUqYnIZaD5pCFPh/d6gfQXOd/utXGgL4mAJmOLMk/JT1NOyYkgpi
wA1T/1QbLL7Ya5vaD8elbrVMqT++6I8hrQToT1dmAcIDFh+X5oI787RQHoIOC9LjVN2kfNGGtpcI
BMvK2fRtB5pI4LgM8WnrCIaRiRtQXIsSjyRAWUAxxvCQ/BJHJJSvc3c9D5OKzNUUGsd6Hvmq5zif
g0NTHGCoFZDZLSsjOkaO3eV3qEIh9VEnelQYHxSmvO9dvwwVCg30AieARFEpNpe5Jp1UFOMshCrx
tidG2zng3GHFtdSs0XJLSy9aCsd4DNmPXpAS2AFsCZYaSb5bNZrZ2Aq1OF937zuEWu2+HOQOfmjG
F2DlqUj1k79pokMCtMGBnyZDe5eBZsFkuGLByU0H+R/6tJPLYHGkwaE/Z9k3agDq7YSLw/LNNn1M
lGuphcmNR7aMK9jy0YJkRHq3yrofGB2cVHalzzD/Ozwde3rC8VWAM56yGLm5tqkj7B+ZOha0++h+
+p7N6BkJncSbKNIU5bkdB7bEozfbu14GUZoWvXqVAEukODI1CzIGHm6la84t5WWjvqT8tx8x2XE4
ktqhz/KQOFSY2u22AtGFc4RCGphcwqxr1w5FS1ThCwkEfVQitMKe56ym4ikDujFU71O/g5H3qrWP
050bG9Bf3qfisA1mhfGYk8VSogyZAO4pAB16CvyOkUEMKCPwL8OpZhdXPXOJrNjB3BcSaw00UYYZ
NQ8ISgojs+hmD4zwHZim48ybaatJEx/vUxOKVx6Yayfh9PhmbxV6WnrMZ2ASJFR6If+LEtHvHUu3
47L1xSMrnzqqKytDdsGBz8USi2IOUlhvOMhtK51ZW+eUZ6ULFChgY7MWbcMwx4llDYvn7PQ+KqKA
JLNdmK3MFLpmqC3dCqiRrkruNNwdTztgV9gOfBu1N1IVwQ60cCzkU9qj9WDg9ywSFM4xZr7+ROWQ
24mGswKhWFQ8KISuH05X4coCr7CY9iTxtzl7udVGW2rNKckzKhd6jwKqzd68vfKMyTNgm48fqdtE
NKuhlAU4+TS6uHIbwyLsAj1V9xia9dT0FaTy2Lr91QzER0EThbM23kL2dvLetSt9qZnXoDREsF/h
mO6R2AVKLgVBrfESeaOo2V8lOox7dE1GVSlAR1Ak4gYq6UAmiZ5hLgijmmRuhKNTqtS8g3w55XUy
BCobYBwfPkLt8y1WIZuD/pBPV+N8R2kpaiJKK7bSG18ziGaX3ORaffmRf8z+2THBkOFcfRFOYv5w
W/q7CP1TgRW3smdFbHQ7kycTuQ2hBOPjH5s5qCNATQ2Y2hBobvu2oEUrIH2x7SnIP8iyqV+IqlFB
pnYsAYXxc38S44Lae2zJTeMmR+kV3uX0bHIofs67Kp0At68+hlsrQqNf1M5xz3VSxlKv1b8QkF86
PN3fLw6GfakUQQ8lp5hV/uZmjVxRuox9/lLtXa8rm9tYHTCu14Grs2f54J41OLM7ylnUTY+7hVj0
ZG6JhiEBpo2URlDoVbxLluhzIUghGjXanqMWFA2y9cp3pMIWDasuBryZffdqtPNewoX53hv21Npq
K2XBbEhjtiYH+1mbo0ScjW6GDqU4FpAqN52ZkPJXDeuF4erQNY7/JRDJoDBrx1RSyvugzt1xwp0z
zvxtylEuXwLf1W5d6oYOA4CpfjV7l4FZALOy1WxaMBYlLdVmkEz5M5cAqeJq74ilHuoDpkTkwF+h
WjxU0G40tfpNP9BzjjFqG1jmaAoKvdiFeS+ktDEWRg2//FhHF1aihPfNjDRh/k2CKrGodlCzILuW
+BaStw1ra8LmTZPgJK2c8FFz4Dl8ladnfJbuudBjCKHC5icePrzRQaBySGzE3lN1NX1TacFBRAP7
3hrNRrfMxHo06yjVD/95zEWFTIiXb3Rx2RjnFX1V8UTTvDEJhepinB3Vdwwfz2KJxPLQ2J1Pk3DM
ige+iNQqj9Gy2+JH7/ZU+DsWS8f7H0byil362yrSett0Iv0Arx3926StPgZBM0YP2rMOGysy3qcO
bfnsYJoYCP8YP2bcYIjr/d2VOaTXRlMUgqQHeFUPg05nuReT8IgQz3kDy1R+uMt6GC3O8U7mlp8S
iWehZr0OBpYhjr9wcTMIzMWtyymsCcvVFxUrtfBaTq6LVlByt0yVy2nwrgOwLcgMEK3tVrfWHPlK
u+fVp9mbf3Xl1dAppSZTG8Wbyr4Mu5rZUDUnNa0NDspFcj50u0I+C+jdFobunOmtEeABC+upJx7b
vaBtgvdUk/3ugXMZ5MW0x1QcHoJFM+XY6Y2Y7t0/vaPXLwJhGJhy4kTolvqESTzZx+WcdLP/b/Ld
LwnKy5HMMW0zC7zB0Tz1qlLqavKLk727XYlq0rkPC6++tPjBl+miTIz7V/rjRT49i1MFYkRs1j5a
t7+ghomdQPGfC86BordoR0r7ZYX4gKtyIZ+ec/F+Q/jH1LfsJerBObwsfJKs4bGi/T4YPHL4YUys
6fXAiq38sdAtCKS+au1SxzY0OoAwA2W+xBfdP4M+WOIYzc4nE1M8qwjldR8/bwP77hh7xon6w/aU
6XG/PWqYWRJWuhdEhFpHX+5C4J7GovUGzfWy2ryZ7xIanoBhL4TZz1FXTdBMjtrtfVjYtSPfie/q
8LeP0jDb58gqlufEUA/Hr7Z88QqM6r/FEn1lTmNFD0wLxsDxDdfYjctpcjb8UxFCw1+wUX5ZWo84
GH9VBsmwJX5xZBfJm01/uxvAN7ehlOK5fbNRYgaAWZQSfOrlRJ73DJF66dsj6KXHC4r67cgIrLNs
CWIq1owReliJ7JlEkvJ0d7mC/oXsDb/IxoXqAXJx+1kjkel1m3QFOW0Wt+iY3AW69X2aZw9B+QaT
+n4E8o59BlvhdoBn91yoePLWConEDHmmmEdLxoPhzxnSWKqmEQV/QpsQzaDtHa8aqz3wkfGOUfEN
33LSIk4GgTduYjRy+FyTfxdC9HwZyJ31S+g+XObzf5nBbZOirwrYBktgBeIH4yiJx+2KEGyimA0P
0PVXd+u7WSubE2Sz3Pauh5Mslwh1RDyMMtkHRzmGiJLjBrDgnKo7rUhMcc7BJvEvribFHTFuveAj
LDuyL6/v+tv9FehjfTWyQ98f4yuVx7vrdBLpMfhrfOEXU8h7upciTFA5/02VhWq5VFPHncH2v5uH
yQVMgisRa5lr5Gx8DurSFG1qIFtJUIyfi+wu+v7gB953GtexC+hRQBQpvwrxMsPWh4ClrmmSlQQj
cGlSPYYC00PP/bzthiufmaCMpp9eW7IT/yfLgG2XLyOglZ1KKppfwDPT38jkvPDevFSij5eng0T5
hxDDHvCh3dyKFe7m8eQiXmwf4Fvh7RAf/Gt1ffOK+c5Vs3CpSPcHp+AtLbpqxCye1LE7BRFgMG/J
1YIwlLnaHY3ZMWGcT/2OvP+mLDLWE7B3/B2eIzjJdIOmJ5w3GEcRzo7QmGBaA/8Z4RDRFJ333ZEe
QNRm33SA6MXuoYw9dbuukmPJrCmFbWh7d+QM/Jo6eRf40SSUe0sFCghkFebNryeU+swgGB06Nf3o
HDuPOl3t0xJb/SNOHFdROnyRoNKrpPrsA4S0UWq6WQb7KLDWIETfDAKdyhY4Zgn+sgw82cioQrUt
greQckXsG5V9t5ClzzyRsWKePnaLlW798b6sRsAhOkiX/q9OmZB2I7Nw9ro8DvXMFnNSZxjyJDE3
BKjtIC+1aoO3QdDKckejXP/634iqbDU+tr1ax1Tk3u+1bkywnAsThPErkBBySPOlH5lTmNViHBHi
gdYCyBABI6cOWzaZzmaPlMbRYRmJsdSjpoZhsuarBSG+iOflfgNQEJ4J9zP1wHaRflxrf1EtIMMF
YcvA3TBj4dnE3F36XQbp8fqaG6kfKDtByDpomVhV4krbsOQdxXtyYBJd8n2hrS6krhMeivfRw5rS
aOpYhZxGDCclgYQE5jqRzgfK7PTCxo3vZprhwfWfMj88GhKQUTwdGUBrV0QplSYCmk9LtOzriJiZ
X+qS0lQtb3WFG8d5HtpgLnWdgLq+Ea/cWhI+jqzcTe2BTD0bCBF74uV7mVy82CN5s49nwUWhUlV2
EIVsmQKADLIm6wC5apj1rUM3an/04DijopLBw7NgLOMYUyfu0IZ2tsSgpFvVtiwalf4dXikZnHSd
ObRIvSa/4Np5Lasl5niYAMMD14iFaMrOwKQ3IF3qAvjPqxk5Fmq4XWBwSxOLGPtSoJF55XQM6gAv
GlpPLcuunOBBqCC5tBWWgihuBw0PFxKDT/xFhgyDuBJJwl06cEhnqVE5xnivL4tHAHPAOsBSBxgp
hJpFXp+RxoqNphSkbl6rc9nalVNu5Gg38tUkrSaHYpr4uYq8zZ0L1iHxZlVD9Ci/ADxIInZ1m4mz
JmigFz5aUBXxmWClqRZ7mWVXQNLxP1QYU3kr3vsHHuYYjTf0HLwyi3ewOQF3HdnEYYKfXULnZiuc
tA2PIgX6Av7hP9Lr/4K0ebSxEZ96AwMJRMyhxsO6rxAmQ3MncXSZMc80Xk1h1UL4Wg7fgz5Gh+LD
9F3nh9psXOFUAttmcDbSa3VqWwp0ic5YTqlquut6Sb1ObbDSfJB9eSSFT/FvMFy6S9fOcyaYtdqn
C3qFxbDzsQFEhvWlJVemxrsXbWg6LQ5G1WSLFxD3UGHxzw8w6jSP9nFK72FCofdQwgp0EC3SW7Y7
jEhOkCpGOx5REw3dwsK/l5Xy7Y2UIFrKMub6ZhY0IOBupDyPI91xQ45IJOv+f3sWbVwHpRCyC8eV
TBxoCKCXs3dAUVPNJos/fkX80xY2xs7r/+CFCZ42H8WWo9k1TTV6p0yaknhHQPrLoSr1H0nFgHsA
zFGSj+hUsgPef39NMulYszkWkStmq2EW3kUQhCvNZUbb/p1FGlS38o86R17VTq7UiPSEgr9bCEgO
oi2LDd9/uy54Hom6jRQrra1Mbtp8sdoZl71DufSZYudQ4xozW1TNjWz2g9lZsQ0NSOYOqrfa4Xyw
TQYPiNIO7uU9vp/rkHddIwotpoFOs7RnGqnnfcW2LUmYMu2bGgP3g+0RpRGMi7eNg1/QLM5HV3AV
NgHbOIVHO7P+HigIL25/9vR7lw2kcT/XHtcRA9G3kL2DyiS2WmAPHZpRb041RZetDScEdkoyaSHi
mMnHUIUbQPi9sp5vyjor+hTKcbJxqdofF76yOj9GPtSb5FsDGhCbEPFuztx6qpbWb3EltqajE1GF
vTapOl8IrOuT7Xveh1s8gwNF4kCJQOrRnYKHbJIK3F9FnUiAuTMFoA9rcMdgcgLmHUisGsn+Y7hJ
Fo9PMZTQzX5MY3S/RhGi5bNwdcDujdtPqHDhi7dNUTHTCl+iu9rVMsaOCwqq/KK1sJj1dbL5QrzY
pCHZUAo411TUqnk4z1jo5+pOD7O8h4XAQPifkFR1fPJBodYc5yHnlRGsqkujajfEJbvIpeirJQgY
iT6MPpf6JzrCvv5xYUQZi0W+VkQBWAhg5Om2kh08OiEld9ivLcfPad4o14ExDWcLQNr1kBZC3ERg
U4bZTgEO19TKHukUzBXXUWL86kT+TQx2/vYO+TRpXK8ljZlwxrRJUpbL3QaPEtwJjBjHDyK9eyVJ
sZSYkt1kVwOOW39CyOrpFZqnhkB71iPvi2oV+V33eFXSwH8++RAtstmPl1NCaQ0ClnuooGeGy/X7
T3xubQbgi7X7RLghoeJlqGPBOzVLtUlqY12pmVqJHBv4+HE2QGX86xR2TJH+0e4bBUGV6cy1nGTh
iG3lOnUOYhA7veLa9ZpB2rOGXW9Ywx9yGEtkXeBydz7Gb62pEBdfBZ3CFVID4kwKkMkMUeSvT+Nu
ehcMB9HWZzEiHdX5s/rMm1gjOeNmRuDQ4ENfLcmueQ++SyfEvNSzlDHnWDJeQnUuZZ8dYJjii6LB
+xuq5vMHe6bPa/DubB9Y/9fOIfKlc4UOZ82TGCq33Bi+eOw6Qw6uALea0z715aKrKJSJT+Mfe7pZ
/uuayQUJIVIjvT0Sq7hOnnWjizwM8BIUOX7+btG6PgjIP7/mzd3+oPhKg6PfWXdai1+5dUNpqpzb
DeQ1DDBWMbz8tjE+SXPLzFN7bPkNCidqUM6v3QB0De1lG4tcgps6N2DfsgTuLPQZazYh7eh64OYq
Sk5efQeJVG81GQjlf5JWfbGSqcpgqdkHUKjiRN73jdtkrs0kGXux1BMrItMDS/XdEADAZIgyTeIr
S7z1GCmxH/QMjH8LfIT0sDGEGKC2x1TXtofHxM9QsyXVwneAqvkIsp0Wp/uvLYtwfvIR/KYAdN70
52GcwozAu3kOS2ljsvqKzzPpL+9uDYd5kO1YlI8kIZKAprt2VtHLtVvjQ8+SK4IUbnLnqTpk1s6Q
Jj8Rlzv6RtcBANzC2TKvo2hCvnyfu/glJHXIik9NdD1z6SHFgMjUDcKJr5/KZwJfUrivoRzZZlVK
bFwnGhY1TlvFskU8EcKWHdncDWE3dqXVWi/eMOpwWQ1SoWOw7eHZvmNYgX4lyBeCRbUQQxPi3Z/N
8Uf28wzdahGqwnjXO0o/BUqkgxrfsd+LgWYhSzV+EQp3NhjjKxqVIhD+d+dQe9kN7vYFwaPTkn6P
QAePKmny3i5XnL7WAR6wF0IHk4tZT8Yp1umOV74hLLX99Pib95CpAB38HmHA4vu+r8vPEK6Bl7ZO
QihEls74eSOd4EXuYH+spYrOOV901NCpFawdbW98BRGDegsyEiDzkugRMWmkRrzF48JXeQb2Q8l2
8V8hHwbYFza1lEt4FqfWCdyB2CtLWe5iSWhAUMDx9oPP53r/cqmd0VtQcdhLKwS/GxGF+8RdA70K
0stHGJbSsB4vcnNFDrXQ+D0wpKVjsnO1Y6cSBobVRMyMh/dNC4K44QNYG1b+g+OAZNlyof2vI8PP
wbMuqgtpPzlxA13Q7HpBMfXqnct2swvjW2PRMbBZWsQw0PVL84Jz+j+ic1wXJzYWBJnyfU+rboJo
0CYFFvYsQr0PuPCsYXVHGkKxWw/9SGWYUYZgMw+DE+bYJjjfr3fbl00wq6ZNt6ktQb8waq+SgxZY
yHGYtTBDsaNhUYrFaQ5VnUsDU/vejsU5OPRsl3nHU7g5CLykshQqHy91ESTD+uuNdsApzMN0Vq8l
znpJHWn41RAGs8wcFOFAKLpo+AuvW5FAG/QitzrS4kyLt6B+pgMxtDriGyz7Oo7BEeCBYSXkozmZ
yRKk0LHa/O8lxDLfUbHjPkgZiARo1yBOePxUwrYqDBANBMD4ZiauyA7iU4riN19GCGbahJn/saCr
fhVjnG6MYjavge8ZazkDojvMAiIQNneRsI5OeWIDO0DvkVLHc5W3k/FOBrhDf/QGi+mM4A/SsNB3
FLLo18dx1k8jKs3Q0l3uqIfQeXrd++bq4QhqehXLg/mAVWtcg4vwi/TQMlDGTRaFj7HUYDe1ifeU
uNlGu0hR9fO9EEa51If5jNmSS2t6dyM/0gwXh8Nm0HCwxiFuNc2iwgXqvT8YK2jnmq1Gps5Fiolk
kjN7hkbejd0tYOUZAOgTh0hDeH4NkuU7kkXm5mxY7pEU+RKdGWCGmSCrjL2I7m0qpfl+1X9AsUup
8AE52d4kZskjH/A8oHA6QHmzu+rFDgJAuQiUrgNKG54YE3WIWVhTzO+0/QLErIN5WHOPxer8qqh+
nu4i5txrI5Xi3TsUoztgn72dotsmH4fMJdrmA0Wepwhs1RbC/4dpN4HBC2Lo2I5AXOy/+GlQaI/4
Z11KTyb2WhVHolC4DNLk3J6TGQjLYw7KHqDOGiO30EMNbzoTtQgiKICkHhU/jOARSNnEkFbXIypX
vp705yfk8JbGeiY5gaedyHrHbeV2owA2bHK66A2O0qOMm8eC5lFbKnGoPDVVfwQB5r1Ar3SzbygJ
cYdGijDxTHFqAE9FmrUiPqwnTGQRnk2dgRVyry12JtS5+S4X25YA1DRG4emD3eyAOtrTrhQRJkxW
wagSyb9lsBqBCz8WQ0wNH6AbZY8gGmjWAyXSkUoME3X3k4CGPHDvg+iNbVHPK8hA7+uam77kYgRL
lDXk42OBGCHhvW4hALeD2eSIz6T3w6XEfhsR1XPCp/q2SO83JY5CdgHOPy0FCeN32lQB7PdEZQR4
GbZh70kUgvjBiecm2zUjDQjormbqPy+0lIAcCqe4m/apivZs5vsG2MgTcBS3CzbZSBcPmQHzr94G
VkbixY46/aez6rXi3z5LOSJ2vicGmK0ugU2djCaSi8Ita1LkjvqEVYLq641+QrnF1E19gbwKkBF4
JvLcQk4o7gN6ajPZexBg0HZHnKFTAZANb2B0FH4a8P8dxwL4kbMbUsugcoWxyAALkeh9B/qMoWGk
hwFl+CpjmFM5ASOpYLzFWsLm7ngd0Knu+w/Rvg2OA2ep2Shwz16OZMsNkx3bqWPCGrF+L0rmc39x
GC84mh0vu/chsBnPfh5U0f4+ksAnMWGEN9cBMk75M9GpnEkbblxZIoRLH/7pxeIxkJ/SWPIpSqwf
+LCMAwcuFdWpaPA10siZcZUD6etBE6rLMDyU3i8wT7TMra3sAyI0RhQZnbbmIWOV2gsWMm4skCZ+
Zaqb48wbSQNbjvjkx6A6JxSeTw9nc6a0bJdm/2bMsfZ/W7Z9KZ8pTdAK7hLoyzL5c5tTYgP06X1H
KvIbbMoQFjVl1ZYoEcDyD1vOfjc7FeEyhxkYDjKSfnl/OJX+NNpLEY5WSH6H0TbfKxQPGwpipyFt
84PI+UdqbI7Z6PNilUmn6/Gd8PNF6iUzGn5j8dgPTPZ5K4FltbG74zomY6FT3IhRNvKzc11vUqzT
JwQ0gaqLA7S/RcP1JLyWO64MjOB/ZbrJUVblA4lQmS9vl2/qbl7mJM/0A6XybAqkqZM0Ya2aojYD
kuxGgskdrVJ4Il6s00J0ucUrSkXHm69BFglQjZCrPkEr8a3m7LwK8flXJI1Adf5xbIVPd4Af6sjt
/0pM1vDpkJ/6tBFamGrJr3DGFBoCTRedv+yTR/GrpnuCqWnj5fuFv2FnD59m7fQ+aG6EsbLIhuwX
Z/9s22Xwwq/t6kYNbFZWii92QIwJms/k8i9AuNnX6yux2qjmGKXPzwawPM89jCifIUbZdrvQStg4
d1C2Jydsiam4hUPPJrHgx1g6oCkQ8kVbTd/xe7nRL2RBpEC4KIYOhYnSPet513gawa6ULtjH7Pg7
KCLhoFxL6VBLZ31K4CsL2yOe/q5Mm01Y6or/q3nxFSvBj/Rw1lRl7bM8+lzOAD3Z394X6ztFXZFD
ryqxaV19citUHMAQ73CgIpsbigvqQ87zbOzSn2Kkx7Mrs2zg6TVaoNxlsKYFWS75n2WgUvQzItfE
dkUrYC2nFjrR2S5tvJhLMwIxqbeFW0EpkfqGDMenNuujW6YaSLCfOsEN8rAijZ3wev3oPBfJjhWi
jNILxRCV/Qj1DArMMy8rIVLfcpmPrOSUHjOAVBIm9hqC78XzwR8JC1NSdk6xAS0tkDaRt6apzmjH
vQ3DJUoYEeyPZ+3z1LjEQ4mfhFxdAi0oKiSY95vCDTIorkIDfZBE29DfQEkbrG1b13lQXvrVMLA4
2jgotFNPjcvFxY5gvu5v113PYiCK6MWnS8t9KgNVVBLoeLj7IEb0p+/8Juc1AJYpnS9vRayPvSay
MXbV7kCte39NoDDiV8udluovNEPIFtk6VLaexU/ur2HiFFcZNDfZdFaxC4lyRlErWlyufjSO4hpd
cD/kz3T5A7sbCwr4mMaGGcPv330DCLN2yem+7ZY66b0dngb77Y3aEmwT3+UvrV0P8vqk+/lZ8ljy
jRK3jraIMRtFdMEgZppCtnAJuGN+FfaWxFV6OzUszYesBmH6Eyes7DlsYVPimPUROirT/47VitUC
l/0p2akpN7tlobqgciwY5XQ91GxOM27cy/IbMc56MZaO3PnEuyx7963pSik/Ba+sJcdi0Y7bCfyS
KGCHmhIL6t+HDraiZeWOQZ0dxF4TmfjMb5iCLVO3liMSi/o5hf/QWAO+FeGVBd+lIWX0jrJBaRWU
j7pTvc/JoinqwhyMmqg2rKCtU8GHCX0BBrtVEMijfSRkeTcuitEIpfF7Q53gu40Jb2hC423xASbc
T1CODANxQq8tEVK8XOSwwuz4wIMwOckQ1gCwp+W6wHDABm0UJ3JEjgI6zHe6cD7KkNPSYu+p2nHR
Tw8xdevFxk77g26GKuawVOSIEUP9Jf9O7BxBxpzwmRFMkUKgrJ4Y1w2qIy0YDfn7mwuDVVcsAqUH
mMYh3IKlZWgRo2z9Cv1d2AFfJCo8OiFOCw53Cd2mT9ZaAckqm3tfiNRImGGokU+vYWncssy/2O3a
ui3KUrKMO6uAuWZ49TGGVK/sp0bK0z2jGA6jm+B4isk7kuPAFRl7IkRp36f9cy8dX42HcouoCLRF
N9eaTM/nwCckTUM9T8CuI328J6HzEqhXC6xwFLF2GpBOLWZNq5UnqzJhZckyeOWsRCrAgqNIach3
AXkl3RVbRct7k4aAsImcsMSe77dkCS0TZEFdFOhKVJ9hmX0gD9axM6pvDPTh4e3VfAD0Opg3Hdsz
XZ1jCjB8zaTLkXl0iKi9V+nJ19v0HcZWgA7pTjGdzJsekfeO3nQraKFYeOIqq1V075bB7Gff6k74
csqMY7ZmddTdtZzX7mRx7j4duLlOhL3ivfWgY/CoiJTsFhJpOehL1ar7qDoKDYLii2A/bp4fH78/
1a5Lz0llqah1mpOpDl86QdsAvJ5Qf0sb7MhwBKERQqGnzq6rwF6onZc441cLblauMy5gZDA6Bvvy
k+m1odrbHrpirZosUfAWiJ9p0d6VXZlohppCxfROvurVM6ITgY4aLLScT6WQLxqcJQOXmKDHI0kk
kPMOhJUkry8H+CYuqovZYsMm5J71SvOBBQl/goS2po/7cOJg6fkctnhU3/sd9stYuc5VsWAGtSfh
jaT/AZZCpD7cm+4ecRuBS9PJ/x/WxrnEFn+kkujfTJ8vck4Z/fwfYN5v7dyiuMngBQAcoBW2g/Dm
NxnnJMhwitznJdBZ4Vmu9G9Rq8M1dHlmn9VhDGJB/GxeBaZKo4eKiqHm0sFVyb9VGqAYEXPL8nb4
3vy5zGAsyo6GAr4Qjuk70bQZe13KEbEoEI1jXLZraZp8VWLO8wg+7NI6imGshsVpxTHYeAaoNnK9
fXIc5ZdJPm/ZdcepQMMpk7EbDIw/My8uPxApT0ZMHfd+aqwJUIiGH5d4znT9enjd7T4WUQUk2LgJ
UwA5aRmmPmZhq26x/nEd8k4Kpck0doMyCHba9jUJKQ6vaXJ6nP/k9to/lwPwVTVBsZTKkf9t81Eb
GD9I551vU9C5xFwxVIdeHSEnEIRrYiHJpEd+YH79exTmqM3Ozs47943PfcROYUtiNofj1FGK0ZHF
bBwV1O+sIq1ZHwXnLfkow2uF1Ly7pdeqZyLd160J6dANJ11dLJOm2IY/7DifhOHGuf3/KUwEKaLr
VXM79j+fjQCiZIvECltEA3o7eI76duKm9HAJ2dq5jR/nzdNI30ILCRpWca9BQ2eork0KjYiBKLWf
4ZpvswAs6zMpv3Pjro83BDlayajnIzIjcY3LqoLcSuR0Uh6bVfRu3/ivlJFaip2NgGLma5Fo5Oiv
REliJNVpMp49pEUo0ClqVEoTeAy+ejqB2/GWGW0RLZRFb4+Xbat9D2HMig/31tLvRfRZMIw1D7s+
6z94VM15sJHFk67EyxUp+re8SwbAK/d8IQjhxorQJk9mPbj2WmRAjzg9/2oLqjUDuYrQn/nqpZsD
jEvHoUy2KYXnDZ/0Aeax8Rj9eF52SOjOm1woi1wUqiYs0sslFZm30Yy/9TTr3GExP1+Nc1hTfi5I
G3qTjHDb25yxIpV9AhCGRsR5QK6YFj0WasXJyomh1dDFNeTcZymDdro3Ym2G3o/ivaDE52Uwb2AW
Jjqz1RIj2B/bmcPYA0iRdFigb7MWvZYebO6xqV/ei5LTfoO+axC6lalhQw4Q8A7cvnZQjeg20iD7
REUoSN2wDETTuY3G/GvLQgZeDbgcAIpaSnr7UvLebLDgft2sPqNQFPLAUBVVgJN7FRoUSAUU8zRP
LzUwi5cVTBL4FNkbCAQxxrwe3M29xnpHkhuQwimddRJINqmJQ1qlaqo0YnSzk1awERp/fKPCys5h
9ZnsWA7LKS7lONkinoKHxKD1kgieG9V5+bOq4IgJk8NpGpOuGJ7i4PieGWCh9DICl9p6z/R3Df1b
9gdmzmRBgKyggnzIh8Ox2iN7vTomRtHdLy3HWiuySOmSAqYqNN3X+KFkHdOVR5NESIkMTPRr/P73
8GOUexSSTvRElllNcOUrDkKon1M/4spKSA5ZaYHjLl3c8XBVMCkypp9+KnnExr5gzdOubZKLNFuW
WQ8FDQ5bzJkTfY5XI4wsJqf5vGqs6Wp3Qy709pDESMu2vMKpUniqLkri4hagQUjdphvd869UTfdb
eybrKKF4q3qUZd+NCOVZr3ma49GrHRgsNwy0Yxqo9xuQIVO/HhCeGz56AEwtAnjSiO+QEJCFdHb7
yS/aZoCxHBW/afPdnEZxRy2dE2yLdbdD197sZibKFW2aSClF3myi5lj9QgsPpZUm8L6XcbHHp5/s
fihWsK8f18WXzq46dB/bB5oC1ym1eEzdlKFTipt09j0JRShMy25/P1aX/VOgApObJSUrdtK3aSXZ
GE4zyLxh8cN5DmQoSg2vOm4eumWX7I78xSX19KE3p7xj2O7g94BRLkIt+HxPr8gQ1Y1oOx0NqOVT
E8N0bd9Fq8KibgaIwrIVn7Wct86FnjyLGnsCSezIng27iBOeqk4TsX6bxo71Nc/Yju8s7lEHgBbN
skr6fWlLPzgwwjqMiulpiSowYalBKw7e6tV0Y2NYe79pDeZ+DYrRuZxwUeSphJek17R0WrRDJQPX
j31WmpWcXy8tErwgpHcDMCbh7s6w6InqDOYVBC+a7TJ4g73ZDv8Np0P7bMgGvJDdN1jrvp+4UaSF
KUNDfGyobXRwpJPqjcItJ/GW5mBnL+txn8xFd6UW92lWMTfjIeYyMcun0KitfJg5e+Zss1wunWzU
fMlPRiix4GTnZX6BpUbsDjDdRHw3bwkHjcdGz5/ZHyJTS8HK5syzeEwXgwrjeA7njwx+Igk0dMrj
ooLKbX+7B7KuJUw3R4GRpGy+NDhI7jjg8KGZo2vZbEad65OpkIlctzUkujvIoW0h2gCBZNZ4CUJ4
1BVglrVFw0J040d05EHSD32FLEbZwTLo+Td6vGO1OpND8kVR4frghyDxu8pKvfTnHYDJlvssEYCJ
kcb2U/upk0i1bMYgwAeHzu1iaKOvSSpJZPO9KAxRDplW7V7O1Qw5muoZvevOiKJQ+WovE8Tu7AXM
1O4MXbSk2VHBq/9GvezQVkyGmRgMIufG1exU4FGrrpbDVP0ZGtSyJH83xE4w7aQZQdEuKr61aR0A
HYJx3XALNf+mSWa3QxRHcZ7YtmRVgwK81JsBHhbnWyWamt0pRcuACM24VI3J2J+KaacVPWGOLNAM
ls8+u1x/Tg5modAGNJX1kJK7YztnNj1NlXR71aADmrzmX3OUorTX48alHZpGkWvgEt5+OmteAyow
enzNIbuHHvBW4gHWpgBGka1Lu0E/ldEajU0xOiLCgzm64Vjr5W7jUWV49z8QNR1dDQ4ZWBql8lK7
B55b/BviPJsct/2MB0D7OKnGbywASInCuasOODuVsNLfbV4AOa4NREeLR+Inhy4emTcYbyzqxWoR
E/rIUlZDWdeJsT9vXFdouuFlShvi8NEXZbr4GT8W5+VZGehnkKlkty7x9UOyhMNPCtr4q3Ey3VdK
XQRFTLbIpUGctWgoG77ax7iKI8qXkvcinxJrZT0WtgRmcC6neLKI97+pRIb75bqCN9SmaQ2cRXV9
/KC4r7uwpoQSaQ81M3G1Co882Cn4iKXbBkmVC2AFms7JeGQdATgglcMx9ohyexWLmNIgdTmIJxBk
fb9ZEB+MHEg7+2MEKWmHbahjY1EUgnxbOej8e7O8OPUXgSpJ393c7dIvwlbaBjW3+mm0aahTKO7v
mqKw6bkWF2Gvc3LnumAOlljU497I4hsJZnYwTq7pDz+EXNYMuw0eFchezYUzWNIrPmof1pAUrnaQ
CTBSXoXZ3aX63JOCL7+n+ppzgqKgQcE4s6BFQxsJRbzApCoHUGGXwSULRnNOLN/SyQDVLqEEyoWi
0PFoGOQmsQHTzoZfEV6j3fvsE/trmFQDqyUW/F/SI0zT/MDOf/TGB9S+/hjSj3sBpitE/e5nhDUU
aLmcGLRexw18ZzTAEcaPk87mchHF0ZOulzSuSNbmgtMPcpTr/tdukXUmaVg9OfFsvv3Yw65PCz4o
Qt5xa6dche7bH2qQJgSbLIdDNOElbt65IcQzDbEjOvmlxcad3D1uc/9kV2O7j2BPH0EcVJbB9jRp
lOQ3ZYP0E89/kc3WKnBbIy6DxCv7qMTYKDc01vD25e8Uobj0dZi07w9xeU/HcTKGlLsibjOXa1Av
PV+IkWLBvB3RC21fNBoMY9Cau0Q+0/YSdjGvB1bXPocadjMJVREEivPLtgWdiShrH1SOpURkOU03
ueiqIFRAjIM2zt2D1a+17lYS8RpIbnJpbmFOKl0M+d6xF5wfj+8axZUJpnthNAGu+LGdEQ3OE15h
21cX0EXsr7kJdP05pv9ZnXk7Vnykk+n2QYjSn+58tGFjx2kIZ0IC8r4h8RnoBqaa3iY7u5GFX16m
i8FHGtltgV4w+q5XQ8ntcbVMwmvR+Fua5JKXNnwcpZKp/0XOFp2POZBFItalTTFpgI2L77oDRWet
jnM1MPXgpCLyK9wUCTL9iaPhmjiUlxJ6JMRh+0kz0CFllCoTLez/13WQntBzbVfKxdUG2SfYDUG/
L3vR88TQfFvP9K6DYJQkPwvh63Uo2q68Thqztyn1zwbo/2INEg5D04lHjuAtA6IX1PF5U2CkOhUZ
LrK1kTvpLBExpvAVaIKCMNu7vCALyVzvetxipqHF06IlwkVEg5aFrbNwqakPmRUJU8QlHzTkYTEt
N2b9Lmnksb0jbHLcGODOgFPUhUDPxbcgr5RSHaPGy3BHGy0r7lgktSyvJ+NhVf6fir3ngVl9koaP
zzYzXru++cylgG68mu5F8GJN34AlGsfwrV5TnxUtomVkhGC6wyLoXZF4xn3g44Zp++gZGyl+s4kD
pE/ZwjgnJmouBEK0xhzBENTWFlBlb9SxddL7HlgWd/kCgkttCzXUZ+p1k1YkeHJES/E4H1a7PvL8
U1ii4Jm/fbqdr/JV5UyfNZRwCVTjsVgmA0hZlTj8WzUuA7OKfWmOXKNU1JHIRBYp4xbVi0PuKtEh
Id0aZ75Ctmh+0VPm9Zo0WD9jmAY6JnRWaRTtFrmvEJvW1CBeDElkXPIj0GTcfeTPX0dC4JsrY7fK
09uy8p6AtxegH2fYoAkqA5/ccI2I+hkbK+rsbUYhbh/r2EBGOkpvHo47zOFfAfTE7+obmqgO0/zJ
6s4x/EzrnJySrKbP7gJNt2FB7hV0q3S8/1qkAkwtKd52cvW3XX7ng3ZH3OuDwyr4PnKU1ZgpNpIn
VA3X+hmBpEC+q7v970N3tYRky3NmqGBmQeVPO9MMu2wbajp33eaPjBw9f5YdQDr7jRSmzKQBLYnv
wki+wd+2zf+vG7GnuL9i/pn4Rw/wlKDBcMZw2ZsrY72PWjuq30Ke88HbII+eSIXo3aPj6sGGzuqt
Lok7jEHSncKTui1TFOaMjcdc553meUquHjdG7wcInYW8zGAJkywArTPmKEbpBO/aEMxFaaFwEM8O
O0o5UpuUFskxB5WuEqCTvOuun0fCRsKRb/g4AEXqZIMnFbZgcBfv+CuFjAiXr5jV3UiPU7LHOFmO
v+IZx5OK2+XhZPcWbo4rQ639YM31C5QQFFxNukbOeR+cUbJfEh2M3O9R02kelumjlE9sgjkfiT1C
iD4rqNoqBBXRUzQzBqBEHjbqLwtw5jAbgZurfsbKg1isYQnUJZmHnN2wTH1QmwpKZrcmYWI4XTK8
jajgMRZNXxiqSNr3b+oU7oyhsiXjkyii4GSouDgYEZXbjHRS+HuVSFv6ml+Ty/sNc0sfwFhibu8t
KKaAykpC0d3yX1etU8jdYxVveMkLwGr+o5br3owrezLmiesYUW7kuX7XqUl+IHlADhETJcAs1lVG
h8tWGpw0kot9+ME5UOWG1cdr/g3S2rfGbSmoOMGLnsWnV+Zwlc+w2vq5636d5CsHbCIGGMPyokyg
S55HmitiwhzrwMr0qXMxrRpRO+ZwsWfSP8+nLnXxaKqYXIq9NYk5PV1PTWvovCmFJO4lH7AiXLNW
8V7hj9GrbDd6qfj0ytf08b/StBZ4kSMVVGuia05VTUXWXENXdmi4KZPhdKabOWb071vHVOpol5up
bgWVWQs35QJlDi5BcR/aL3mlEpafyBkOpX4XnwYnkOGcuxweG6KYapqN+UaOy1IyOnPTgN6ynyKU
SSmOBaeshHH/7yHTZ1gigWfY4WZ451jhnqJn08WEo+PP9qFqbmve3R4xfWKPFgo3VGIKCTV1MfeF
YSHkRaobmM6drxGaq8jRy8b/zjgIF2CzaFMLBTQJa2/vHL2OvUH9liAmFVHD9HErbyOdHI6IY/da
S+25XirVfG36wcnw4WqncDWAxGSJsHVHvS+W9PTRKSCg6aVUN21EvdS1Ml/sVHmsqzBPSNI2JFbj
9EzFiKiX1Hzq30TDqX83tvBgI/epePr/UWPvZDOvPnKBxDBaegf1o0OezbzQjKRggu7lwbw77pKm
1stfE+a61vgqP6I1dz8J5U9owFh8CTPY2WGBmUkFXeVawTKmBQ/i2Wcay3tI+Hp/PNIgEtMWjShr
dgem7YJlVLdvtgr/UU3J/4KELzNrZkm3nOpq/d6MsJ4w3lOWBFlZ7ENoz0hBy9mLjhnKIy6UdjF/
j26Al68z/LQsMS1BQLft7V1YIRP5rhulWwIq8lSpIuKfkEk3FBBSQhRJ+HBKwWAL/um8V9Z+YzWa
tqOeknnaNXTjvtHfHtbExAbOHxYxQfrLR6uZoiPZaWX4vB/9QGUhZfCddAbpMc4XK7XhNhH+O4xM
2C3K7l87Tfffz1Dy1T/7lHeP5ht+VE8Hw+cmN6dS2Xd0WfKtRJfFC9sZFWzIcdjNcN/DW2F8TAzW
tbONy/hpP4IfR+443SEg2GSeA8DbElEfUaEyP5ZFeTYouTGS98XjMnaHfqmw3/itkoMgEOFCEq91
8k36EcbbF66md0bEsqRsU2/4zvjrIff0ZUIVhhk2sI5mHRgnLY+d2faoa4Cle1eLSONZ6/iYChEa
gka8lszjo5KSYcuZh6y1UdOfjsKTilmy7JI16NyNwk70YdYyU7PXCD1zEI1gwci+dHVcoax0QgGK
qK3LPuXkO5i+waSSlAGBZc1MpmI0YAs53SCkOWbxwopPOQPDw9cffarVsZlEXVd2OX2/FdxXD0Rq
NZ7+WPJxXCQS28IYl6e0I1d0wgRQWJNw7RLmcvBHOA9NEJcM9Z2P96TK0KAyjky+HOZVZ6KoeA7F
4Sk3cn8Kxer9ghuxWwl592aW6iYxeMR7D/zddrBXKnFfYeTRh9nkUOV4Am1ka9+pCyvXiCX+KGh9
keb8C5prpnTiZC+vFRc3GtBqEWiGXG5BCQ+3lpWl/jz+n1BfDEXqgkm8d9AnTsF82I/E9RYv+tUw
s/Ij+svTuuVvgrzqJopfn8ywlQW6Jnrjiu8B8PCrUpPr04P3G6SON583mtOMyU6XPxS2Gzg/Gafx
cplhzBPI3JlouDsm/an3i2V/N5A5wLRIuxOnKrXk9a29d15qquriFT7+P9sm9kQybulGgiHBJ/rC
lUW2Gx42csRLfLARL3HsTm37xuBCMzfHyVJdXJbTNhmFBENMtkadLLTPYFL3ldDGDEFR1u0D4RvJ
/KCSTK5QOQy8dVHOzEKsAs/sYg5vGnlQB04SU4J5kKGVCz4AicBxy3DNH8pmXs13spzjpYs7jyvp
WXOXSXCVNFG2ibMZbACvNV3xx+r8w0itzlaaCIy4KRNmQCXnPnPbhM4DZ56iNLyXcjvfctmUyHnI
JzurWuhKqr0eKuevZcn1KYcY6vn+vJkU8iRW0LIbmCM5Y3Kdt+Tcpli1JxDt9TaCXCZcsYen4Qgr
FPP7rDagI353fjDCU4BaUZZkcSHdmC7KcxlF+TTP9g4W+tzmX8Cz+NMpvcqfy4QqjOQYCdcVIZ0N
C1xZ36XthhJwmHfLzzluIyJvVtCCeJOdCSHSrTwQXibNnN7tBbZSs19a0wpo6ZNx0YpqLyaeMFr6
nrKEgNI3vaYeNelbLhXk/P+UUI8ACK3/52IovxVL3fZNL/Cj9hq8DWq/zbjOQf/n0BW55RG03k36
NkSmp4L05114ZvMcXWnKVSyWGnPbm5tHOcMCiEe0ThGj3xth2cZVCFn8HUIZm+bgZzn4mNCS9u7m
IWqCjYUuJL57PjIMlrm4atB61hw8qIBBCSc3+1G08AQEB7Ps9TCMrK7DkslhVx/FT4h0LjZ2BSU/
HJ0ZGamxNXowut0yu4RlPRJ5Zg3i8wZJ2zbzNGWzSECg5T29L4UeiDyqYgfJdxQz3bKiP2NYsI9k
fucofhK5hc8P7LiiuLGFV8WeA85aRdtLNvmvlULCE3vLX1kngNolkUK/Iv/uGaFFz+LR7LMEdDUf
OD3vpAFErYnrQJ/ZSQqcsGCI9pYJUWaQimTKmteDP9/ji3Jb+4Zt4YAjaP3l/Sv5Uef7DQ4Cyame
bConspZPl8CNS5ERhfoQN4nMkS6hIrKvnpszUy37bqVGv5usjcV2aWfU29alGxPE4p3saBVAonZj
ooSMnfV+QFRdYWLN/k1fkjxIaxp6t4V/yxjs8Fvnny1KCUXt2AzgHIbTe1q9z/dG6NG/VrKchVsY
rivZthG01sJmRyybi9czSBRbKVEp1QHa9OCpItpIGT9kGbyhF9a3RpJH2CHOMBVG4rzPgA4APKXx
f9vod7qbIwHd75VmSHJFg0WkjDJkIFcdiS43yhWEgM7kt+MKGUdKwfQLa2Kz7//MVHfcxOgXyfzQ
QE3daPESGK3ufvJAvARzBFy4D7HcbUOJ2T/dVG4j7aLd64aVWJMHCdIMS0un71mbAZnQGmQfzNvS
J/cgz1KfzJyswL5S6GXd9/cLigyw2fQ0llvBSg0XaxZokXV3Rrvl60JmnEFQIxZZfXAtgVo5VB6q
8gACe33SlOy9qxwmg7PP3uGDOF5bisH9qyvUIsg8BdIsPtp7DQVj9203j2a3icU09HQqzJaR70tZ
J9ajbYJN7baLJYDCVZ+mwfXL3Zkuasc907mOcr7jkEBwbYR9+p7+FB3kRu0j+71Qr1GaW0T2YkRt
zm2IzBQ9IED9jVO0V5aoVJenC3WCjw1SO18aejWiQef5y+Chp35ecscDwnCx7gLGe5C22CoQBVT6
eq1nBwkoFaRKikEzc7xCRitN5T7dvuODvaR79T/m1MNRvITQUS+ml+6uVlxJGk/k/IaDK5WvajUw
KP4RufqZxxLFD6tC9iD8cADfeThspuRh/5pr+p+GbzeV/l/tt++RxMPufaikcUlfD4nNK8EfZkyS
hJSJQuGzXTUmAHVY5UgdO7bVyK9zbvUggjgObf9ncNNLteB6NjF21zvdnfMJ81d0vizw3/47kNSR
XKFzIyx+YfaziQfphaTnbRaRyhGrIVCMgOfNNo9GT/9Ki3VcoqCKFM01nqIlsv9sKUnzySZRfMGH
gMOHjVbnmzsQoKDm4wIzDCZ34l1+lpHt98mK//7C5wXVzG1UfCMMkmVU55pUB1bvIejhOgEyV7wK
iseQd6I773d1bSRTpDqqpi7U53n84t7FomRzl6uzoLi+zmHvkC6HcwFbhrMnlF7vZ6AHpYIjHD6K
kwxTX5ll1WOP0ufpYmIgkJDGYlLaKRQNnXkBCX/aWzB1g92ITInQxRBly2VoFtVji1m/LzNg736r
hlcsoG22RY5d0u5bP2yDTqrKZwMFRUeQD3ZpX8BLeyXPgcigSs2MKkfBD9++UvyTBM3hXPkZT5Ji
yovVawsPMNIDYCHbzyo9c6WEazv+dJvtYtLzNd+S2en1zUKHrHP8K8ySTh7WW/6OA65ig2T/FUEC
7n4a0B+IgOsxl9EzqkjH41QMJzWfk6l8GXFVLvI2hz0+EcpeozOkhQGY0eDQdgxUJuT3QluFotD/
P+dxunEtMIEGva8uzSwxg3YkE6SC3b4E7KiEmvyWJqKlwAlZ/KylsVPKxZKVJ0uZ6G166fy6xlqG
oydU/DP3REEt4C8oKfeyFMGehErzWe9rKWhtgx7f3fOdZYsJ3nRwu5oM1lC8jekpNLadBUmPO+ux
KtFyXcseF3llXReFLe8rviKcaYjMG01Grj911LmQ81sfk0czzpIfaWXI0zCBy+nc7hwRBDLUV8n2
r4FD8wLDdGypQ/VeHNvxj3qX14YPgi97O/yrAb1Z2DBKnXdYr5lu6H3Yez/mmdwPwGNhY1LQsfaf
+H2ztYR0XKcKhr+KYcIfIamIM7+B0BUX9Vs+weqJiqa3vdvRCdmLc4+ZLvXieokh6v0e5naNXiBb
Rc8t1C/bmoQ0dE3FvnUWN5cqVIwRsCGkTGvH1oW5vM/WXXNLa25MJJMwtkVtgXqns7QDpXnrMsbb
Fhb+2zCn6G7q/GGz8oCPlOlFS3ZZ8xkO4OlOUCVhZtO4mTUzdtCHL9YAEPc4OpwZhcKBDdPZi6O2
U1irLYI8XUsB7EzGs0FgMMxDL7qmZst2oZJ6aXn4T8fTw07HSG/LB42OTOlsA7IS8G3YI6FIQHvy
/Iil314TdxHgx45LjVZEynfDuQs1WWbAkmkG4bYxWslUIRaBFO9Vrtk8Vk9/iZqZhqFhv7BhqZcK
avUGb9GLvFUqWYdVY9ouLYN/eg5iOjfiEnsfnetITyj4sUJthAKmgJEhGt+aaVGs3mIbNDRuzd3c
rr21c5b9HoWmhsG4DvpFXt7nWcUp6xAxTJqNgw9q5wwQlmgoHu2wKhMAPhUWhNtRMFs+06FPYtKJ
QnZ1kGnJnc5V4yPihr753vV9fHfMyDLBsAjdP6s7VsERiZDrbqEUtdR5wmi2OXxDhMtAtHrnIZsC
YfSo7En1kYELC0+f7t9dJMAT1l1QrxXi2PM6f14tIekghAoI6PX8v+oAY4QN+6ao950ON47q2iS7
4hsoNPWXfc3nbhjDThPZu0RhD8RRKJ2pp2Ylr8qQ0G0KUbGj8byvNzAcDu7YnmN532YuVCrI4kNy
T6vyMpNTtN/pD3egkQmBnCvwGqfhtKVVAohgHdF4YEZiHFo3okBlLBY8znFRvfutTjy+MSl1zEBQ
/P4kQi7Q5Bvj2j+lzYZSRZfTwEAdzoK8Do1XlnlMaIjpwNhxOkenlNikWmOxaMUPQC2UITzk57Zi
lJ+gTZ3ja8ySW/6Q6fJW9DMK4ZM1XYlDt3hDvS6gdYl32W2n/zkRqcaAFqb7ohu+J9JDn+0Smfjf
MkbvKhVk55iDkfFiAWiirK81NJHMErEYOKryhy7K43g7L5NomfH2bUpk1zVz/93yrFxxlHebZ6Ce
jJrFdoKmWmATUxHaLr9mButBFWxA0fsiKqE1Mx+XsrtzofbJ1U5kC0ql3XhBS9N5uE2yG9O6/f/K
K+mQ+pGXamb3IebVl2OZq1Qu1k7vKscIseJybwfVUWPW82i3ALUJPvZ2YFzFQCGfvKlg+2l6nyhD
5oIp/FwxIz33dYMmUm3KzpcyVe0m/X0eO1yUOda4eFQYGD/AduQTbx29oP1FVMox8UwpRRJvdFJh
osTGGriJa2wYr5oiIAKzjf9M+Ic8g+84qX6fqrkjkhxt/61W5sCGlaoHuQ6Hwtl3c9M5HS/jfVm/
K7NXfxK6u0Xd99A+w7PLZBLQgIKPgN0YM9UH5xnqqNT88rM9/2+ELQ11Jlh/QHFt4sfoHPY+ww0w
zMxXQYsE2YPuWZVPyipRQxK/ynTfMEhSEipa+ijoZ4Bh2NFsRK1Nan8Tw5rjzcuU35TmuSeyAe0k
hBQfCamLsWlqd82U+wRaheQVxuZ0MwSET2rgBg6D8ipeh/oGD4PtrQInAShlw2OApZULqX7EUFrn
xehpXoLcPSFr7AvsCdX4XhxQNhp4rFQI5aS5yjIbeUrLJO8GawNWJwmt+HfyCidNVoX3Y83Ud4/2
o+DHMHvHqAYngDeaENPf+saS0MN/uQJ/iY/hi4I7OPKt0v5+eGHqJO38WRKLN58qfNHH2PXAFISi
8HZPrw+oc7UNJVHi/pSF4I/MLUmZd3MD6J9r+MeeEy8NL8sCvce3UHQXOY/9ChW5Zh09tClWGupL
D1cQ0UkTjdYzl3mGsoOS5M19KXpGk29Xi45d12IDuiFbzSARB+GqpwKg9l5JFIs1c0aEjeZdfD3q
/aO/GGJRfTDVtUB1MBpIvaPnukUWnboZQFDen5653UjMHK3vZfPM5rNYmBX34YnBlLDGlGWkWhsH
mnGCm98EDDwcU7cZVEZvGm9KqXpQjvrzfT/0a/GQLnavN01Yjk5naIrx9NynLhWpLS6jMcTeB3mA
P1rotW7nsdWsll88vIBjtdzSyotx6Naey4ZArH4fsQbu7gvpVgUkQe4clnO/Z1892NdImgyfzzZ4
9duUwyGMCIIBQMLF6ib3/fWaovM0a3Abp72PdYRpm4HH7Ui7jEnCSxoNBmgiIHOy7TfE8zqGokYY
vnMF3+K2IgdnQfW0BhYrVUumLxcqYg4BSTL5clF1TWEym1jGVSTTxdKRBY8HokN6tZc9XwqcfJqx
PmAO2viyFwI3BO5ORtJePR+WqhL6Vij/6sFj+T73MdrJKGrwb2pwp8Sr0n9NbPN5erXb/KgEgCRO
geNh2AERtqrFbRNNpp+qmNavbAscm0jAJ/mlz6ZZ2JN1GQSOIkyhFSZygtbWStarzgcAwBdgdk1S
nP1cHdcmFwks2NBoLLrp2/m8DDkbc50ZyrfICbZskt72yu1Ni5xfKIvXF7cla+wSciebIRJotrvK
oaDpgbdEFA8ZH2Kuat9+rRx3FxN5GYr+3wcM68/yt2XonNTgFohcaMSJh09l2Vm36DYqBAf4r7ai
KbY20XBFbhnrsv1c/F5/B5Z+4M81NSgJVv4B2F4ly1d6jMSGsB701uAGLdbJyFnyElfT4Zac2f0S
7+/2x4SeC2Ba1NF/FykZNevwJyCaiBb0r6qiZvMumMouVMQeUby8NPHeRdld2IJyF+SZhuXN4Whm
FohReg4EbwBgnx0nZz/KCNACPKzf1MZUpczqRisIzjrl2VKy2oG86alz/qjZ7LOEb+D1JUKW5CcS
vgTlsi+gyncRUbMUbhE28nykAvb4xk5K15gokl9iWUx9TnskXNHafJ9z+/MgmOlFVti2PQF2odGs
+c29j540qJGFBozY0G8oOVMD5pRXlhRAk+zrYVhnML4Ak2yDiN82WUohyvOvLwho3nJegumOwH5Q
DI0Z4yEZKJ+v43+OxHTH7eCW8lOI0m8M9cEo4pqySgKRAiyUCI+9n3vmN8Ua3pNj4kU7GaWihVzl
AU6Neudlw+tFcqluNvKq/DuWypjZm9LZLeF9BKTYM7ypRm9OzBysnqiSO/83GQpVBGbF67TAvwnb
tG2b2IA2dCbkAX/VXCangI55UKBK1Nug8o4+zVX3W9ywCi4adE8r/GnlbAFm+DNNYt6uMcY0ypRZ
8dWFgqy6dkeHk7qc5p/cU8BMZqj8mM9ExFk82n+LHBg4wH9LVMJK4NYO+mr7l7CbJTBavN01a5Db
DwwCrFFNo5gFrbMW3wVn+8qtU4bSZ8gy2b/67zjAyAINRzRh3GpqTgBVUwgjmM9/VFxJUHDWgp/M
x8WTSJU4gxx8DqItFzYJCRvdcppYqUq3rqum/RNjbMT7b7LtrWPHudecvR3entohzMtunJFlLO0z
q/DkokRFZW+65TLfTthDnyGvFoj00VHHphZ8pzCKkMixDEtB6ElbkNY37lKoQGRiqUNb/pr6xWqd
V2ADQ1ZW6QhKIOJJv80JjmlbwzHgyzVHMR/wm20E5fxdv1ZrcRaklEzZDaMgJWCYcmKfXFuQehvx
9jhvRz2hPvPdS00bG6mANbU0FWslEVI2qk14GwHDI7mAiWM8GRO2PTdU0M4KZsY0u4FFEqOecp6O
0U2RyxGu2jJ5E5BjgNT4QLHbW3I8Vj3Lxg6FQ2INWr7F502NuzKUT3F7c04el0nkN45Zhbx6BiOE
GWRMtfiA0AB1es+WTBnADtK+FwHZqOWrWkRGhSK/OF5CkUM3zld8K3uoXOUNhLqXwdbWTUm6sbOV
KwLL7Lxn67+o0eI8D7RS0ABajwzBnEEusF/+Vo6b2VlZi44u49bH/WX0YwL/vYRhdm3/srbJZLDC
pT3RjFBxu9XWIoyDjynsneVEsvkoZ/kCVMCSL8zOZJbmv5JiQ3lUxR/tb061poP6gawKk1AUB9oi
HE/SQPfN0AQDcOVC7mwZERecGhFelJykEveNHDYcwX1n6DvfYZGjR5FnOyzDdOltEAGRU1Wm9vFg
eJar08Mr7qxOvOG3duvnLYm2nMiS7KHuifQf3HG/7O7hv5RcMjzS2nEDJFDrTiOM5wKjRPBNXRgE
QhZe/T1tyItZnzb4mxPN+/8scK4GFajo74xKMRUGhw18bXbxk6QZ9TYLKooMhDw7ZD0CdfGpnhRB
uGimaMua+hRrz8BGDXy5w1BMW6LtvH6nVxxkhQw+HYjrfX6E/zdnEnLLnPbiuqqsfwObeaUXVwZD
zrBhYevCJFx1/+/UPfQniCw61M3WxjA0vW0Zq6FHo7JjoUGC1Tx9xXjj4DRNau1NuDe8MHpC3Lq3
4UIS0+5g+iqx0hKxd4Q7IcViMkPbzvEZir2pBW4OKOVKANvLCw320Idu6MGoYkzc0WRvUS7BOMX6
CksuHd4k0qaXrSzomw0W1Q3rhIbHSGOhwMcWtA61wv14ZmH1vJCOpNhFwv11wM2sXWpIF0TnD9F4
iE1C+Qj7E/V2iUrJze5FiNqbvYCTE+3Gzf6P42tqW+AcWdh0QuexQuSkHDjJgJl2CYHRjdQxxO+q
qmu1dqo3CXNA62rCcRsrf0+7QcINrEc3qW2lPYLrYnCtxszdWh48Zxo4AN2L+9UCUd8rlzJkCnMK
0ItjXDV3fzFjEQOcGcaihNeeniZIcQ7vpEQnbAiG3X2ojLzlOqkykQH9KcgDjWTRh7Idhxr1RauK
ycXy4mBupchq/ESaX/8n9mTNuMBG26QQACEQipOSpwbGH53yhju2rNPTp1/PBtyRzQM4PM+DmZs6
CgvSfARKEDLA3IDDd7+0XAMUBZwtRbA4Wf6XdT1YNo7p3WZXIKFv/hBQC59GHf3CtexfGy3hpIB4
QMvHHtkVNeiOBOGBYJzZdN14IKDm/0AHPRQ8v3J1qWLMXrgjNzyXbFNxnk681SUCepPkF7J2PZ3p
dRHAruHPNICTuys3KUWToxHZyi/dKwnRY2PtsFzihOpcMpaug2GK+m6ybcJVYZvMIIgLW/Y454KI
01T0W2da5MHBzYffx67kvhleyHuk8YLOZZsTYJeuPs6z5S25rUnpuJf1dzsO0H4wedN0mLNxK+3X
ThED/OQhe8O7vWJQWkl+pnu7GmFRD25suPI4WMZZLRvtEhhxL6YLaQx6VzbfXEQG+2JHRbDlk5kG
TWFlRICYzAeYXlIYtbtt86Aq8IR4qwDE4KXcg6Jf+aN2sRRc9ZQvKUKseb30bXfvxJ4SYY4GkbYE
FuK9X8DF1pZWsweL685NsN/FPeL1dzb7g1EAyMvH4pAoKOWnJDZL8C+C3vqAhcWVtrhOc8OgMvED
IhS5SNtsrS/xZQZViB2YkuAVkxHNTkkWQ0l0WXLdmgMrtGbZlOe78FUkhTleUJAAAk+BNfmTgclp
lE1ReFSaTFzG4e/B2KYW6e8WQ2t0eA6QEIpmxUZgVe22AgRLc35oxZbQpyAS7We5UfV5cjaMM8GO
BgGwNvJrVKcEegdABbidvavb6G28C3vdaY1pA7VEMnyc9b6ZZsINtjN5v9eh+jJelPKiPC+4J5MC
l3swe7FNiAuuVJ93SMkGfUDZVpgqQlBqFpKzjiGnQaoGrT6v67CGMS+Yen8jIKYxVIrOJPjcJwwp
ATehCITbn4Xr9J9hVCKN2t5PAGQRTBa7g/EqtXwK4A+OKJ1CHAS5T+3jfE3QR8Uk6UK0K8ScfVGX
UpZJRRZhpQmBak0+BEjBrZrl2KCemFLHZK1pnfQFe7iwcDavMKeGU5g1gD7Lb34j2tGzd2vX9qs2
ayHw8yToISWOxBbVDznILnf7nNiqIOpYqsVJpBgSgeonv6gfGXfqUDVw20ZPAay+9buracIAMpnV
Lp7bPU28K3xyRjgOUwmu/Ce67UTfKYomdzNDl/rrpnxk1ZA17EFqYRpIqBzMgogNHt5svCOdJ0BV
W4k0rxgDkTA9njdoj9Wn7BnBcG2S9c0SRQCVkvDyTDi5sN8yFFPLab9FG1zAqqRg4sfQXwDRMSbJ
EnEpgyiBAuGkqRUaV/vrQm6Z8iLKocaQ8CxJpI0mC92yMzD92hX5BKow45Sc0uz+vr9MgCX0X5Q8
uUFUCQbVbdW7xiTszUJqic61UbFgcttYIBvjxG6CNqqHzrt0SjSCBuQtdFTN8EOLUJ/uNyQea2G8
Dp9udhzkWy70Cwu1qqnhcLnz9sXl0mza2FJHBVT5RDO7CtORi67P4Am7YXGqW0eh1Pz9+6J6wfdi
4RHuAid3CchLfPomb3yqe8a/IZ5Sjti1VK0x8QYkZDiTon3KVpfMivM2TpKAb8ZeATFTkXISUSoc
I4CpmRPGk7i2u0o0bgVbVA8/dBhfMeT0fFbf8dzEEoDK67ptOztjB9Wbh1zYxLtXN2TKUPS8XdTr
oL17x7w5iHVoiaTnEVNdRux9NCvwx9BAR9DjFfD03SgHVirrTTab1BTk9XAK1AmASgVgm5bfKAaB
6fkO85ovNcInNbDbQ5mAD6SxJqAVe9YR4YyFi4NbbGnqsPApuKI8DzKt2B77+K0siNAi8A0ewNGI
9wojpcrThee32pmwUewFj4Q4XN6WTCB0gYqOjVuliMc2QCkncr3dUwzwNSrWlp1C7IPghWmOoWMo
r5Rp6qEEXRUgOz8qizZlJYvymOTWmtSN+C+nl/jGxWzRIZ7wwQU8WuwbKoActQS0pQIS695hqmFT
bFswdqRF24FXMWvwONU5hEK6vxhfK/VB7MYXs+Us72OLQZVYRXLz6Sd+PLi1afjJwKDgmzFObqH7
Uwmk6fEHn8M+mm416w7+ob79jQnxzY+RuCbjGRFJAEbKqTrX9XaRGfYC7y3m87rY1qYTM9AJ6sTB
Z/9kJA7ChNlPrwu1SJ7F2xtoF0sDoSG/xyZgZLbtugqSd9Iio4FXNBhpvTiVPK7L87qiYorgd/m6
5EAoWdhFSGp4HCbQPQQ4fSTdDbPyIjbYdH8RFE53Yb5FmfGAGRoUrOvl4zKSUYS9rr0ida+w4tRE
tV1L6vfrKJAPPc424Qjeu4hfGu/yPgdtSN+egXfAsvDFNOIZxiv9Zomxl/Cdg+eyAUYH3sNY75Fq
M+d3hDhfYxZl+cWGd/KogPslz6JGo6OWgzo9Ovny5/nBSD+7vy8BNflVQ9wx893s3f0a1y0biGRm
JfeXH+vEGHZgbTtS1onjKKDr93ga03ATO6FyyDR0MmkjPHnegwzgDQPi1/3jxfBkffnt+aCIudYz
gQERNxAI5okpCCnUbJ7jXdtcEWXBSvc5HBsYGrQcFl4qURuLNzdmVhv34JoczjcM1cq6xQnV27uD
HonXfJCoW9ZvXEiBwtJtbTUBv4w+XXfSFFLRw4LzwLaKnyt200oYqQmuH8SKgyFg2uLrr4N86L0L
1iWTnMdaekmF06TkaARDyKRrMsh5AwCW5wlxhAYF9jyczavT6Kn1GqhqcI9fo77c4UCqfbok/3SS
m8OKTk0C4A9owjPnM+DGORFrEQy/X8Uq9Z6pIFpw/O0V30wt00lx4qiNBqgrP1AV4Drkw07VVDGr
zenbtUC2zqagtBGVggQ7QXUmT7ARMnWm7VtCs7ODZwXnqME883VIWIRuQ59y+xrAH+9e034l45MC
qqCcZhXNcGAMHhLNu/Ro17EDB5QEjPo+eQSmHZn5t9cORtEaWTVsV5Wn6FV2sjkZ3VKRr/EISpjE
xZpbM3d6w7GJhou9lfmrRN3BrsuJADJu5EcL4FnxHUxQjWdYZXQdHAOofBzv0bHvxt16UsIYq1DQ
Ps/Uy/hVZ/K2pYROhhuL9SOdmajSsoXx6hfxzRuNdvxDKLzDurqJm6HW2CalDFi1MAg5RTYfAnnO
WwLzp/XMOA26oiWBGIKwqe20JxBci+ktS5gD7HoudrpEcptvyYv/+JVsGNccaVOxrF3i1foqhW3I
uFTVyLk51HXFmKkkh3gKXPiGw6ftAv4nmOok59BKv4K2o4g80UwUfEepvubZIOLz/VVHxscwN1lh
EYevGlfBwH4TWDfhjShP5n77Af0zaJQAq/2rieW2FF5aBskgeB1PAhkwF7s+weZWyAVDRyYT6EYF
VvaUgB/752zuuCMu8ye6Qgu3BuuzDo2VL8dKZiPpGvenokH6y/lHvA0EOHuosjoUpm4a9k8aCr6i
uvXJNbf6XGjdIkQymtpGFMzGLOb4EVwo9Zbw66MBXbcZuG5vtYceBobHFrzmlf/wC99h8fOEhuaQ
bakXVT1KQaqAfdP8GdtAoVykbcyw4PqwywGMOqAHJMMvLJczdCxt/sAnDpYjBmAEFvExT3WoxhPF
mxzmw3YfcfRSB1adPrFsLwY7mGW+xbX/FY1Pc8AayEBdE8NWFJHHYyqlVu20l0AOcRGjg492s58P
dyVq7D/lPFm2XRJSF/h5+VVE93ecGGnoN6yQHAr2CRlfhpRnWPz8Vl95YbNUXiYHd05AwBS4viQu
NGI/5nczBdtWnDci2PnnwlnU+oW9xu/n/4ivQfsG87jgO0qoE020i6vDERaQAgtNkorVDfVmB9b+
decs7wVsh0tSlqp1GOd1rD+YA6WJdr9KHlju71aqjqAuJr00KrbOZbhaJ2F9VkFI3+hKcE4C1vqC
uRZMTlhsIKXkdV/7NvPcqI8f7jM+HrCHC4UT8t6Z9SAEWsQ/LCsJVysInOE6hIUTeGAdk2AlDq12
sYj/ZrzdlS/mhU/h0o+JRo/wqZioJHLNNyfJTx9BDS/8+h2oxXRzMMopvnp8Jqw/zwV5BI5Z1MrO
aGtnzMEpNP4quveOglyDpHNjZ+XURxh6/yrKttIIfIsSoE5eDXDfGnrBzRE+gtcPhNGNzoyCJkdY
1BQFdm5J0IuOt8mK/p8Qbk5B/gPZDDnXghmB5PjxPLuNOtM4WOaaNTX2u6B1PkqFkX24XryeOzi1
v6EOWp9ABK5a4qQoOmSMyoXuWugyVodSmcczqwdiawbRJh6RB+Xby4fuylBRNg0eM4Ssz3oNs5CM
FvCMJ3mybpJCIn5d9u+sLe+2LLVrEY3BZyTGygVcLYtvtRPiwVlto5ZhKx7psBBeFaxln7lm32yj
CiNq+EUX6hpEtCgHFvf0zgdw/v9VK6lv5ZJ9Dxgq3WvWV/xfG5eD42J8FsAPjWRuzE9gAk6F06SP
F+OQcho2t4ph7aPlMZtMeFWbcMnHDRShpZd21wNPjVnnQiUdpauPMsULiG3ieIqEyZj2g1JD65F6
NXT3w/qoyix/upJN2V0mw3Iq3lM/NkCZ2pa8Rh5kXE3a5tejGgrQ4edgIIYXWXejOvc5z+YdyPG6
CaJ1KCnHJqzKj42JEL0RbXuUndTyoP/dPuFC8EbVDA+HuECsCCikc4GIeChx1DShKPkRO1teAqIv
UEQewppA4ANDOGB06ffSQtH1v6nM5p0JGtwRe1UpE0ImO+IGpc3sNrLA8/cqkzlKEyjCNBDx5Zcq
wPzrIgLwPgePyQejTV5UvNzRt4nARc7OCAeWE2Q0+PJovJe8jgyp6sWLWZsy5Gi2EpQLXlQviXFX
MvKX9gBFgJeOVYNuaZfNHY/omiftzelp44GYUaG4x+nXlTUObKEw6bdQW7h0vDkoBnQA+zSDgjtt
4SvovL5LnSyAIDGEMBKciJx4zC7aqYZ34f0XxrZTOhJXzP42F6LquRRg2cFmt4ZJZrWhicEWLE25
KbLJxzLdvvA/KvoTdKu/HEz1GdWdLQ92XfjKWKcnYzvj6cQ5Kcpnhe/CHXvaB1P9qZU7AZcrS8Ad
L63Js6cegRVUoNaZ56R1/7nZl0uYdMbayl6qhH0MPHh3g3qty4ZtJoQbGPkoWmXvKXvmCU/iOqgv
rVqh399LgYZzfH0l3pXEyXCfTzViuKpB4sAonhTQQi2LHslCjEhGiSYevrgicbuv9U40flnis+0a
jBfdNvu0E0RcpnSodUyfU+3qH4cZTABm5A/JwCBOmGWrVdrOpC0bKTDz1dmntJ/QBvgCAVzv/k4f
7AYYUagKYy8OEatlVt0kfScoY+PHxhw0ZZD86k0qgU8a+SF2bkv21kmBYHpUkhXN1Ac+NmygCwB4
FfL/1q1CHZpM/uDE/kd6kT6BYvd7uwKiJG6C0EYijFBOFYvGYUSoGIbzVxga7CtXSPRcrSs7boey
pp/E0iuhuppEn847JY/OoYgXRHBZMesQU4ZyEO0iHKdDBjfdqRM6Uv+K4ggJjhI+QdQ7s/1AfZUX
suDb4BR2h3e87pDyFxmfdAgZOTNunTeZDGjD9KHpZeaTPyBfF/nI5kzSEnDklzctP+tbgv3sClZs
6Xn3vUrO7hH9apH1KjA39rY4nTQ+rJqtXACv9ucVdpY2zsHjUeFzyZee0p2Xsrs7wUXr2N2tnyRE
DDdJp0/L2XCY9Hp/D5pYJ561pNedvNoPiwwaZlSo2e/fqrdYPLi9EQq4PKS0EhDb5JoBt8iagJFj
uh6pmNeP5Zzd3NukQbkv4C9qlvU79mspt3a5/xKbauiGSc2tNUPyKtW6wi52PnEskDp9gV3wk5vm
Euklo7CpqSuxe+ylXMDoVLH7UEdcBWtKqM2T246XcRcYM/6/IiVJedpNazu5dNNKEPudy9XvUydP
ae0AMNoYaAmReGz6oD2t22p+eTVUW648pBrctsPVE3JKXXzAxvQizlhxdteK+agAtrSeVfK9EtK+
BOSOwqza4j3qu/wn2V94Bx724bkipptmkQchjMg3S1xskPX8+bWKccESxNeEvVyN7hWSjBJWkbTg
WqBX61C8DB7Xh3H9qHz8AmtfvYPuVnmmBBeJbuTdStXP3s7JeyB6FWeYfSsUGEz73DVJIwvQuFzW
xqDzdQy2OUdATUHoxIGyuZHxrMVb74ojAFAu9ACzLPZSlzPPOXOCRK07mfOobhU7BDG/xeTNefeZ
qpyrc55jiGla0kEx3xq4jFpUpfyDhIuj1Z6DUeVHp3/fUXyL+78TZwSgKkxzbt1oC/Mh6LjZhNck
PiSmalwZqAsUBSsLatC2zopfUaMg4WLEObr0tz+y61G7Yuh7ywHYmdUpRgIe17OaVefuRvXeIvcc
CGeEZ/KIGdpntz4NAZWHScw8yDValeojAWSpuiMBd5O75H665ndCeY1gW+PZFioMhKXPkgCApqBz
BS30vWKBVzOjmW4OrhqhhNySQS7bK23sO2bsR+OI4SMZKZnSu29IWAGzOJkjiE4ZVfY4VTrcMy2V
5dq/kF5caRfJwOTUzXs22SUWRA0Q1TkqXqeiv3Qjp33Q01KH0EJg6QyCfBQzrd5gdNPRxugUXeNw
Q0/d8enh+Ml2gpeuM4KP9nQVL2hWgUP7N31RkijTfJh27LgInUCeYfSQz8JLDe1xwlom4tGARmuq
B726bcq5BpYS0q/GESxrxolnHvPXwjAvK73lFt0lADU1ofr+59CpfnLs/dIRLOChk2w9WS/HiA0G
CtvPzBD+4sjLHWmRDq9FAe7jHIw7xkxnkK8rjeyGUCsKgpYrmfgQ3ojDzZIBAyewPduvpd8a01xa
zi6pyMAZM/y89YT/+c++6FYmBFg0c3vuJVOs10CYuMEKNR69NbQ7DfUns60rPqJkkTd3JDIidyKy
U71W9aM58KTZ2HRdLYc7K/pz2wPeWabjMqAh5R5BMQq2c0EfVkLm6Bev+M90+nWG+0T61A8z+3Tp
C4q3RxOFA4qEHTIqbbG/u3WfRVSEuSjEhXNC+kPUTSkAfnvnHccIRThc13D5mku2k+Oy7SWQ2XBf
WFn0VPGg5EFQMFr8kQ47T2emG4v7NONL3uz7MKNg7gsuy6coUHgybGHOwqaK+PQfRASTjiM1fWkg
Ivin4ri+GwSavMMIuu6u7GU3HVU/IEEQtHjRF1veCEPY0ZGoXfXWDqf5p3ayo92vRm6wM4auC9ki
/quh9l2lt1nlPP9VPo+4xmDx7CyWChrPyJ8p1Tpt7ycFgWk4HLLxHtRUXv6ZHuYl6iXLaTGkpvrg
scRBlF/1y1WObkXsP9J/HIko6VuooH0Zmex9LdxjzuhA+rgHNeU7Wsv0e5pyZfYJ6ECLk9HuAoQw
2wI+cWUrmRxQB9rQ9fa7qN9Y10SZoXuZe06r5OudbyGWvYVaZqaYt+6Ac5167JoGBg4Q1YHWCMGQ
siqUbsWJ7ZdCn9nPIOcSKoHQUsyJnVmV7Z/edc1qbwZRBjH0kwfyZ7sB0cBQVVFeo7FRu4Z3TPn9
vDykFF0o9JknqWjFtfnsf8ySZgizW7ydi9l42WlnE0naYgDhJvlSlogFP57m8uUlxRQeIA0pviIR
bYqSjGuxZoq4rqC5XmjRHHGLWxzk4ybqGMRpG6KwfX6570lUjp5d1jZ34sHg8pTd0I0msAzuIqPx
TBvbU9sxXhi6B0ebOAxHa4Z64KHGTymUnbxnhhc/YMNEV8zwy/MPsLgcFDklnMTA9OyzoosGyhFS
viG01EL4DeQle6QeN6pZbhIhTZzsl662twYbpB42HYAj5SeVx7WTKv0m2digg4tFne7aCMnlapQu
GVTqD45LlRf7z6lcD/Dpvc+gQ5rxxEqI0vpM6yRh7ti1dTVUj3jT6gDZF1YaGVg/OKPkuvInYw/p
esoxxrdL6xR32TYSnBDtBwoO9uvDEBzvxEwPbXEKM34U6muXW4T7uEMfnnrukNiPQi9SlnhBp8IO
JlTf7IFzj4Utu2f9ZRol2W58Lm5ffa2RxqQYdmff0e/JCU4RJ2wamzrMqoNgJY0v12T79qAC5E8l
wxKnZaHpQ7ZDD76Ve8sF70G18urfPIL8oldgGLkWmpHdXin1AvbqSBd0Qz7a3BTj03OVkcDBFK2l
G9ULW0uBaypNGYgtG7w2G5toxJg2MraGzMtRIwramxenVPsLokvP9bCyGY0M0eFWfLBQF5wrJmAA
tX8MP6p0H6pBbJrQrMzzykTMeLWJODxC0osJv7MznixKJ62BJriw8ELur49eCgbOlfHEv6sF8pLv
VRO7HQKcjgiz+OQR6iV23TvbTZnf0Co8cHmeOa695HOP33lRoGRCVASJZzutijBHZBltgREYhNYT
meoYfMtyRKuwf3T82lQ7RxlOTki/Q1N/QDYJ21DHj96f8jzbvqdpb3KmLVWAq7oB+5CFMRYbprUg
XpnhVp0Lm17xn0LYYnBCc2P0KVpBf3fVe2IhXzojNaIddqZ+rzOYyg1lVGAwq6I6OqVVNAWlWczi
BdSgLUuf8GLVjMmp5glUXldO8/hZVj62UbU1gQxopsxyMHRxSikR4WH0cJCVZFc4lFReLtFLdvx2
aqM3tFHWx3RDysRfMKWdcOZQXlNb+1s8eT4A2Ch7xyljjnnF3dr3xsG3+snV2N2f3QnyCxNUgRAO
RyIIJo9jPiH5ahqr6hOugtgpLe0loh8PyRw202VCXXCWuQ3Sm5q2c2zNjKkTNrNCe3LWH5oiM4d+
wuBPlZmRMRra6u6rGhohRC8SU0xmLxaVvfwWxrqrdiOtkw2N/jfEfYfDFjw5gov5L/QzA3Q4z+7i
xAifgakz4Luv1aipShMLMPToC0FRpeoxss9/WuSL9pDzWdbK3UMoIo8GH/iufb4StibYpq8HBgld
eAfzUHL6XdpAj+uAlDx+cYaYjSMLT2l0Dd2VaJcQkvb24Xn1AqxQy0M8LSwJ/PHjgIVy1avUQf0I
UFuvTjl/opSkeTordJhRyejKrMefQsJdcfsshO+LYN7IUj0NKRv8F1YbfI+6j5QGElSpBvDckTFU
qYP+SNJN8DEcQ0iRWdQa63EFtncHjGJUXwhkgwmoeoQ/CHT5NffcxXjvVwOw+BPY3ozGCD76POvi
VzNy6eRbQTXHlILlgcQuIBTcQEa91dDqyqnZJ4KYjE+YCJMJ55tOlNGW86AsRPuEBfBw+rEJMVNY
i4PFoukR0pFcJRu53O5cqif/ZDvoM016wkqhKkiwzcVnOUUITCylLg9w1mdAuhsGVXbppGVplcRs
akUPa8UA1mqYKloa9mP8XcGkgc/1YJlh6q9piOgbFkwaitajfK8DVfcpaqZHggB0WsefFd5JbnRH
SkWh2+wSLD9sqO8p3X3v9tO8CKYdhCUNUZJLd5o0iBXSkwBebJeoq+yZ0cUqL7yrE1TGECJA5NS7
WOJcmb0vuxyG21egep88d1IkpSbIVqyrKJUwUZ1kUnrdPD+jQfna+wCrqhFnIpHTFefMBlcjVS8q
0Zed8nbMcoluTJDwikcFa0aazaMhpMQ/2ScMGjdATkk/jbOiADcIyo0pVs9leZaQ+G3L33k7UL/3
u78vlNHLrDp4mwVBk7VFXec60LVekt+/DhPxjpbVWP5M8SDC1HAphK8x6PRwJvWLuaQGdu849K9G
QCcyfCXq6yZqGi2I9OGaPSKT0gymqm6E2jqA+/QWmgthlUDXX5RY59ajB6GRTI4JFPkUO9FuJcZj
NHn7dEiJoSZg+UItl8449RcpoZC/xvW35LTbMYljRHkD5TeLF0bXTT/6IAbdlHruxT6HYaM8ShHI
u2eWD2ZjJXVuWBCGNd424eJGVHNjZ0cQnPahDD0ZM2qWW9+5GA+81MWdF55PNR+0z+5hhbR9p28X
ksCUoHwxUQszBrFV4XZbH2Y+wIIfgmIEOgScnfTFZFTAp22+JY6oi2V4XeuWldHP3947w5eWRry+
5JXIAFf0H2AhGPT0MoPirZULhd7lG30El7zX/QWS1Ugs4wmv08YzHNQeF9EqxrZXmnYmafFtSeFU
ZwqJTpzOn4/xFS9mSCeUk/5CcObJYMvo6lpQxoaoviXJ9noq0cN01pF348x388vXddPALQttmBAU
wT94RaypihsYKVmf7AWdTUk6LvvSHkARoVG5K43QsNEn1FWuJtos6/Q7OKSwVOh3mhlNAIgx6GO3
xG+fJTwVmkHvgtMu+so+rCJbam005SXXq+iSwyOviCp4kCuhiJg4fNZEN26/Y4isEOAumAEKYn5F
fYgo7Me3OBtiJ27APJ6Yi6TVXtLlhd2arYCMlkYtE4CJ+KrKq5o5fNcZ2/xS7/ZGM8o3Pb88VVhi
e7Kuigr6BbfzJWZmmVP9mAw4Ee6EKDho7fS4jwPtvBwgyZ6z8Ebi2pTFyAdoVNkS+coly43/ARSh
svgF2S/G9gYCPk+TnfmrQ4Mcr9+nv1YI/7+639ufzZvRGHIdlI0l3NVifMnvd5E5C37heAilZZPA
5bYgZVvFVGK+3Gbe5hQpbyKmRJhHuDdfvwsSk/Oxi8uxSll/kDNOi1ic1tWJzaUF+swaTNHW0rCR
6RoTh4gm3pd4lIXZDxz8c0IY9OrB3/W/eEPttxXWe4CG8FgEM2+0HAFEXpKJ8W9jFnn3cjYNPxOr
P4c0mKY1xeFQajJLvviJKEZS+GSzw3lPOvWj4e1jEaHOfcMGoPmObEmXuGH4Ek3LRKmhbKVRAO58
Bkg80h9sSwYb625TBpesT/QLAFsujD31LO9nflSMU98yZOjn/FPXksuF2BjSiI32z/DJtjQYbg/f
qbGj+6+GDTDymFz3ArLqipJ2n/Aq4Y0uTBrzNeYPszsbXq9dDiZ/DwDjJbbDAcULWcNiKd3p48Im
zJEK2YtQxJBsOkFOX8NfZZJ0feHiI6i/qQWIAVj2yHU86Q0UsAtx+S/7r2KlHVHe3mGtVZqRDWx/
asurcJgm9GzW2qxj2PHOmBK+qBkBHaDxR18256tlrW5OIDBPuQLxlepLSEpNE1XgvpsehhVCZAMZ
FYup+hmKP+Wci58WnuVJ3TYZQrdygqPivGR0DN/B4AlSJdoXhpLLhAyGX7l1ggStD2XMqO6L5LDB
FXtoe1AHA3H8c4N8z3xW5JxQmhj+RDSfneiVz/AeKpFwjkTOkRZi8FRMhylj/fqcyXt1h9a2B/hO
OQhmsAGXrJ0RF5v8BmJ0m51JaMC3SrQbcxJy3jT+7eAByQsIQfO6VT7f3NqBmuZTbBEpRaEzCEwS
/Q4zYZmAzz7NBfR6+3x4KXjmYY95RadC2VD/yF7Qhlcps683CnmiAz+Qw84KbewU74T1RUiOpnKS
pmli4jLtMt2cUGp0/FfFWr5O42EG3a4lafFH49btFGJ73NyGSQN3RJkkAIOETFUqV6GjR2tunRbB
5HBJwhmtmB0l6JAQ5/WdPQTvjrqsuGn4JZWtp36oj2ONBZY9/8oOMatFxwIDtJPNXWxfhlLYzMP0
dHzR8cvLKBbiOSKcqDPFq+4xHkaAdyp1YH+wFelSAnigsEqbXyfcwNu5DpRVJMZhG2SvRCwkVddm
6drFJ+yhLBkznmVZFjk+vCWMKH9N5W3NOpENIyJzf7LxFqP404aViMSeaxLVIcogKtyDr2JxZwFj
QEP2B9Hdl7Fq9lZ+8/1l+S6SE/TVRaq0m4Nr+i2vbqLp0NXi78BRNh+cKesjHV6Sutx17ypU1uCy
VkX+23yYcPI4p+z+EkInpGm0kAA4nJvM9LF+7p5WICk/0Kot4fgTThFvnjGr4m7kST1tThHBF3Mc
n8oywSRWyysJwbC11ehtqwLNvXg97XNdDrHhD0/O51+nX7gSCtgvkemOOuER30PHDM3MvO2fMwp8
IUNWHmWy2itfcprFOosvDj/fn8rht47qtD/ej9YGs80MRVJkZwkQu0If3bWS5wCdcu1M5+NkcsVf
r3oRQueUjzHqZl7K/q5F3+KI8hDDmAkiAuFPERol7s4wmrVML4whhw9Fc3MKgWhxtsK1ISY+7RBg
G+s4OFW8F/1UhBPPH/L9eraUSae1V562Q+JanX+y4GUSE+GKfVlMOisKTy6TozctEirXEhJLRljO
J5hlyLfumxn7CEfvxPjoUUTcOB8kHZLtK30X2PB+BaZ1AOBo3T8TdPszWQGz0fMQuI3dOiqoz7A6
JqIfAjqkEy0+abQNhLrMTdjHTzBFFe/JUYQ6+USIm9XCoKvyg1vPxs2vRwS5M8tvZsypTjYnh63/
A5dV+uowxF48ciiZtG1m1j/PuYO4NbqnEWEBlAObZqf7ntei8CuF/jn0tHLNy8I7IeZEsegVMEGt
EfZM+X5DnhMvP4tYAFoZFAlY42+YP8CUcqJ93sawbtNoYWO5FHvNg7jVCeEraKK/3W9X8UPEiwYF
FgxWBeuDOyvodfK7UvctSlGTv9apKb8iDZpXi0vWIRT0yQrfw9pytZ/G0k9vfGC3Wz5SxC7bM0TH
D4Uz3fDc4Y9Nz3oHdFgSrht3IdnrT/J/lFdllZHy3cUnLKM5fuyVCGd9aV/feLbWzGp1J2ew2dKv
cc/i/r/RffnLqWqGkXsESRtQcpAvb+7wHT/hKPFfd+UmST07mRr/kWs6VVp5C2ZE3ITl1Gkiiun1
T4MvvEgN7hRNlquQHWcee4w2Q3hw/g8Ch5ozVT6Hvyt9blUPxqYteKVDIml6Tw7ynqrc0SpHbxAA
cVlZBRino5Wr/D2OjQS8btdyL1pyVA3VZ/wnFJ49tFrsSquY1mzqcQJRLdZTH6Ya3/05ZOHqqsyV
2tzoNgPI8v4KvFO2hUpfeSFmgnSRiGojYl5ym4Dy9MXU7M1bdlxlPmuK9OkACndoiIwPmVF01Dgp
6DjhMTdhv8fmlL27hVK0edZP3OFafZmmXiClj5ubEW3w7ALQ8t+o8z+INsrdANy5nZR7c791ZXKw
fPxtbIQOeV7JeSTjLyaoB5fAOqU48NJudzMSRj91J3H5lZQ1aDpMwA3KcXjcCB/upmBsfNHwTjkC
0DMyY2IISNFn6x1Euz9WXAG2P9uqFizawzRhMw5CyroNWTnWp/g9mMBIvYGCEphBgwEa0BGUJUlV
YwTQ7fe/AosFoMaBT4pq4ZyvCMrP5onXq5KNxpHK9V4/zElJX4qDU7gY825PVUsrHEh7y68g6iA8
XW2BBOfSnZft0yIdSj+x64fNCI9/MKal4KylnflXS/sHVVWQp7I8IHEAFXKqiYgMVSyAzD/Sw87N
bpLZsZUy/cCSZftwmsJsP7eIUXqloGDaKDfSAUH1vpp3o00iQBHTRs0QGrkNEtYn8T48h0P4m8cN
t5iPGbAu95euSW3EFk8962YjJixW1Cdc7cmV22xKm4wiFlD2cKgYy7Phb5WaQKa4dnIF0vEjT84V
cii+0xZ8IL8NpL1F3A0VhLa+ZMqEtn8JzTm0poycjM8E6rTyIbQv0jy2TqKMGhyzUGDCbqSS2nFO
pouxlpDBjK/G12Itwd6JivNXt+pOkHZq1ljfr5FzZHvFagXs+pmzxBUGfQaBNjrwqZ9uQeuBYQQr
SzlE6TTJOKx+EgLsZU664dfmIvJn3AdM3wVtQxuLAyLnvy1TH1+5cCO+SZqI4XBEnMvHwGEJRX+3
9Wqgjj+zHm2xyuBg4OYikiuKHssc1XbsfxQ1CyIQyuEV4feh7O47hpvj7Yt0FyuQFjm5+0CCF6sp
RyvMX0YXHODe6kNc4sQaFf84dQPOR0uhc5rfjHYr86lng+3tfSFcKFKC9L7UVWQNHyWX1J17wPMq
BlGBkVGmAKBQlE6FxDZXj0zQDw1/UAQDr6mlRDV8zi7AWD6xzBWvtJo0pFvX4r9/CkHPxSAY3BCM
uG1ej9toWSSu/V0mdV7ompCt0cNsRRA0oEOTOKdI8Qaqa0QG8lfja157y5iLf1iLmPaTFJxSeGw9
KFiRQqDmJFqV7XIJSH+iZ8wPTvLgjEf3AFpK6EAUgEZG6wnAQkuxnPZ6WrdrdWfp7CLUBo/u4z7u
A3JAo9Gh7ePaDASHHjxiowRE/JSW04/iqBWBmCcsz4cu+KNtufngiCQxmivj3jnnQQLSEJYnzA6G
MYjm8SLpeyB3WrwZnBDS+VLopvgmnMw24DLOE6xBNyulKRJ4P887H8PmDgbyG55DWVjC+HK7+Oof
gIGj3bU6gRyvdJ+0FLGuVgDQaLfbnkzEC7tj94Y7O+iD9GGLbCp+/s7fFC6wZK2uurd2NZhcNpqK
QCQ7IEyyZNUNODOQrM3Vct6aTcN6dVr+CHaDvsWYoq0DJ5/VU8pkuzuTFe89pVHpE7fmF0dKszfc
MThD9PiTCRmEHKa/YlGK2+UjL60/cuoOllpWxBW7Iw74Njn/x7RLhKlubhqxpEr6xyiveWYdM24a
N2VYVEKtzuiXjA4oEOlqkc6nmO1TztSCzQ1eoKL1lAJMYu5RKlbYPgydHv3eHEPD0+x/cKSPkfWz
rTAOS246B9HEqK2asFRshWP8MDh7J0nFu8IHshvbA9hdiQOMo7wOtHNkm4dIFkc+hVgmFurG5anU
Wz0brehSONgdIT/OxdyemO7dGJsFcmeq/ANY09U61iLVOOvGS8tKLQW7fdkpBMXNw6GSKzXZk1mr
xo2q/go1lxJhZhAE1TRtGZBUMcV4wECMJ7GNq1Si4ljBTkkMfH/0OKg5fVCA+bzu1nBJvg6o4zBB
VT64+6tAQsKbGWLU5ubkWVBZfH0JufghZUtktuXVwnfEqR31whpXq6DfZK4Y0NOLvwAS5aNPgY8u
VQ82ILR3Xdv0FPDqmb8UCKKtBNK6jOVMJEbqeMivn7mcSYylELVMSZ5rXSOlNg6vcpbxkD2pYdUr
wCqPraAfq4ZGAdmOOWdDYLCfFQcKuIhoD7694kphWisbJ4fNCt9Bn0b7VoT+gOAkIRULTxWdvw5T
thvEq6f2kaKLoBQeo7pfHDHlp1rK+MtqKZ03jJ3Ceu7J1kTyZndIiy4ubw2mL+t++22p4/wNfEm7
sAdomsg+7SxnDbfh0XzygeSY4KYrEB/J8p6hlCdWhBc86N7wrKMgEOvnHMOUwbasD05C4y9SQs46
1Pc/oTQ4AcEWop8By4yyOgsF9X7e6RvCkyQEqP6ueXDi7AA+5Q6iy1jBEuYDkMld5WmFBZcluC2y
t28GbL9hwLgDkZe3NQKaT+C7gtyiL6UWz1sZKywLL2XM2cvC6eI93OSGlxdrzIsxNPteb0J5Oogb
3O4QkDCaz37FIOq96dUzJxNXz4kVV2LtVsibaczwFPl+q3GQ1YHhI2KA2TtQ2aepIftOk15Jp+E5
Eprg2Yg6JcxrTCeLGF5p+t8ZCj50zjBnTm0b96vp+90bKc8GhTxYshhn2wNPCJ65oBBmFb5GFltT
qmL1lkiCCgFFYqeo0N0msYMT3wu/98M1GtIbDpeesm8Aw/trH3tW1zAnr7viu3dAAcQBRD4YHRxt
YZmveFIWb4NwwUpylGpaQ4eKNnjlJ9su3FuUJ2Un7KmWAqF6LQOYUwU3htzAs042dQewAbMA5LZT
ZySdm48EmhyNv3T+l/rNMzTuOGMG65rYODkDmrznueLtaNZeSoUIgr+CvQaSNfFea6XVshfQZSOA
Xk01OJkg8hTWMEQhOMwhftEDfNF6Jbjz9sC4kaF07zrAXat97adxcTKLeE8nNDu/+JrjPRJK48gO
1NEzjZWg+VG8HbCiGLA24NQKYGQ1DSLtdQBYV9XO+EjY47fe1EthNV+YvGNWap5DQzxvJYWC+A62
kTULBFh7E7JU5Z5GTRlt4ws6abSNr958fF8H7lzlWTG3Mhh2Cj6k3IOAQrhJ6VQWuHSqF14+fzMb
4BLF8TZczcvNc8EOFLPRZAuDsxXJGKqTdMetNEpMUyQi3vldK+rG7lReOvDL3Au8zu5E9/qGqkTt
A+2UKTtkeESBBj4/XMU8JZW4a4KW6Jnv3Wxx6TlZb5Y9ih4Tix5HF6HMAZ6oXLKFznJGMKxhmNBm
rhbP7nZc5b1BKIeRSSELKKsh9A3dhgyZNQDMX4zZSue+o1KXgdO8kaG/K6PpSWUN6hcCUQxVCweG
mFqz0qFMA5LHNiz+K0S33wo79+eRDK02dEf64Saxlnp/522ONPsl7yExSfN7iVaUsDOt+3RqUFz0
EC9tWtP/MKdSLYz4JuIwnXH44gw1ilzcsmRuoe1kh85VSXZ24GrpJXMjhREFNt6jVybevpE/5HY4
ydyKQgm4i/Og53/EnHC6BZ0vul3CV67dEcR4mHSjo+1HaAzfoIis/nuoFiR8pj3ce3bfS66i36V7
PvzSZTM6Vvp6ESsjm/H1E1E51PzV/gTr+rIXrKkFleiOTcqkk1HiIMp14yn0E0qiUNRTnEJvuoNr
q6Qwl4Q9tVF9AouQGa3PVJFeEfO3Ah23TQhQbgUbsGBfPkcSZqXr81dJ/taQGlBk6G/r6LnR6hNT
ka4bQsux0Y0MxsSLbkCVbeqJv39xGz5zAQeGPAsy+ExPJmJzigPfI6XJJMJ+Xsvni44ij7gls8iH
ovTtlhw8DKTmdUmuSLsoj2sWykRliWk1jGenaOcSBZkgFWHBShvMI9EwTZRLlZiB2tnyvTQKfsAk
4LGMERP/Nr0zPiNwcZXBmuPwJGNjYKZHqFG9b/L/SSBgg0absxV+xadtmrXf8qNbZbKszwBdmpkt
CP0zTHAGGWP3H5j86Yep/rvwdjaWUAp+ZHYVCry61sc2Q+SQA4rlOsSnimCSkF3gQ3kLCM6j46Zi
YMlfBlC6w6nVy0EjLwVJEuPrasBRRsnw225W2So3dnXU1reIRMLY5t804vFUNMe5iMmFJjKR2HDK
UKl6ueB8crovsGx2nOKvgNhaTLj7TIjJP50GfUf0hKf1NFyhu65npTBN985ZpDmK+vrOK87q73UM
mRjXhMhgnm4u2V3I2eKEh+EKo07uL1/gdl7SA5oYg0qklTDVzUaJTKUnL7Kh7+iJv/6cN5A/U3zp
StLHl8VuvdA+RqaW+b8HtGdr4l/UhPn35xW5Q1EVq1x61Eflj3rBuMzdymdxPNlH3UlfaTzGVXoh
y+Sjr+jJibvcUNlUEcazNd2tsDHVS1C0kXngM/axThFYFHQ3EXOV1D4boRx9zD2fRjYMYmU07Vmh
1gDRpQo2kE1E0zcu9BRhroRIwj2cUX3vfpi9vElcACUTuvFtFskbYzSyn38wLnJGXHVUjxbF4/yk
SAuFRmz6JcabX/NeyCgqynNz+iPfG2wqQi1024ltkz66lh+2cviWPgJZOppEFApcNyFsH5tVW4qM
mAXuAXpreOJXKQpVl3RPuF8K/y8OAEeYdd9lb4OACazHTKg0MMVWKo+/DI42C9Uv9EqcepgTRieu
0nsBerKIITC9XAplVXy/HPSSzS045SQ9Kuee1+Jexac5+5qd8zICXaN2vueYRb0X4i1eBMtCuhaa
2pYw5F3mIfh/fK5HoYl7oQJvKbpo7/n3z995JjHEFm2Npm/jNDHoak30+/0u+fxFjQ48YXA4IctJ
dHT/lbjvJSMBi3hjp7O2OZ2WL9WIDDLpHXnAHudUKAeQSw6+Iw1z9vJtnJ9woObGWJkjm9xuTJY6
GQzKRwDofa4/NnDTcuyTYby6S7bGnJ1kiM+Wnq5k+qZT/sIkVPt/PwdHnjWlxcrm+1EKV4wWDasd
zNMVumJ7rYtYiiLQHvHgDaRMObGZ0lrjbPzZ065YQHWbMJKDoJf397/Rzh939zmOuGVFekZ2pTWL
oEDfLqyH3nk7srcxthP8EibGN4k4qO1PUuV3EehyurA0MDEr6JldJcF1QEay3EWPuk4HWuIJC4Rw
kpDlZfDsn+n5gw3QUqS19ypJBTIf8NZofkRjxWnTK+rFLCpzpf4QaNYGO9T5oHnTKEx1ykHSeJiw
EBBLUD/3O8v0XVeTVZuzP8G7aZKuPTO7qM6C+INI3Z00mr9swkudZ8b3s2v1SAYAh7fjxfgSZHTw
tMkvtJkYFcgByJ3S0RRtHc6ulGIt2hHhzju2fIo0GZmlNcYJi4KCdbWq2nF2obpxvw8OW52DNxp+
d65opmHTwDXOwPq29AZTYhc37AxBSj0AEazG2aNgCYEzZELDLwsbfvsDRai9J6/MnPv5yERxK4KO
XbW05PxrsSPMzRspSyHK6XaB9BZjpkTWjctbi1oU1s5IBkJdLmDFdHECYuSL5nRp260yFUs/FkeF
b7oDWDYvSoMnCJDT7sZESiB5s5x8Ului0jCJNiyIy8nijHzYRNLnmT6HKbRvraLwKdtC/qDTDmyA
4eHXpzjKcDWNuJ/8qnlqoGtbVQwT/gY3vxyjZUQ4q7iTaD9lrJZxZR7qGiiCshAVLXpW7y90k1pN
pNz07VaqOuLNOVUZsfrpoLBh3DRZDkViR4G8xPKDzp2qLHH4aU4k/+J8DCIdnQtCpOzg6qtWb+mp
cnxQ4LViqxlmp+1VDMqbe1O5i8xWnYbXQ9PqnhcIEeZLSN6sjDr28/GlRs1SL5rzByJruXFlBUX2
+5N656UhoU2UZh6iaVQQ2FLiTJbDR/doShGDgRdInfpveaL04qHu6p7AvdZALAvsYVpyVB291BSN
SEN+TiH9AGOFnBd3kMYNLKZVdcO6YJdS+22BbUCRfOzblZuqJpHCL9kZV8omLkE6wqymp7slOqyi
EjO86AouBdpXQTry1huJgJWmsB/dVJtKzFXT3P5Pp+Kegna+cUj/Cg1AiZgW4IIYDCRfIWhmgQw6
biXdl51++my6G+tjzDGRKED5r2lI2lazmxdJLr7eNx9mJRQ1YnCUH7QPZK0oC4SofEhLDVjAFVDp
fiWtG+rNOQWtGo4pJvURrhGqWA+RlEfKXvdDpJ7dh2WmligdYgsCbTiZRCzSPG+nB25QIcZU6ZGQ
aGjzrD2+z8ju5RYpRyTuQl+mIOHnhcxgk5sN3414SIaRUhwNtRmEiyAdEZWiZI2K8lPgkQvl95si
tdcb18W4k/mDeBzjUPzNk0pgbkvRYMtid0OLtHPP0145jYiDSgF9/buqG351mhR2/YYL0itHIyOm
FcS4YzDVz34tR1wN181Qqhon1UR7wv9VlZZJsKGEQJeqiRctG0Ha4ERp5pnmLrYkbnVo9iGmzExb
VvA5RY3ybgta0X2u2Ii6oRZ8vy5jaZMMgAzWPC/8h/kZzOzWlwKOEQzah/UDbVUeH5B8EkiL/qtb
4c/dhCIUIdcu8SUy5dBv89gHtj1Eqpk/9U21yjtonzYAKUA2D3O/yoVCfhkkmH2wivtQB24as7wo
KRW+fDfTGCXPhg1R6kgjov4HGYblgxZQ00/2CXS/IzB1/ydoe97g0BCXDN+aRsWQD76PqbHTN9wK
216EeSmJfd/j7ZK04zrdaOGzYmIV8KqbJL4jRu6DDCwWxuuhdK8fnHpj7u7x6zPjKcREyLZyRUec
+rJsq4+DzktDo7Hmcd+3Ask1Ys/akSwcK3zLHD6Dy80+/sQI7OgFQCnurAfOX2rkeFemePkxTpwe
cjxPD5Ec3qNgxrXCtvG71hb9DN3JflYDI9NKYdIx086rnChEs+BAItiuDDKW1WSdhsdw9uKnlkRY
ZkypM+CBM6hSNj7VaPuo19RzIJvCm/m6LAS7+KuyZyCUs5/Tem8bVXULu+QD5GCE7KOy3eBJxNe0
rl/G8nqzugtiYCqWOBGv/k9zpwve/sZJumDwWsAwa02udN34kccEaG4T7RzWzHLD2QnXbYyEtoow
NhqaMbPDSMM+XEXgfKpgQxN+oRrgZwNikR5Bl+B77XdnvjVQT5UwPls5XvOt22AaEzvKkwK4pqxm
+9rw1Fd+z9N5IJkkyLAd3cRd7uDQlpal051Cb+MgUD0WLpNkljRSwMxOiI0tf21iNA+pSRSCOh/w
g30ADxLXERC7MPIB4YI2GXH96ySPsjhTwZsB3pR2LN9HgnvwQGNVLnueUPt2BdB/bGUvWjVriyuu
UbrmZIvxkSPA+T4H5nL0MD5seatLY57Nzlan2owF/0M3aFiCOfVTXtdz900iQ2qdRv8ZwTzu8rae
BqxZznNJ1DURaK8KtHTT8A5PPfkMsF83FQp+O2fVzOv/opOj6Ff+kBhmKvdNh2HChWaV+rGQ2Ixr
77ReSNPBO4asXfSW9g/VURSXJb137hvLpd+Zzrg2ttj39TlDMar8zmlGwNXfrMi/EPn9aeqCKRw0
aS4ziKv0JmzLsajj3TDlQz5jXv9CKEShLmRk5q0prW6NlPQFXTmmPXwZQWoeLDr865srfphXZUgj
KXjcUsC0pDtWXNwiQzDvXnjcszgBzumWAPOvGRV11zdOSjOlA9xfidG6S0emj31mC5UTMeIu8BxF
7txnny4aoQ66YnwL5h9H0f1gZSlnQmA+5YMpguRiyj+6HT0mklvN0mCvEPPWjR92qWGIt3/1N5X9
iNKm3Xt7vOIlnQ/zaLn5LNfwglGbjRDbmYkm89hmf7q2lXutZazmZoC8QMFXOk5PG/4DBWuh/g6P
zu3cnAhD19UNFuBfPYP8NW2X7lfTrtDd3jfCjI6C3lEBvr9PBIwX/hUhHJr1RWKHES37k+ks8STj
/GVu6/sXiiRecAjPKR+CtCJYyFZr7oMTmPAyb0kD0+iTEYDOGrl3w82GxQNyIgigjC32Kd0ri9M/
fTAlczVjAVfP1XvWjry9N/yqfUnxpHvtIZMOpuN16PR3ws6ASFhwNTRvDQt1dVYC6Iu5IC5ECLAP
NB149jRO7rAOBMVVE3ZEB02i2hHREyCqzd/hZrIu+m6G0bCDl7ZEmq6MaZjeaxhYyc1KJACdyGAF
T/OJKXMwCe9V8GUvvzRXjqKCslCoetmha2kS7diRm0z2R6FImbf+FtUz2t3XdwtyEKvHJGH8hhKx
QM2L7l3G/y5oLLa2N01gRbWVQbZ8+sX5LSdm9XMyxzhkIJcjFqq1Yu7wYug9BrfDrUKgMIAGnN1x
deGO5dFsMfadyzlzG5zcU/LZkJzM+R8IPB7kTEgv06oTuDN6X1eKt7+7vJx1vQY8HvdOqbgu3RI/
7hGUkM/4ZEsacUfil5yiXUb1I1B5v0IDPHUOEXmXVzJP9kkTjPtrJ4hVqRG1LBL7N5NRAdcPQepU
aJS8tDQlSg5ysVHO6zPhrlti1jOGIk944Ij8621KDGbu+PW5GrX75bJiDuUgNgp2wFCUh2l+YhT7
wr77JPC59jdCJ/89a4SivVYjuCHaiddgc9Kiavz+CqLpveCUVkPhmRJZa4SVpDZfcwkNONCSgCDQ
4SV6x2eaZZNktxasy2wIFhV8Dg2VANpbnm/yrVAVAWflBi/Ed13NbrY7vFY6rPbPHwXSNp1LxUvY
ECfTGu25PWBzH7N7sUX+rMF/7D7WpvpHAuoUkBAO9b1HKKkUt8z9AgDwdG33oBvCzkT3IrJj24Lk
zepeoEmQfKqJR/IC/JGM5OpM0XvZ0KTLPC1tsVTs/5Xwi/vhJ3DtLdnVCe8pbkDes6EvltQ382nL
iOy6iyLWYRMErrP+VS7Ru6ogacfjZZS1b0dIaweG8XwbAEaKCYRh75q/cqRamYVMWpFAC0WCMHCr
xksoqUw9QwLSvj2ek9QImGYPRPeqgZmYMEBD467rh5zZv+3MxgmwYelS6qSr4oNUzsY8g07CTS5f
JS28oZfH4BPqZW/wfpLl0LwJDLU8nJZpUJ/VimBLUpfQGMowWLH/CDHgNNpekAAMAnktl+03unav
Xlg3mSm+cw4AlDJyR9l3pwTptt1jESHiyrIEcJW7RDNS05/LeLxiMxJxjLBF8/S3hyRaskZ6W2NV
WcU9gmDHb3gLNs9iM86tFk9tidD+quw6yvbfFT8IIZvJ59drqGsaXecgZQMtjdj/Do0EpdYelkdH
y0QAFsCn+OPLASOhfWmuAJ9XVamb65bWuhDL9Cys0F/cF5BWInuKfgveBF6qWcKX8Nx+NPfeVgx2
O8ygOwrVj5xZWqfK5VqmEPE2GxjLOtUvzhoHkmsCvUuxc3lIyAie88H9r7MdJmgxYT3KxMGN9g4+
ObZ9K9aRTUpo3TUXKIs7VD3nOQD1O+jovGzU2RI+udSRCFyHe2my2pSX7zItbdgrmMC9PQuhVJoL
MiTNI8rGI3U/yBkJ++G/E2nzQCpDLnc+mpsdLYPD/N0u6QCI+LHOsOjWwBrn+ULVKu7u3y/BXJwK
pZNMuv5ihTgJJBwOwCDzbhdvpywtONyTUdS0n1DcWvZXsbVklqOF4B5Xx5ZnVzmqVwC52lZBepSN
YTL6+quokhsqzW0fVXkJSM9C5dVChfbwLZxmvd3ZKghrJ19hcdZ3ROm/QazKIFfao+9Oc5LXMNjX
bVfQXntUxi5bO4gwIwnBoQ2qoYBNaan9auZte8kDcDw/NkUKWMWo+YMSJuFra0zkX6USzC7lMvrL
dG3hOdSgn5MiEySCLoFk6KSipWGutAp5xtx6iGiTMDGVvYyWuLF7cR7cfT6WAQ/h6MIN4IknV4Xk
D1sRkdFxmnfeS6lu7aaTqdZ7diCkHowy+fcTyhlzKE78F7ni4nslkl0syL1V1EzxhjbNqhuff26p
oyR9gjVC86XK6Cd8ANSk/ufOFxkIvCg9NCwfp6gXBI60XpINeXEGAuzfEt4IWetOvNhEWhN9TImA
LusguIfA56fvEjTrCQhM5ztUK3pXVe9+GGRtc3y20yDR63tjEdGPNEzvcPDJr421sXlm1679FxQC
58+34bVAa/C5ohNF5q6SR8rnoI4RuxdCJ/XnctufuXwR6ggOn3uDp/jzF/LDYTdoIv7IpUe1qjeF
Y829lrhibEq6gV99lliyTkrizHpzBo0U/75ruXTXHt6LOB3xtyjtiBOoW8i8eB5/NAk77BCx3fGU
EKNZWKl1EKd9jA4SGnyQt4LraGflE8pk8piOZVuK/c0P7UJk9RX/52sWaV1GzxYcFdqNaYU7v6m9
ChRCbMhly/9qjar1T+YeW2tB376zJ07MAnoH5XxuepsMrpkGBRYno0/deg9IZRbNpNq8YzZKZJfS
BCwsWqzJO6YXg5qOuD24gkmuQU+xI7PgBfzkQUb+rPv4CRHqRMH/Nt2Wng8Dj1akyPsj/E6eFsKF
UFQIa+m1ZAaoxOPDh4bnSMt6HunW1FWOqYFnAVRngIAuw9TnqZ5d8dVhXn/DO1kcsxYIBk4UFIj+
+oUU4NRv68jkWdC7rAKlPrRyg3IUi8+Gp3pcFzLSNocvKssGS16ibsSQ1xLWsgmXiyZRejShTvpx
OcL9ZQ2ZSkXfe30ttjINsTlQzSjIyFzTO73+nQM32QBzhfITfstL+cL40trEo2982ZNGAMQBEUS0
QumdC3KJJGQB3MH4D3HWl8JnSEd4yvL4JygUfX9q8xw0z6kKa2XibBhiggcqxt29KUDrK8LJj0Ww
t5f5OhT2HK6QFtxUzJ9zlnd+9xe2K7wJ4feh742mSYeGFS2HJ1HHNSFiANqvURSwl3nxyTRHhhYD
IxZYPCvnNQg4oX4ld41hRtMsy9/7w9NjdZnv5PUgBdEYebvSgm8UZuMazhpqZdodFm1CR3GIXc+F
OD6iD1LBWPRZgYZsbHhO9qMzL+UP7pZJA/KYNXyu4TsLgqOOCNxBw/O2tqCjKp2jePDE/eLmSPZu
xdn//PUFzAknKWhze/1FS3W1u3eE1ucafFyJ12+thO/imdVyB0vzxosPgYpjyTFMp2bFH8wpD/Uy
QahIPkJY1+608NN0PY1dDJA+o7j7ozu2QbvWwbpf2paPeKWkx9UlEoSTdWUsS+DU7Ifr06mRT56m
Q19ANOsHaEy3M2U8PM51IqDaZjVuQ5qT87lMMsgzLa5oWE4llmFsS7SAyxlS0v9inLXbHjwpIP5S
HOLjiCSeYR3WutbHxvfPxu1R5ZofZvI5+OP+w/lkLdM0M8yw+Pv1au5vAgXJrQ6RfXzNhSH821mg
WsH6oxxTq9m/kncHhHxJMAYOnkiD8+qH5NHJuLL6mM4k0GRu4bLl/cbUmN2bKdQ6eOGe7al67Slk
JTnd+UC64mn4vo18QZct7c04Wfk5/VJbLcNG3+2/qe/iDoJLUWfjNTDUU+hOdEc/Toc4DUUtXyFc
M3WdQAEPHHyoxCAZn8M0A2ygUNRXswpDMsK/xNMAEyVzA9cOir9iGJCp1RbJ1kqgwnWsY39lh3Hr
AellPnWZ9+Abs6jASzSzicybUKA/vJeowydrarR1lGmX8c4aqzPHu1s5sR+ExH+iaE+VhONW/dYa
/MYA8g7I27JJWsu4l93bE7OD/OeImJViM8iBAjcuNFiZ68eH7oXYULPuLRFh/5eZ5RjC8pS9K265
df+f9sMi/utla3WxdC3oe83sfmPwabG2DKGO2G7DvMK+NCPYxIc+SNcbsPqXFovO9rKONKDvi6Vz
uXp8MbFyJ+1Rkwty9Zoq93OYfFDflepmGV/DaBtGspwiksAPWDgo4N25T2AbotiECOc9sklGcwNp
+rVSv0eUCgfheuvXdwtjxiOOBZ8SfiI4MGusG381ws7TfEmq3ZoLublAmgAOYryFXWOyPyBIoLKo
YL4ZjGgSJVDCpU2dDH8zQdIPaecWpS3r95afLyy/RKWOwcHzyTZ3f4cacESq49yGPm7fm8k1HBnm
YBrCoxpbsfx1fBXRTRhIG4zoBaHW0wGyRH2WEGZAIet6JvepTpsiFQ6tveWkffPrRhzGePx9XPUV
1FaJ6tdAMmj5AhuZSGh7wvU3hjgMhIEwvTXSWB227gfCTibW7zInJw3YhLWyFLo+wNFZq7NURoHw
STc178/FvgBAkcLyho+CAG8ZT0ucfwMzKEJlyQdFCKa3dHFbHj5QxOdnN+sLRHkXv16fcthG16wd
vQzOZPsYtRMepQxrmdsaTZByUj6EAxLwEpmvv4pdTvFG3ctmt5Oa9obmw+CMZ1Xid+Y5ztXRAosn
sjUjYadbO1++yWqtgSj/Nw+VCQp/60Wq7mAUBIQDrkyrtyE2KLDQPWhc5cMMQfDNf0ZRxttnp2VU
oVWrphcmOUrXMVXAENuPROy3uthnAQnNS2kYMKzHTScXR34SYI/3ozD05DtNypa2QB7cTosfZz/y
PZabBCmMYi3oKu/DtVBkbRqVw74I2968WaDUWQxoPxqoTwgX06Zmfog71fb0vNC4iiNt23GGTkgz
stXwGwpTEvRFoQLF3Vop4SHyofAoOH4Prk5wEONzz2azeAHJjFsnGCcApNqQOqrop1+9Bs6omA0r
K1JMl1f+wc+phTE6l1prMeHkyahs5yB70PJDrxGP7xY2RNvwg4i489eVsGK40kgYtWGRnLbWNPVi
fjKZzJIZZkYbAcCOSIpTS+fbrRlAsExhvLq5ZUwK9C2t5vScQ4oTAt97va7p6gU+1Lrxe3IZER6W
X9KONIjgvBkuNh0Iw6kJYYxRx5xM+LnCw6B4uRTpVHZDKFBqKE7jFiXZgT07tzVOH3qYX5dmFxsy
XaMzHqx1F7tOm78K1ZBRrSSDBcbHSVHED4vZqxMs8RjbzhomFuBV32himvrsbOR7XKd0QQfbP0Ff
bdl0mzO0590LqHZ4/+hgBk+XwFglaqnO87K0bCKdgXBjTiVkY/VCSD9+0YNvIcn/oHnOWEBbxoex
44JdYXXpR03LCk5NP4JAQPwFGMGJarHINEtVUaBYgpmwnjufZLsQW79X+u6EOlGo6ozYxyFM3amW
uMkcVgp4AdArT/ByI3vufQG6O6AtNMH6jxhZFW8IyTJDIcTBS8p6JbPYaZlkajSvjrjBFOyzBQYX
a0DjP1xrD4ozol1PpES4K8qO8hGP4Fgo7I5zZ+cPOuGaLPXliyE+WEAmrSjJyGmN475Y49JHipy2
zcx/4Yo5nfvlYTJHrGBOehrznH3oKgaIINgU44kq1wHAh9Tj1KDBeP/kkminCHH7JEpPQ3i0V+aI
y0OvOikQhPqSvyGKKlfW07VFObv5Y9LpBxefTtDSELlOML2ahMZb+x5u08mIwkmTaWpTNVWqQlik
Xf17r9amw9NkZ5cQtwMpF2KBCSPQcEIZbbXNVo9SmfkwpgtVDkK47IIyPcf79xZeei9pAAsDfMVM
BRW1kE9vaC38mJ0YYzqhhUV/q4hG4pgWSZ+/dTWR76D3f+8vVGqpmu+EKq3JvObFUooTDVK73quQ
qBlpfnx+0DmLHCq1Y1uZ/83/mywukTkvqDvmsxBOge91Mu7l1JyLzcp4uXN/TfDWKdhzJaQkqcm0
ausINx6BUsOb+YO8xk1f5jnZoB5BKJyFpcqodIzVrti8frA5TwNxFR+GRMxUaax071tGRtGuzE47
lBM3STLWlxhOgVmx4uk75+hPBwV3ydNoOjvw4CdqBsqJzuiONhU+OwfHFO/y9rqlq/JoM+QhiuZl
EvFgWRtBBeqkj7zc4WCYmVokPOG5C0x9Ml+upp+pw7HijlrUGcmowiqUFXCHRabppvkunQ9uNQC2
vI6C1SFFIkDz6Y9ikdah5FFbkeIwnaW0i7Pf0ZKcANIqlF6tq8O5GDnE7RkhSooX6gbQ2bzIGcBy
45MAN8UxlEoBSs4zbrYz3pfBGhcQeoijYw76YH/sw0cuQ+oV9lxuZxOuS71+4bEGFY4Nvx9XKDr7
KCX8GqDMe7rh2usb/fRf/9Wl1AnnqauYMAU7b6UFXLcqGDdov844ptHpAmKvkCAvQob/3/moLDYY
FjgIKzX0jowXUCbrajrL+rwk0MsMKTHJ3J6kUeMWMLuVzQ6HdhN/s2vL+siSkurJvlPTUz66R1Jp
onytGGBgHTYurRz51lnZYwj5OBVqk8jUbpd2cF3YV3+vQf6u68O2Ny68NXBLbGjAhMPOrJtVag9o
eXqa7LYEoKlEgzmn25uzNDFQ9WFiKNmvmVit6DtyDJriTvOhqip3LQ2uCdofwiHgXfe041U4Zv2/
hK0XGiDEd5+xjbyAtaZaoWV5yTOKyI5GQlz+iuu2sW6i5K3Z9aChOCWAQICgPc5tTEhfxyHpD1Un
iy7Pjo2zfiCB+HFHk8ICT5URXHbD4If2Sj90U+8a/u51YEwSi20hIxL89FmHiPgpmEzr11zowyHZ
Snw/BMOKtkk32xiPEfX0D8fIuzRcIuolPqRFHUT1DWuCTd7s+PuR31Jmha2D1jKG33T1o1U77Wmi
kdPKUnF3aAjr7AVdXa++j5E25nJehjWu/cyfDbQV3wPVFo74glXnW+YEnr6+eImBzeqrJD+JiG38
0RjiFNxUPqReiBmSiOvbdWcHhvC9b3fXhvWA44w9keZpsmK0wzPT9phNwItxacy1nQnqXqQlWXw+
4pZHGc2NypoliMoG3kC7PEOG4kJ/sXsTgw6zajs62NntjrLd9Ksu2x9xerJgy/QBFil1JTlOWuKn
ZHeNUmN4YqzOWoqGZ/xBKwCH0t2Zvg0XNuf86BleCcdgPsxsnmSzAfBLPBxHKtkO/hHCX9h8P91H
925WY905WUWjYDrln7UVADo4P1zfijliCBuRQPreUB2QrfmCViwPSWCW99yyrursJIbQbb0jq204
FK5JYtTgU3TxQHlwJb9E+UsbIKat9LZRaQIsoXGZmrcmkNOq3r4qP3NinZogeHEL/AkKLxpDVMw8
mwhKkUPLeKJopvu5VLDEZo00At2S1EowAsdX2Yt767LPe8bdpxydrdhBaWTUMb/I34siLRNLI0r2
hDc3vpVFhkz8nLY5AjPoNpE17jCYOIJJwMUHctsCuLF6ZPTAkPrDF9N+1E18harzst920hBBcQdL
CjxrK8GVRQz8gsUk6HhWJUxKWelSBiDr+yHvlPxN2HqDouUT7qKzadjTn8b7nOVZfQGT8G22/wPz
8QtHcBbYUs0ae96IcNUUQhKAy7fbm+hBTLPnjOK5AQ2a/tm0Toh9QQNV+Q+trKKHYuGx19qeJARg
ozX4X+WcDhUU9fPiGUKqzSvUFYlL9x1U1xw1BM6ppTa14c/2kLi1xHkBoWtNfWUsPh2Wx60s4Q7/
njVXtazS2cXoxc7Ck8JKV1k7oiL5YGWyj8c8lcfkeMVYVNr/E4AdR6fYxZae2KvPOcbbcRQ+29cO
+Un1sjqxWxx83mIzHZNl7XNDVPA6zVqCbcKkN0PmyBGlRzGUlXHiftlYB8ghMqYToiI72QRu1dXK
Bnwrj7/hHdf5Nxv7/xsc+DHDyr0TJ2PSWMzuK/j8h3wJDj1PkwVO0lJGB0lghdNNpn4sZn6Fcrb9
7g7NbIdCEKs+OeLDDMQ8ioHVlYaLN3j2821Xb8tL8lOIncyGbng6CRiUNyV22DrwoozziNk6fWyK
IAXGYaxPnMgdNBbOXkpGsZRX6aCwStBDJnGDesn7sTrrGHXohPnW2Op3QEp8GfwiWs16kzC23baB
u5Jhm3f1CUNQgWrF+k+6hQdHhVaPxtnGQQoT8WpQumsDT0jy2SZ/FEOH0NZJwqshh/DoVYTeygvW
NByWAqvUiDy3/i3petNuTcY+d0WN7/hfp1yanSoZe1YNNmt/sGw9un5ocBvHlLjf53aWL/73ZcFt
c73AtcbbcAtJWfW44BoGbbS1WUNGq311uYW0YYSn199A/KMIH2KD0MrUIfbPpNcRK3o24W+Y0nr2
u+xXZQd27SeOL4fNF5mkuSS005ih82O4fXocyQ0XKK7CT1FBnJgReExILM/oKqm9i9Op7McjF7kV
7PYgXtorrh48IYn8oSBYnNnOyZgP3dkG8zqwbM6gbkfuYgOpgB1aSQpsMvGyYE4QYsFS20LfVDbz
f+L+zX5yhSPA2FtGLlfqG6ImP+zBpHSd8xM7EARnSLZr1p4MQWuFjJn++fpD0IzbPYDWwItY+oMn
BxZ5R2zv9uOApxZNqWeNZA1LzYaLSsipLS/FSm9/Ol0T2veSULXRqt/UphAXCBc/U9DxVrcwBOfe
luVQ1PLHgUtk0SgScwhjvi10+GfTz74tSmtEKPwfdIBUeo/nvjy15a8VaBiMm9NhS2BLCKg4zlVx
zK5kPPTPUYYhtl5Qr1v2PWaNRUB0QlH1nF1O4LKzvitD4ObeMy9E2Of5qd/EpgItwv3yIZxJcKOu
BABRUIvI/21Lp2+Bjw/YDi7m1gpJpd9luzZmL19lyBb/P444XbhdZbYG1mfHYOwGKDp3ljXSGrO5
kBXbum1H4O+XV2FPPsmSWtDFS5S7+i1mH1NmvPa9SoFivPZWzHxV29Roc05xKkxMFLVErd0RHx/E
iSHV+3JfU4/MZT9qf/jTSOqoxTt6XAluTckMfS0pskdlDGU6nEco5rza1McBgl8bbvhhLkZVamL+
TvaOyCPyc8cBkDRW+qYV23c3jFJBIW4bsK3J82kqSm7PCQpOQsxJ6KXyklnD5u9ZOqPAwjKa0JeX
SD8oMqspt1Xk4AL5KiJf0AR4uaq+oRn3mBOKEA33Bw0EDYB6VbrRxgP/Eja1dF0xzV88GAJSEaHC
L2gdsdfSfARL/FRr8eRSsvKArFysi1jxbk37FCqsj2uoYk3xDcnMGgongXAgkanK8HrJ/rt4AE6p
RWQvPMO8Kez2soSq4JeWfUncSTGVVAYdqqZuqCS2252gq8o7YLGJHNwwGQmbxXWliSOT9Ba21XN1
PupIR9Op4KpOQV9vYhEDu7fOeFmE0hAMehouZYMKNSqEJeZSAFWtxFDI10H5jSklJnuImV55nCLh
he0iHe5Nv2YgTIqbPpLcXWS6w1o4JVtdrHAJwoxIbIv8nVN7G78AkskarK1ntwzcRGNL1/ba2wfL
LmWjo0xNw3+ixYEQW7QpIn+qtwFCtBa9og8gjBU6WnBjdl968gH1XzX9eYxLApWisP29RkA48SwS
IvE2J9FEQGnZxE1ce3oR4CDxxfalxxcPgo1YpvJpnYOvN59hP4GC6hC7VZA24e757cAgxOxnoLS1
QoftZT1yZ1VKBj6n3yZoaTRZqbuv7HlG9gaQxWltcZCZxGoJw2OyMIGTaSk7906wOyIo5u3uCcR8
tPdE0oeie8mVRf3aHX0uZpQZjg53PDBeFn3wisT+S+j3glPqrWTjn4mhKXjehLxKX4McbNPYt/OP
7JhtQCG8d2kxjyruePqw4dp4Xkrwciu10nLSIYnLRFCg8uh1RtPj6sUN+1TtfXQUuuX/MgPWMw0U
Zzz5+Q6LBz1Dld66wPCtRqQBQUJRWkawMIB08bxneynGjI4NHIJSAjMLxslFf4gAncKsm1pGrS7g
2sbxXDZRkpIkIN/8HTk4tToXHqhsjVUiSwHo1T958KmV/8WdyyYVtJZr4pMVEMkBKaSQbJeLx3r6
OVe+2sIMwDjNU/4XE/OBVyjDHnVjA50gCa44DiDGQySop7xN3ypBz+e2XPmtR/4xf/aKVK4qELqE
//27t1+Nf4V4NiOxHa4N+B+axnzBUSFVkMjoWko8CZIsZDOu/Z+psY/6bqOd+g53Uhe+O4ecVQpo
ltFkYxj6RX7MCf5mytJuI9p/7kdoYJDzCXM0+G2tt5/Q0zj2U4NAfTI2gQkn4Lv1vXAAZTwmkHeN
Idp9QlG6IPZVokZA33L26/g+l2jhou/jdImVlt08bgYGLwlbaokJ2+8ZDdJHUwCQSm+go5axSowr
20s5g9drKz9SVQteazBfboVcXmviOoyuPPpN6bWK6RblPva5OQ/bKnsrgzc+zjVA9Ym5jo6qsWyC
PluaezAwqLCxLoWO2sxN4AQUtakskpYIHaO2CjFLCLJtyyeiA4W+U1AUbsVIIHoulA4/z0hiqd74
iFqAZ2BNsfW1ZCQYywEn3CQhC8WOidUjAN4sz9lXLUCBjWiIcX2zYj4/8WEMgG4cKUBjT6yq4gAd
owMIpKMW46YqZRZAx53utjydCCj9RGtfGhoiblQ3dDh7TmTSiLubX4zjxeumZTstB4OcGYkx2GH+
g7WidTcE14ihr/hp2fxVFu9HnY0nz5QRqxZ64xFQO+OdelGgi+BpkTHqJQEGgCo/bcUJVuMwOhAG
jCZ5rr/lkb12kxpno6XbRqnk95/kc16V8h7M8zMNXkfm5dXel39zRGUd5WhXu4BMPI4RcI1/Q8j3
XBA5Uw63JqOkFCkiEoyQUyc7rkjVQoV7pg48Oo7EqDPtMW/Q7Ymk6VzT9Q9fZxfs6minum61sGwb
poXhfnCEFG38UVKwTENUjzlxWI7TaGy2dyIkJP5lQZNbwCW+W09e10ZVq77jRTm/YgSNch6cppBh
+iF+vFmL2Z8XkCQXuao6jSlJ40KYHl9qtQfFRJGB+NKSs3ZnVsjBICTWX+5biZrSYq3vN0OlGn4a
rzAtdPpsfbDiW9pCAsOqOR5bgr27B2XwEawAF/5nF2Ygw0X6OJpFHgdLF8bNRPRq/2Lqj4LfgSdL
6qXMm5eBoDhmoYwWgaKUZ1NXbhQmRuZ/7axi6f5CC+0Kxk12FyeImdSOov9aaL/AgfDlhA0rJxhO
RSIEZiqjSyabRlweSIkccuzHvPde1gh2gYu9YjbJJkxVFu/fGN2FXd92Fc02BrOH3KZwQHoAsXf5
yB42SaYD6rzUVjX4fMyQ2c6M/e+ETl33vY34S9ncjTQj16UQ+7F2UsKwLutC/Redx1t9mcLChTVi
z3Mmc+klyjUiKwwqH9NZiHKLBr3kAGg4+j+Gs5s2qGT8sw/sdvwW+EwoTQdZVXom4xCSOasKKXwX
bSsekFh9hbZSK6h0ZPxnNGZe6rNGIoeC3fXeSSIe4owVH4PDkpGqA/Ee0HlL1NvO5eQMTzSfN6s2
2POWYNNEnCIWBW0mL7Z7t3PriRCww+OK0uXDq9ElLYMJtvCYYr0huO0h2cFgmBDoqV443W0HNu0U
/h97YUZtz7WVMN77RNe3968lr2vnJ+9uVc3IrYc1YrVNUQfBnLe1G357YRDS7eHXalVZJfmTR3NJ
ldPl1LNkD1X0+EgjiU4RopdYs37rxPJi30+lR6BLY9KRMnbQnMR8FkB//58spm2hp6PiqGOQzAC3
jXCvK5cdv5Q2bICmEatR4/VeliUVkpvFYQq7riG4ZxVkOTYXxloED+I3l2QfV+IfoiPboqMU19KO
2d3h5lsYv0e68xvjkE3ktewKstQnA+LGeepWMKS7S7RKPQ+wRSkRkFtJi/mlDvCzCmRq2UwQMKD8
4jch5RcvfoaqLoVUnB59+SjxOsVFC/fUkGtygc3usLAE5jmCQ4wqwaQqUIhO0yuwHSut8XSmygh0
+HS1cEU7HGggme1QfKWqk1QgCoZM1eWMTAWJX69VuZSDJvW/PHSHYDxLT/Ikc0HciBSr0eqgJFVa
ic/4Zx1p1f1X6JAKfE3+U/pLUWZcn9pGG2CVlOqj0/TxDhgaUvppsHYK0/KIP/lKCGrQmAe84HU2
Z6O0NeRv+QsBH8kNH8Jl8LDdcqdtGobBKVrIYi19WeWCKp6bDY4qaLHg2aP0iJAovoz8YwBD3vZa
I4OVgaQzOPF6TDgjPFGgqZ9+VGuTqzERnTWZ7qj2TbyPnFKZP/FkD+adKU9ThpciTuHn/81lk7dd
AVZ6WMV08Fe0deHi+Yfp7S9ZZesEz9JxbLrVOSko1/guC2TIkpOkobw4Y2ErmhUtWocJ95a5cDF8
bfuRLJXty94THWYx1oUDjq4MLXzM5Do1wY69y1U0QxPrFEMAPQSoBg7HFL6or0rgkG/JXgxYXeuc
NkV7Pc4sn439qu/4fT/hAhJutO5amtzDNOIujzhANF8ChyXYwuJuDIKAuUhw0sZtq1BhriPTm6Dc
+xgInw/xgyPPFe4m6qLfkpcRlieoERBpYFYEjjHEvqy71cYRXX9bH4ibnk376PLHjlu2Z6HeLf6i
aJb25Qs73eRjOY8V8GnvkvxIw8IabsGmVYyygGaMfVnngy0cn/lXgsieMS1hpp8kNuSIsMdGevAi
iMGTXwtljJZwKTcjaGLX2waXWRdAF7E3RxjC+fvIXQ62gjpv9ZTypJEb6VCwYq2jiQ8kTo6LtOMs
ic2czo1/aiAmTqhYAZKNglqUf7NS4b7wYNM3z/SV7IO6ad8xWYDdd5MEceqG9DlqnLaJAGbewpwF
ETtCdWAy25k7Ncsp9rYfWEpd3LFtkua/gnrOzqfXJGHTzMZD0tVmucz7aek1a8BIR4V2jh79MwNH
N1i5myCk1g27rYck0tm0HJqGpquz8w8SLopByWLgLHfQfKx0uHro29o9VZ58OXZLrgr/rmacsfdF
4R2b/nRhcFkzP9jMOAI4ylJN41JCBKhWk3hVRLJ/qZidCkPH9xTWdPEaMOV3QQsl1IKuxLFveZ7u
BlA+FLkpWPqTJZuAJ10dunSTlVk9/EfqcfDFsTm/7scPyhYX8zQJ4VwlUW20d/ZrC5t+jB1W0AFQ
SqBm/D9JdKcuRYhVW5CfUGxS0AW1y23QpLMHddAYT9LX4WKf6kjEc4p9lTJZiuVBeE1j/GU5ehnr
fjbv5QZ6QxRL2r4+IPWMRzzuCPyWx9HIyPGatzkRyQOKgJROyURSb3kAckM5chPSdhXzUql7wwDw
/hNeAExiRN30Ch+K1AVDq6mC79JkQPPAm0hZJQdNishBhefuToVMZCxyYckE45/icy3njgTZa8mw
NT8V1LJWvis+XV4NtFl1yIsYV2YZBrQdtA5HNfyFOFzBgO9AJS4A1hK+DnFVbggc1UrcxnXOfaDs
lq1ZFC0MVhDsGgHLP47gL+KGHPpirZ6Cd6My1SrYx3IWHoaxHKuHRvyJj9schiZ8o3hKY+w8zSxf
b+ehmqRg4JSIyHIC1KAqkVi3wH1i77rl3h21G13kjaib9yVLdY8q8PJIYWg+LC6oc9OfhXSdb5Tw
shlQhgqvwf27nw/0UxygE1LQE7M2+c5pchGmiHQKLhpYyCOTA6JhbY3fukPwN6QxaDDGo7y81QV5
lF2SrATiy696ks9AG1Zdss6M/1C1SIuRW501Aof+9wMh9qpIdpafJYDfGm0BrmKzB9zCMzlpxQRS
CBLRRlOLqMHsxs/YwIwFDZLLA45SA93RJHv+SEiSsXLmMXTEUW1OOxJMSNDm5S7E4CLmiBp77VKR
zqFD6fPzWehcURoIK8x/VDbf/5grR0XmvTIjfiwQ9gV723RVsELzWwlgxITCoN5h6MovLgvuu6DE
eLNs74ZHT/TKSEBwsT+UaH0vu9G5qZ3ScoZkK35NFjmE4VXNeZjLpHo8RNQBbKT4gOMgY0+ECmDe
gqBcXYk4Y73AP33/jWmjt7AYfcNfJgKSn9MVf1YamcZec3xNNAC1RBbIpQyBxlbVmkVWCCc+N646
eMKItF34fmVeQ7IR5TKalGilO7iYJHufVg3EQsGBAmOnLNE3qAtTBOVtCtrnrsLe1fZ4YXMoV+m1
1lWCLvDcqvOFWlF4bYR5RdZ9JxyzRzEUGmhrPcd4TbboJX1sPc4925duymBHXPfUALaYqhrQm5z1
VzETvmCw3v/sP5/YmDtU8QYNoguXJC9hO4tZo2wKiaP9m0c9X7V1hPh9oKMyWlzA+TCcin6Wjak9
5YGNL9aTTleM/Uln0UFpnw/ZVqyYxCrXs3DqnElzfL5kV462rSx7733pLummPzy9J64xgCOzC4EN
QIyoIE0AUBCChfsUhoTA/lQl1KmjNdvTa0ZEFIMf3yk1KB+6Nxs2b6No3YFrgffDIAQs20H8wH5G
OwJ/Io81m/nOVeDPi/WGIZ/gQ2/0fWL3wW/4+inojinVSkUDI4MzVskEWTQdcOS48Lv7G7VAEXYV
CBVlstDJjcB0xFEg208BMJkGfamnLojyMV25bBQJohazIVth16NXYvh7FDVtaL23ap7Y/rR2WkMM
I2rZoYXUrc7ozH5yhdlF60sLXrJxFPAT3AQ8MW0dF8VR1oyD2Y/NxHN6sA+41Ngyy1Di1EVpC14y
H/sHT+6MyQ+ScjOtuQr9c7wfN9Mw7PqtQK2C/IyiPVLLa0O7wF8QGuRIGAkPjHcMau8Ey3TxvcP0
mCfjHd2htk/PT6ezVQJbmeoJU3J8d78O7b4H9IvabNeMv4w6Nr0CkDrQ7hjazuT6Llnzo81INspV
u3JezjTE2D+MH8GIMaNhuHay3FcLCOGhoHcyq4qvBVy/hnkvip/lS3O3dhisMSmdLPlD+ifGAdxM
trdnndDAwO9mHSsOgh7p+Foh5Z0prQHfeXrGQAmifR6L/T1Rlz45K1OGQn1UxwWLAqYWHStzcq60
yZTBRu+9FH408cuIr0zyr19y4CBLTZY6lfV396uoU03ZHtegt6V7fBx0Ft1/sALZGa1VI88yqkZz
jHMQ7dAi2CGQRAQ8pMRPXNkS0Dw0MRhC+yWUtYSoK0FVQEMIQ1vY/WxCF+rFBo64yqg8RwlTtGRn
1uCFa+LXnN0+0zoELtrxrUhbvvqHYhGmDHT5Nl0LH2vWhgLDCfgvSRFkTCH2dnE9LRadSnKkr0DC
RpB1pdyx4HQnuIVApMGDf3QFHKFjy6U4T0KAC5y7hdKWmRU0ksG+df43PUsjbT7Gp9WcWlJOWde0
ky0pXunvAKwHjFPGaNO0TxslawkCT9a+8JbLCNF82cW5ch5X6WDTjW0Ut4jA1eV6AzOUhOxLZMuv
kY/57r+ss35S1ARNyqJfsMshgyTWK2pNJOgKJCwsOSqbFx6Ro0YF39H1DrebdXLR59iiC2RUeQS4
RFnRlceHq1OYPXPQHr13ovbukFSnx9D+Bp6bSqM9a8YbtXusIx4Hqq3AlBpuAGZnWzK/PgmRGzGF
OJnbJ1k1hmZ0BJOzisD5IvVv2ps1BGOZWOEmL4pTFOyeij6Xh16r6r3gKuBhDYZHwlE+ioegYsK2
xjPY+wdl7Mfra9btnpyjfILnA/yw0Y+XaAsQ6kFt/lp29FlRlmhw9Zna3mEiIf4z5tmdBAjQOlXy
NZWNEwij7ZDVmFqoFXWiB1tB9137pHnD1DGsXGxV0RtSKRqgtyVwjr/ygxA+ujIM0cLE3R5hRL+u
n8pJlvvMDPk7RhEwGYBMmg0hc2udpOOqcRbVNybENfkrKUDMEBsKIqfulxNa5C/X4MAe3HB5ud78
aHh7RcE4OmESn7nKoO3ZcdI+9FfmYxJpt0fujegIorYjXCxhqUPWo0gNESbc2t/iiKO4j45YGzrt
mRHXt5HiRO8Srnza1v2rLzbcJbC66ncR40vtAgQol6lw+swh26qi+dEdSmjV/dt3fEzyedRe0omW
dkIabgT9xlavzFZvyi7Pxnohh6KJ+tIXVcvl3qknB6wSQ1KWQdlDa0jP5iRH2hDhucbGrsuaEYiN
5H0Ak2o9eI9B2vMJQg68+zMzgIVDbcwo6I4M7YxYcKdwhTPLWmMGyu7f+QXs5mXF1bk6f/DrZcrX
Hzr7GNHMhEDHo9aDcwIQR/1RttdevIWDM6eHJIoPMPSwXxlOXD4JXbPydyPjol5+aLYoAvnHca+b
wnsxMK6FWZJ3CVD/IkS1HXLCskbI+dwl61U1Nfrq9nWttM1qs6RzT9daIcL3hglByNWLGkVQPC5D
ummectSxYENBYneyMyi7cxTs4xBrhlHd+js2YD/SHEpmtQkhkoOMbumhgjiw7reQOwmHaI9CyifP
WRSrZmxB/lIm4Im5TbsNvk65CtGAU8uR5nlJOwbhgpe/jSTDoMO0lvwgXkmXs1ETrH1OcbvljXg3
ZgItg9kns9FKezslfYuj8IaGpHcwV458GkpFuJiFn/mcyk/xKWUBcA3L+U0QxI/kUgxq1hcpm+qw
P2i8DbBCYKqkgAVbmcUKuv4PPt+zDEvS47SfGdngNkgvnAq2L/YnPL8/Ym7LRBIXSotwvBSM+CUC
gSwJGtlmLUHRHWS5xvukSKwg+//5nzaK53Y5tfLDBHtVDisEz0uCa6cpR/V1W9Bw0ncR3nTYZaE6
EJa61kCjp2zWFdo3OF+hv6QNuKqY/Zs4aqAI+1x5UHtKvCxX0+ZhB8HsdRTcE1PnbU+1K3EpheZ1
tNbSKFB1gZgrPsOb2TUwaTLeohbABIzuAhVT3W/uXlFH/Fz0SXZnevx/uUMJXxaxrYDwnJduA3Rm
obNh1TRooQLoYnH1QGYiUwNuoDU+WCCBd4a6E+AaV8WXZfWviPwxErgNaj2jaPBGySSsLvByWrGf
cs+LtPsjdSWjLb4HPQf4k89+NQ/DVanbpRNE/z+TNoTb41jAZZRbF4miWqsT2GAMx6HvRbubf1Q7
IgY72U+RnCiwmMolEl8CakYjd/Ic2BFut8e80Wd0pg7uMZBJQ2SZog79kBMiJE9oZGbbCIZsMlmv
kX+VYNbvAyP4p5IQBdhUC/xr+eUZzdKpESYP7PRww62R5FMlWQi5H5eDQZQT+lETNtXVeWoJfUXY
vCsjuXT3/pR9rNFJHa/V9eueWOcM8kfq7ahdqm+ri7OFnhC/ooUrUGDLjnpdaBMEN89AaUv8JfzV
AAAlZIKu1YXHo6Nry/9cae3ln+WWHAdSTmYRQIWwvZnntscnkM5oPa0XToOO8V1D5Jn+yCNky/mH
+9N1yFwus/nVABLS8lr/ykBoTan9DIRyhLnTSgXGhpvfj1gp50fui554QblBDKOuYcYi0yGiPDfQ
uQHwilK/TTYN1rRpuwkA6ZyCqGfZsW6N+QL91N8sbhWC9LhJ25XInWhgdfSqSn4scyxVwGG4UE0Z
RMAejvGpQgBAaawqBtKg5AgvrO+3tX4HkFkVGtPV+jZcRgxzecoXXE5TAxBp//mnddbKatHO15+6
C0xRS7YT+RG7wT7GMBobluiOAMJDVH8x538YPQCeE7pB0FGYtSaehXe7ILZTG/Sl5YyeX8Rt8oB0
EfB2QUHJ56YJ/4/b58mLxgdHBAE3XpIHygEBtU5ROlQsaihghegiqWH7f8CM2RN2yiJBx6m41r+R
Ghwy3FWn9C4oULZ8ELDSrfzdog2UqbkJsUuAr9JP5aH320BssymUzHoYecIexJDjb7rAshxNSg0A
ggYhRHctMQN1t4+EbPMIIWpuo9XOD2mOw4Ql2IrqbKYsq28+x1gvpxFsQh8H6wmmEaOMO1Po/Pde
cweRi2owa/EpTO76HS+gITCWudnIds+i5Lyzq97brNtV4JQCGM+YHc13M/GLgyhA/kSKZMwh8AhO
VeDX6vUTuw8As1LlQp5w65hQ9E2RIgef3tODaL7ey/nyMIp+Wtx2XJVEXYF5wVZNYosGbix8yffx
+561Vl+7M1Lv4XGJjEUQcfqBRFX7MQiTcTbAYrUFglaeb7mrh/AKN6XkZt/ZOE0DazQIGIf9roNX
fepvn24vbqxI3iSd+CJVkPg4BJJQNNxTPZoCd7Zhb2ap8mLlabuYmtMtIQJk3D5I61JMls66PwOa
C7OqkzHiRaB/zkL8h9BPWNnAYbrpzg1qOv8XL1snjatxyRZoP/j6fw+cJ79Dy98aW4JrWOjLYI0R
oaUWwsGhOI3u9wI1hnX3QQ+H2Q6cR3rcQioTJz4EpvllgeiuLd9T500k/i3w3tazgYP0HXu+z+rR
OMPROWKsGthVvjIijv1087A+N+kvPW+4ij4ZSZvUw6VfHuLgyLbdBYugWj4SYS+FdxQsFx0+UIQh
t/5ulTRhW9oalwdM5D7C6AWmO14lnWcFrdeZDWuFj2MyzbRYr+XPB5pubQRKC7spcIE86J37AV9f
sCA8TE5O24zLr50J6n6VJuP+dyymIFT6rnm845Q2IX684ivXU8SF08fXVKIzPoieS9bCZZdCFu8t
W4JucC+tQOdIRKjphkEzbrkX07UCzLZEiMVuaj8QbtR1NCQ+XRk3e25Hdls1dMAOVgWKF3Rygjv0
2D4YgqTPtdqqgQ+jydQ4RVnaRCjIJQ6DW+oeHuAbOB9uej5VaVy6b+c1pse/6IIg2IcNWdIJ0a5d
9m3hYwScW1vvKCCYcmSxDaGHKrqfhQio5/NZrjFe+nO7be1LFOK92zVXXTBas5xTFFbZIFVnaW6/
s93ZZ58R/DgL1PPdu8jXhZmSGEks0lMj+e/QGK62Tp+TOYnTXcX3tRNrI41LNpW1DbVDcNgn/s9q
N6ggVi3kBD5c5mBp8UGIkw5HdF7R3G+H7U0DZy0WaUSvFX0PQTjvqW21tG+uZBz/pYnRs6F78h5h
gzZVRnOluy9XHZ6hPc2YrH8NBax0OmQqqC4Rnx6gMt1oxfTtuyXlECAIV8fyDdldBhyUVzrzWqQ7
lDzU5YczPkaxYdADXPiIwvVwzoNms9EOlVYgxcpZROjlowou3hBiBXg0cs56yN9329KBE8KFzhe4
AU29l3gHbguJlkuwVqnYtlaSgAS+OatTsnwTSoyZeTqz8Sf/svZuCqrwS+GcyUTdMtvFgmQ44DDZ
N2oGeTbh2UzdwFD1qyJKVyFNh7fa9KX+eWUw14GN7FKsk8T6dflFAOWmKcBCWtDnj9l+6lyI3/X2
dRjmoWuVpwQxdKBh3hsSKjOYtWOItjZKx1ln5XTicNfD9jyf6a4jT6pqnh/2mminqJtGLa5Fzajr
zpOoeQnnhp1DoXpP88ARKEVKSIYxjVuJUmEltVjPO8wXsBdyYVACC/4in5+oPRfPNzQU7GRLMNn1
F6CgNV1QDZo97tMWoNhICKXo5Nlr/ognIMKa2NXyOuRwhD4LgH55P5wKBDK07nz1KF55x+yn1Vzo
Nm3jobaiI4W4mwu5sqP5478rhZJ+4I6VQFTMcivRIweAlU09tVnt8uPX7Q6hv7JoMNu/b8kZmuea
dagmvk7WPb7W9S8GB8x8Fft+HIHubtbmjn/QB+aRURl6Ad3VEwyu7+yVDldcW3v6ZaRx229PVQLv
2rf7/TIXda5CuXXsk6qvbMX35W/OZhtRKj1LBSTl4ZWJMZdts2Ji/89NLbqNl1NqIgxFyVCIRWzK
OWe+0a0HH+wAQKOa2IxT6kcVFMbhYWBl4WamEAg6mIs4HzTfSfP4lEfTQ71mwGsajKwz9wbcCcuw
tK/IJnBq2hUSU/iAeu+TaVVRbvFBfOi9YOqaGcsZjbZuhe09S2+K7wDi/orm8PFWnu+Zeu/kTdBd
cfmsDn6plOtcnGmH8ea71FcK9OPtM53ISY+4L8bwnlulN3bVd5j4qMaRoYWahmcmv0qScjobPpqB
aEEThkc8fknrAe13Fj2g0ag1EQuOnYw9E9G2mOusa0ordKa1jdVr9pM2jLofaPw1gLZ5XoeGcmKm
Nr80kwFMzLUdJnyfrVs2gH6dVBt0iYmLRx9xUAB/h2gPLoUnV9cKQb6OI5KfNP++qsyHyo3uJdhy
Lt66RB14tF4vnzCFtXXnq/2QuP+SikS0tWcNCMaChaIzRamD5QKkMm0UEjwDJA4yACx+GK4L9Sbq
oGkaWWSOg3wgNDhUXj0UtaQIXTvxjhveW4LT+HzbBF0IhPsff50xj8jUD0Wo0DX5VxNOnIP9lBQL
BEAvdvERZTxaWTdD5keHgtQ2y5NXq2OhZcb0v6I11iRhu+dk2/0fnNC7uJCMpL6R41vNIaRFm4ao
fzL0ZPG28XCFoQ7PAT0DxaK3AvC+BMvG7n+irdCwrJp9z5P0XgnFzwGgl9XbmcEBC39Yz612WMVd
rQj3ya+RDCSnVfA+UpZJ0C/PUJMVDcXjrDWt4MSF2Pso8aAKo8iCDtshDCHcwI6fRNDCcUT4vxPd
168FCU3sRZv/zba62gqy+V8PVLStsXuCtH87JQYB4TQB85cuuAqqNpM59DKaaJi83AUiXbNTes3S
OgAy901tnINfqtNowh7uYR64KYJi1o4k/XhFLUqrRpcFEc2ObJDOeHnbo61bAFYb79AoNh0zln25
z8gFOP+o2EO2MXEW6dALhqxRkYg24BQfGXIVSH6eHyFPDTBoU0qR1N1iv+zNaedGavNYsZ9n4Ea7
LpVWqa8x1YEbAkgMqYc0C5qF/y5QOI/KugVNhp/9dxCQJv8VC5jGQ/vk2AEBYNroJFkeE+8i1VeT
7WQyLKl1IzEn2r8PVxKRyHpF0m1mNlUulY509cXOf0cIlBMve5LsVAz6Fw0pA55R1MBir1AlXF2a
wxvragoaAmB3xSoUf/ts10RdO1iSSo8wiK2SVDoNgnP3mwk02XFsvy0Xz/THzQXSLiKxKVTsDE2T
7Xa9cP5QUkD/2st2q9Bu3NfT+LmpEsgrk+r778zwCNGX3XJgb7fWNekPyJ3U5lxDMbPNBJXQKxyb
IAKVl+JNemXsQIw2w10PZ7oPYhLpu0kGFDn21RJF/xlOfFvNYFqmBK0c2Xw8OImUvEAV/UoPy+tY
Z9JDtd9lBdPA3FBxvJytecmvZax1ei5YyR5YUy+DGb9SgpP1Kw0JyPlM1rMYsz2SZcLC0EMYB5yq
REubjzYrK4+bAXDWy+qLTH3exug5hWl3qOJVQH9jSJe8Bm2bSD0IMNYh3DN1jXr0k2P16v0eGrVD
6LA0oUDgj4DdQ4oGF30zSt7aKDBQfd7ANfq3F3zBrMeei/gg1uX9TwAjNmsizNleA4QwvQ/d07hD
kigzWaG9FEVjfYYCC59lljJTrK0Q99I3OHh9O22wWYzRyIXR/n2uWZ6DFHKoyN78fnQGEdfzfFLp
ULyX4AirtMr0BDsl/fd5fUxU7vEFxT4R6Fg/HtxN1J2eJDeS1YqSsH7fGMlwYihsM1HA5WSfN3vI
lWZ5GKcyTRf6Us4PCImSItUZbnlTW+nr7MHtsqciZANzfWxoIm9hHgawGd7Swaswu+lExqUK535T
54826ZYX8M5LR8Kpgg4Zk7HkaXVNGJ3kS1DvQFQl/DLZWHHOBFJ7TTPfJEcNRLmOYIFtXddL7AvP
NUsJHihYRXswaY/DaiCUzn8y4FF9+w9zvaUh3THA/xB8YaKY2LA1R72KnrKu5aJe1lWpqhcSkU/A
vzrlgXmgRbWmmtSTjDVa03v0bo6kI4d1g5HTSr3LeVrcnjI7grfp2bWqCbHi8NBg1K+2ZU18ewcc
beKPo2/Bt/Cf+vkBWpoZohT3kbCg+gqHzWDTFsle5BIAtNX2Uy8o9ysoPyBZJhGQRdM7ZD4YmmfB
fbw5p07DgAiOxJshanZ3E1HeuBdthDBqQWTniQ6IFA/hMznPuCOYF17rahmPWvWldGwDEyKB599A
I8ph/4OjYumHSHa36c85a2T/jAH4S1uN4rAzjCHc/DOjWipt03gCFHbVzH+grgVKxgaVyzyAz18e
mP3anMoYuRx9JQA+WCiWji+c3nGlpPUAdBS0YC6rUZnLULveR72kdy16B8DBV3aAPL5XQQ9xszzo
HM2Ey4JTO5/NwIl1wRFn7YB0WJqCnoeGgOdVM93cEq0vKLWx0whoyQmgdSdV8feCSi2KGo5aPp5X
rnptzTS/bYKnj9iPobYm/DAEFRc8qwEhwxiBrNiaRZAQIY4N/bdsGuzHeNjNGf0Dk4ewa3ecXxly
Aw5ijxUBdT0KdilYxjKW5mB8s0uIEbySePKX6W6TzI/n9EnFKvA+kqxP0cieYCWRMb8jZKk7gi99
BADeJlsHYgbuLXpaVDIF5GmtG6PpWsKPQuf8vxI88K3qS3SzR1TCSDuaG2fVHFgiyQ2qJSbltzT7
9jjdo7OUXBR+1Ck+uwNwfmKPIeddNQM8KP7D+/YjtHQqpRjJFd++jpkfV7NrSEtHkw++dRQ8pmcr
f6Oc3vjqKrQBsjkIJXnaGwWCK9/VxFMXBpvwXVfQk9qeQ1Eftfnu6R3BDQ/qEFEzo0Wgo5SGNJG3
STg3PbSoxBW7VY9NQDNDWPCzj1dOQuTLzNuM1KtNFyrLsH1YTEz7yE4NnWFcw3Iqgt/WDIE65L/v
B1VYlW3PnWF6aWiGPLCk7FY8SGjExEFrwI/bdHe4ilDSLHjraKkzRnd6EztKlGaAgXTFZaduM69E
LmSDkn0PSV+FLXuUpscUk/jNAN96usZmwZDdb1P38XQC0A5bQIKDEM0Cv7jzXxdkt1rc15QIVn1c
iIIoPUn4IGg6NCOf5RIdVPxdrF6Gor0+sAuVf/HFTBSesDgoUskSvOiZpMffQxfCml8kDgnK351M
pWwzvfgZKe7BwB0pS3j9FpP0MlCBmKRP6TeWpvWJiBHUqCRARD3olxV1DS4XDpGyimh0wcwovI7p
gBdvjDQNxHKQL483ImrKz31kszbjRj+jIOZo6b434JGMCoTdqtc513CJ3chnp49FwlbzHTZxLyI1
fAM2btb+d0Ykxbom+0v3LTXrve7UrvQA5grcklpQ8mr7aX1LL3ZJifiAnKiWe1a3wofh3wciYHUL
MNpYBtEjGJcBFDT4ueBNkc0z4sySPMh1ztvKJWx8dm5HD0ajD+vEoSaG31/ZKfkbCC1heUlSWpPN
Ms2CUKAmoeXXgL/OE5RwfJaP8OkGY0eFbCNgFZM5BZrMVdzKx/1D4voj4Ik+4UZ3e70GlJ9yz+oO
EyCgmZ/AkNesSXlCidMfcluOXXf7yoI8A9ckz0/w+QolhUOyBxW6g9xWQFEXiY+m1fQfmNqGlb/M
RVcO44oIUkzaj2n5+JJcIgF/+iB5nh4V06QjDju6OnmA/wYrPyGLfzfmBCDtyCGLpC2negBxSDRC
DonAdCuJDdLJkQDlsl/cF8ZKtnGl/8mFWzxefR+R98WZN5GolB9l2wEfBtAhV0kCIWhS5Xkm7GM3
ACJ0wnzIv+MtZkrjwaFPKVoqqE7ZIpvDGP2Ao5RBqae1nUktNGD6lRS8elD6YmrfZThMqwOVK/pz
BQ56LUBGX1hJGPocL8JJ/LMfg3gyB/efRiT9p1h9bX/ca+fEOmvRbiZaha6jSSSwDriMdNpmHw2v
dJu1YeLUGWv19zeIt0YhOKQv6upzHhu4Zbol9/2kFKxfACB34+peXiokFXeVAdwu/GpCp0QIV0lY
/UGvd0e+Cy6nzrA1RfxSLMj0bsidCXd+ByFVFPSbNurRpKHPI3qeD2M8BGGzWME5jXscO8zXWR/1
VpKE1cnWBTpTX2cd+3PBfQXHSDiQeod4X1izSFTE8AEK6t+KqHOX/bwtYhcFn9GED/nfvTSy8q21
ICHAciU4dZxX2SqfFc1k9Z2O8aGPdRHumZB0d2h/hrTJzjj+D/nc+gOTi7+lWYK5QmjyH4HeST8+
x0uXXkuzLeuV4MobKiySJtkO0FQwQ+aUx34XFBJPTqSub0ChWxno+Hrj/BAq80V0n/BZdNlZs3kP
gvmO5ZwlSxh80+SluekkMypNEW5IauMpNbpAJQ0b4a1tHiKQTGfi6Z92yj4WKxA/42LwsABWLXRH
h0B1KbzUKGtLC5GdA8S1fwPf8wDnbr7LuiXaZUs8sTJ5V6qLcw0fhHCpKSeBnkWeThoGh7hsU44p
FQknjrqjYFiSJ7djAPON5Te62lyZvH4TMJjAtxbA/Q/KnLzCXk7zqmo7cxLutum5EhKIrrpCwnbb
TET8TG6T4LgcnT/L0xy9mrXb6S0N+GIxIYl0Uq9fQhURiRLgOA2teYmXmGL0JSho5g0VArx4rZeB
S/SkvN1ZrVG6h2pMGFYyaQ3sh8FARvFUeGAwn9iIQPI+2WatACMXzg15SihuoZQFWqZpQ3sPOB0p
KSa2FN2cE00cdUQUESwD49RDFGAgf+mypB4hWNJbL1m+FSKz6oDEdrtxtHc1vvgUwcO7mk1wpVzQ
7AHITwZopoZqGoNEq2oIm43YRtIH/FfleOOLLensmtQbIMqShgl0UspxpycBo2xy/kFob18iphbU
Dz9/nEQW3Fp1TDeSiUVB8kZjra1dSp8X9nZERvdKxvQ7d4kGeTmV0N1VkyOYD5x6cJULMqSKffoG
VS0P1oOPYBrgMfHQoGi7DF017HXd2qo0RmEBl3sGvWmhurZIfhaz3AonprnC1/pP3sNanNu3QWnb
p0kfwoCkg788EY85wMW46et+7T60W0Zn2JgQuWsh0bora4LtY6q6p4WN2qfDiSklTYCSVcQcLiPX
mpjApjyFcDyRhTqITo+gLkc2Zk59xW7xCxeUka1E7+VACKykEb+IzokHpxvEDF6V/GV561Ror3lR
xhAxYN97KxZh89MblNCXXGwXmA5qH9k3wSdNmQSddnNAuqdzRtp65RweVk1cJ5rjWIb8Q0qERp+5
N/qiqZCixn5oMtNFDO/q95BkC4rLWlKj0sJUuifqjtJdhS13L97VGeLx0VuCam4VJSrXJtQSSWNX
lwTM0POn07X4xgecYfJtfVF8y804tRzm0bThSU8Wy58TLLwQqeBIfClpaSb/yjiHOwAjem0+G8ba
OwpYjt5XuVuIT+WT0CEvQzJoqwKFjFApJKWnsTkerjVa746fwotaQZRcSZHmmUO5ISlZSRQAef3c
uccbB70SLODKDyxKHzKz4jx81VPuFov3Vbfv/48dkus0pRFAuDU6UZLuI9janjo50+Q6qA2+EEb/
YeY8r5DwrFFzTma11Reg7a2tyXgAKkUjTsSQT1EmNpgwRpQlaWsneo8saCe9n2E82lMFScxS/Mja
HSq1n4AeptAdqm71YZCvVhL42dKAM07vE1RJ0VFMtdhrc4m3cFonCSdW+yS0xYLvcH8u8cq6B6S5
nRShW9yhQjlrxxyED/l0wrDOWMJz7w+WPKdhumH1qoVONJhxrtlvMNnIohrXr2qBwIJHyI/omrQW
o+bIh5C88cDx7ttUK+94aptslln8RXmXpQNaRX5DDqQbI7HFe0yDSi2jr8SXD7hQseYx4Du2hPuU
u7ZnzLXWG/8+KPV2zGAP+0+40FHjacKiUlOfkqmkKLHka78pmIYFYSaW56HNkdzRxO/Y2O8qjfG8
f+mwOLAUJ+AO9VwxIhLZga9BNso1ibuohFzjpq+LnvVa7xbOeSI2uMsd4zeYBEtyQ1Cu2j3SNPp7
/dXL04SyxKMAYJelEreof2mu/6BzmhurVS+TyRgXBajQPtTOfsPJEjHpEzphj0+5q2A8JutbAyMq
mkI6CR0myuIbv+ShguQK5JudfYyOARu8da82INCh6kpm7KoWcP3Mm86fm/A6t4x9oHpo5xAMPS2I
YHbU61bxrxeAb+/Yv39J+jp/Y/ycJ0piabTVw9lnOIaHgyqcuvmxQ0p2Hy+GlF7/QAgTMKQtNrT7
hqpIC0LEijQ/kRY5CFxeoEhfGfLgJHdLCPa6Uqvfgh2Bg5DAlcZWmBEuKhyWueCOAxtMmxDCWika
euDUxvf4PDySVcnuFI7eYaQGvg1HZvQK1PpX8XFB3miKYlHfrKm9gUdQ5ulCKxowsljeKuPtVWZ5
8NZeOs3pexskjN3nQnyZb5XrSe0L2UqqEmEB4negFRGiB/1XeZVGZ5Rvq4QjkcISWoPDrT8865ak
POj+3aW+Dm8ScE5lA/G5YU9rR7kkau3ngyEDhtkBys3HxlNv97TrxA/pgdsGg3vhPJK9Pq2CXkVd
7TFWdCjPs+GVCWx6wnKdGvJjI8lnZrC9EN1dlUn1mustPx/fy/nR6EB5W3FpI6o2ab11vPUG61pH
S/LfQ6vA1tmuoNDoIU7rIm1qg8vIrc9/M8uVyX1D7eY4M0kMqnDUSLTxP58AA2rGCVXc4YLgjthJ
dqk3r29Epg71WmQjX+N64dXztbrWwti2DWuTB3Y9mllYgQKMF9xeU30z7yF/w5SypcpRBNdiYI8y
+nzC8cVfJULz0Yt92YFfwXzdbJLe6JYc4JsEPwDbILXCgNwrO3MW6DTkSdtHW21vjZd7TPvvoMit
xCMEzDcKxqs6cn3n823bidnZZTuGFewtiZ9Ay41RgclRHwAszKVS3Z7Ht9Ji/4leoL4XrZobsjFq
qYotBUMqQdkZf2paGLnCQ06wrY7HsehCP4qvZ/rgjIibr4ERBpTlPj7Qw1pBxbdJ9ql7ywgZiaIO
WrwcBZZd0Iv2QCwtHADK0tOvqFVt2pxMFl0dE8J5OronD1q8VDEZH0TyJrjiBbBdSdrLrinAYCoN
D/zCmQhcUT3b02VXu+ZmUDxHH9AFRubbkZA7DhYC8TvvPreXMVZtUl8nPvhDb8sQKdiOE8wfbp0k
nWWcNADoKLHHTPgkx/ZeBrIPoTQ6xRtlU3MLjdHbOJ8IAqxawvBuTtVYnt0BqkELV0w9/RvSnNY5
Bww8+ACjSG3RjEkVt83o5gYvhfR8hac33aKvL/43rbRnlQVZ5aGTU7PHVYipKeb40E0xeJTr2ydO
LzQJYsyWwQfa6V4uonB0Bm7v63QE3QTSLQE/uTJg+LbxKWcMYfRdMZC4kAWSVvZZ7F/pRsYSd6vG
ei2u/8dEqyGcs/Hb3F2nvMy+1ZSsql6Y2EE5O4Ay0i6f7HzlSwkuR2Ie1C0dNL4c+IVKEAK/eN40
yBEhkjLjqlyG4zkKvnCiP2cWRbDLSH/wy++CU4u4vdf1XtNifZlMYs5fTz2DjyNruLXKJrDRpBCe
HU4RtJZXCsbUHjDZhftIrVdktV7Bkan3AkmbIuayaPyjO/WIJom1QzNWXBHZJlYuTLSfM/ZPZfhQ
ngoMDYuwVt2F6SZepzBgdRLEi6+f+XHDfjvOz/dP6+/rEAHX2PTog6x8554QWcqBLdW2QNVhDkyL
TgOpgijf6gF7p3lXgEyx+cN6NgGB612MrZztqXU+ZpC7XZGemXeOO91cmF1Dm13YZCXq6+WR+D1d
xqQ+4k4Jl4MPXI8mui718YIUZbS5ub9pgSTtK1b/K5p3S6ca4ndNPM5gN8Ia03Y+I1jDBt1k+zJY
av7k4V8gC0/zRd8ECSHAZNzUibh8q755LpfnbyLeEqySPONhHKu33W2dmsB3Eg0moO9ZYas1xRqV
uBhk8XxE0/siQwQv9wfFrBNJdiB80pf0vaODAreq4gsUx+rt5yl8+v9MqiPWeo/Ifbar1a9qYz4a
SmI6cgW5vrCvtSTZyjwyzhTtEDRpdr78Hry+GcnrOPUETXVTMAfckMyYCUUWrMfBTH4GHvN1ykBs
AoZ8/zgwRaE388w12pjj587HgQf1aJsGiC1TQW4/v+eREGo8rtchLfAnDr+OQ7tgGiohlUqqMA/2
aaXmyrj+JnbHla660gdVQQEW7P/abz50lwgSJodRfMb5pNMpDFyydvUkESThdNsZw61t2YtMKyiM
JduNfLpVyTUhujtDir/7CT7Mq+EoL+2uLPmXFNXli2JjRVObVuJmp8ApbXnZrFdeP8cuiE8hzxO7
+cDHHklxbpW9GBbyR4ISlud6UMztoBpWbEKqYQgPpqytVykzT0JeqOqpMf3hQUB0fLMiavBYXnHX
IVt7xPAlNSxMd3fOGlsPM5yY6qEJeeiCbWf7RxQ145opoQmYAyBXVVMW2zxBfUA8f9sK1OvuED1G
/BMeyM9pfN4MgZTMqfKu9xDRzfZ3R8HfTdhJZMupg8KkLH85Pi4/Lf/QMWkuNbgYDqB7136726lN
Z6kXJS0RLAwIuyVNp5mUfcPO1TRpxJrYRi99pfqkKMPR5vsvPm2HTxoV2BbAmbz3p8uwtHAuwydK
O+kWZmhLXYlvEStLTYF6r35jTL6RavCuIVEHIVqEpaFuGXNE/4CMzN7ljW/jPCwyfYhPk9BU+nLB
NIwZ5bb1xMZoNBGb6hYRq1MK36CPSxUF4r95QEeR2jEPXGC0f0tdqEcmaic/I6GWj7Wtn9sunN5K
uMuKf86VQAoAg0peraVsRx8d/jcyl9tWpSfA15Vhr5a3jeyEb3NormnnbY8T7pDk8todAkAwPTZT
Ug40G6AlIIEzKxzmZfLfSA164Tz3g4Q4AxygtQ+LiJErzj/NnRjWnoePXh6TZL1UpgPRehthlozB
hO24zPRtdPCn4Tk9cMH9j81QrichZ8p60r50KvuApIwJ5N/EeRx6ZPLILfYh3feI1uUaltO6Ctov
1LrnINQtVs50XwhNLpKCk1oL79MOw402sQeeSbyr2fTIVOiXpoQqsFBMdr55dWhsKZUaNMt6IJih
kdoOrCtyAj2DtfNs5iy02DwBdu3sTu1+bMRmu6BGONf2aNW+q/Jbq6x0vy9rINyMHM6MR69Sj30Q
HZjqQ6bAUn/Lyfq+Vgo3mkufbdJDS5RMftwUOiWdVFfPYUyBifeVjG4GcbQJoar2Krf1whx/MeGO
2z/HWfifrVfKv9YWTC4bN0lHDaRueNIRr/+W36/Sua+aaJWOZRgOJ7Pfmrp4uSoQkwDVpKryVfBM
8loOIl2gU6yaawotZsnldjAQRCRams/2379jcJxt404bgi6g2OX4JSEKguh6opEedjimza7NIB/G
7bmYm2UIraAP/JT0Poctrmz3oWB1WdLPiMRV+zN5OYlh2m1l1wRqxBazHssrYsVzpL8nDec3maHx
mbF8HnAkTiBHpRlUQkCezUryIveCoEwdeGUz1BJyxdc5RpQvBV8FWhhem4Mn402rzsjVbOrzJ0Zt
YU8zeLlPUkeerTMcFiX+mPTUMXio4Ss9B6TNBnjfrdBYSCSO0Z5j6g6+wWYRyyQPJqnjn563/SlF
D3KCn9UhMIJpRFjlWhWWL8WkOcM3R5oz6IBYbcZeAVZxX7a0mWaCawA8brBNHkHXNralnrmZCdX3
17v7H46fTZBhVS2tdyHlM1eO8s6eU0d72wvn8/3dMrmZG94ZcSLXzi8ng7TQFu+Cvn7m96+Ps39/
blMWsH/FqhLHBy64JoAH/eo4MMUSh+U31y5vBoTXEzDoRL9VHrLMe4a2cYEiGha0P36z709vL6Jo
mhbfG+F3HS6U9PTa9r5J8kXW/ZJDEeZRXK9+42EZ884Hg5/qcMoVRVoJXK3nRz4EGEPLIEd+aqq9
Ll0k6v8M1P1j/g3EYG6e338g6GypZC8H9Nyw7Ynh9QqNFhb3JD6FRAsu52D7cKR379S7Z6OkUkLU
Mgoi7MVQjf1DbYJkaIdoOIz3QaHbl/XYB7NkVTvv+aPk7/f2F1rFP63vKcrhzoXauGnAcPvIQayo
h1ZZKNmfC87C532NX7iw/5R62Q4PPo4FaySB4J+jcD0jXvzuiTd6lT2tvFa9F2k6R+VlZuOn1QLJ
MwmqO4oQuDwxGF20A4WQvKD20tHTQF1oPtmQW1Cn53fMtNSIMW7bkg1cXRP9iq9tlyvplxfuAAk0
aEBB/OKjeF5rgbuY08mV51UcUAQbnq8FYFtxEjgoaiQrF/CgnkZnBLsijexXi18jl67Ar5j4Iret
7OzLzKuE8/eOB62AeXnn4b8PHJ7GGrfOJ4mwOLhx5PGpMa6D1G2L5jUYWw3jGcPbNDoQCYo0ElQe
AHQIu9/og3iOyzoyiiyjcRgeSg/8nCTfu31/xENt7Z4znru6/WvGR4m+ZdFg8FHJll9Nuh2QX2Z4
RwWqiXNweW+0HLIQZVRVPIYj2WbBhUJnBDt5MWPdfoTQH6jqZ80w/zczDLAAYP36haYMzQuRWCwH
jSE9nvYYfjIlDN4piX+yh7A70Oun4Z2vpfkTMb/n3stzLswKda1Clw06/uYsrj3ufWAwdH8+Pn9r
AoFfdJlMY0yo9+8US0mdxBnSZlNbirgnqeaJw96CQdnRKrxmGCjgbhxwF3zJavu39A0iNC6KWm5a
co3UQ/iUuNa0vVqHElzjdrJBH2Ry20Myadrwh3UQga6ipTK96IvAVkAwniXLp9XYM106ax1riWOR
l1b2xHDjTKt/JmI1OMVFaS2a5hpGRup93uAScHW7VdQgnaKADsTpSivO/Kr7LYUhvylx6D6MMqdn
DdANkv3HjxQrHyAtmWcNQsu5VPo8I2VeN+oWuLqLr90Id5IiUAObFKfdoFGL2N6l18bmEMDmHfRf
NsQ2WxViuckcuQoZyikhyUDvx7QcEnxA7ElzqddLIy9VQGkPSbXixmJc+fX2QNsMxa/QQa947Mmg
LREgyRtHECSIjcI65StQMAJ3Q3LPENZ+oYyNlYWQUwIJeuksRJPFNV0CIbx/OaITD2QoyOyfdtsf
z1qy6RbwFiYty0QtZEzTfKMEklM8VmRR7VPJtY56AtH6ufZPMebbHdshFYryIhaFJHndDUdohhpH
eCopMOx+akinAj4uix7YQEkU1ch3LVADGu8/+Zt1/b6FZRu2+UtFHYErE3qfpdDyiAy2oBY82GEK
1tgTKIoRIfCQssBNYK0E7jvdu0uOBbla4jIKYSurBMh11jPDodsTOwFCjT28hOlODwrsB0Ih8v8O
n5NtEKR/tNbNgk3rsr0RI9Nj1usX0ghCo3ool+wytqfhiNzdNZIfVQPNv9FzpLhqkEj51/DoEYc3
P4nIuAvznd9ZXfch5yw2h/KSqoRpLqt3cgQ+S0WRzgjT6N63MRd5zmOsLse4AzuKTIhPVRAdnynL
hbAoANn3mlxL0Kg2swkCZcYhZmi7vePfKKWrV0Yco2WsGpUuMX++2pvEcXf81VPdG9x6oGh8hHNg
5WXTY6cxqhA3wWdn/wZfPXUzQl/h8DS7ogk2VsNZIKdK+D5RnbK89FQcQV2uaI1wOP2DM+RGxWF0
s/cwYkYxq1bLPuZtEpgx58TuPRMpMGiAHMHQMz47DTK7dxnZ33ujc4zYXlmSlk62qOWQ82SfaWXS
ioFxVuPAuJOOOav/agWAVKqC4qtw1dmaeBPI4tdQ0fezVKSmMzW1gWn7zKrRyhaeAOgl6jVfSESj
mSNRZLgsXVyNFzM4pUi8+7t9gcFXUP+a/gXUV9DhLSIltukDUS9OsQGJb9f3bl6cnY2NdndVgHMW
DGkbrWjmTbaEkOnbhWVt+t325uSb2mY1GgLPRvwiDgwLJQBk2Jlrn9E7n8/z8mfYPP0qsXPKTxy9
hzEjmfUMdo5mY6wweFw/QI/SGN+9LxzoJtoem8YsibmcN9q3aZa5CHlB7vTzPgiw/YVHQ/lW1gq0
zuvGiImY+kigU5eSrDQ/n2ChTwCeUUcQjxDzvdujsIyxJgjmpeqzQg4HJnRLrdroc3cbnzXZd0iD
Y8JLy8WHBTLU493WxGVRToyAy2ZOAEDZR17QTupF51s9Ev7RKq/pLw42hoqXbXxBMNZddLsNG41l
c5LHwjSwAIAo1BoEBtMhHVWF+yPU/CWeXC04Yp3oTgmEV2EhPP9SfexZBEmbqXRQLQnbPj0rGpbk
SaC2aL0S/FNObswoCQa3TyLv4p0K3+buOUEPOJ2+PUUpB4WEdmMVrE1uyyyfbh37cIUXlgQqng8/
7sASgF+RcK6xmHg1901hI+0QPlLYQhkxwqG7pznUIQDcVBPuPCaR21PTvLmVZOjBNUjMApupEReR
OeAAoKoKDDdiA2Rl26OZq6H8LvcBtwOKAaDDSLCuelBXTay6kQEz5Gyx8T4Jk2d/bUAvmmOLtRbv
7geA2JqvicozIc7PrKsPxDWfskkDlnI6J6fc02kDMd7sGvNcUMEihbFpyvlUl58hzD+jcZrXc7jx
L7UZ8zSJKmacalaGKR7kRHF+c2YmjmkqAcJOnyZNSHX1T5omjZhrp2eg2fCBbyzrNnTmpsiaiE9I
VjwkFZtthwbodT+au9VD/xD7VWqyF8V3KkOi1daXo9gaTN+ledb70GHIrGBtujHA9lwGIWtj3Iep
UgEHbrxiGlXUlCZ2ZQLxGye9EmAbn0SvUol/M8khS3V/VrGia7E9ZxdKxyo9xofVmahiv9KZ6XcM
vYo6bUhmVU1wyZ7XWLMptCMSzIOs8O7eDnJbRDGD9zymBVujiffnTQyPIMgBXUqiIvfaA2AMk09F
HSoE9aIiIQVb57/jZjiuNCmtEeMBBOJBY0/IFt4uuk7bDgDBLEIe/i2x2bZaimYKkSKctV+a3osz
h8dDuVP8tgNJVNFPdv8MxxPStzjTWc7YvRxMbSY1CO8+thU0DsMCTCXSKPq60jDs2lX0WdAcJOVr
OU4ZMjRjrRiz6ZUOUm2ivz6oHlsJXTabtMqK9G0c/Na2hyMhRSwUpt3u8QL5tZvygVDCC9HbMJIY
vSoxEeLUTdv6vg6YiyV+v0Bcd2HaO2oysTZvholj6No1KdSpJDZnBNLL8zrId+fPIL9HB3BmtR/w
ETD1rm73p/Q7IdBehfjML2Z4k/ZS6OtSJgH6Vod3fkQxUgH62AEgY7Ths/pf6CYW+cbHNbCv89CD
Kqp9o8aQF//DgN/A8fmx4O4B1Fg3XSc/XGG7PejpKlajyKTTHIGJMGlWG+QUlULIXy4pV4qT9IyY
2boGqooquz8nCGr4ErQXZGmbS7sMekeUxgBGJTfitk5ev/xiTYuoA+Vvwwz38RXO0Q7u6MsrJysc
zmO9enhjnwbL5FX3HkO+Q9VAA1ljCpeqy2y0PXXrRp/O0T5hQdzAurSSsa+HLRTGRPvu0KNy+bns
A+XAx27IlOOCNwDg+Oox62zDixh+Zz4xzdCv3CvjJ1V3aP2wQKZGdLajwMWplH0nmLdbyGHUffA9
aXu+CsbLuRuB0zZrSQXRMl0w0yKm5y1MvT06OUP0JZ+aXyTOVV8oWAxjh5aTOS2iMkg1OJcYEBFJ
WTeD6ulNyFZzy7LZFXs5W6/3qv6Zs2BxhTKL4Nez3HSgggkPajwegXL5zbRk6eB73a7I7q0IxB80
NdS+PrQ9fMfULTxV5iJKJwaEuW3JSm/9jCm9plkElDz0P1kZTJBNLx9OWZdJGE+KRT4JnooHkVM0
JZGg0TVWTwUOZOMFgUTcHFe3vDVfNgMMyy+NWGz/66h1yXFuewhedqGrNnYmX6HlRLxBHLFNEUvv
pS3PsKSpzJ8NNX+1lMrpNrXNpubu9QjpSFdZIvJe6ww6xf5j9cF91gPBrJA17oj27o4wekX6lMwr
ZD4stnRVzATiCJPdVm5ZxtCyq9uCDbiG2YZ/Ny3DYEQ9k30gZ0+R6sqCIGk216E8HD2zOKM0fwc7
jIBxQ5Ii2NZ4w01bJIV96cJ9KA49FXyBl0beufoKaEqh7L9z5/l5IWR3RURU79Lc68ZbJxmxgl0t
q57HI5TPJaBw28ktdErC0e7z/kwVoMgblfRYAbqc0r6dw8EynsOGv7fjpgNrXkyJvxeiCY8zbtus
bzHcd5SiZnW6MKp45mMI/rptqMkcJv5TMOwatVRuGW6mAfvZzCHaJqZxwk/Qi8ifkl+7aTLvqSXA
U55CiLZa8xEJobbH7o6glopaF7y0cLRg1Qp9zQnk0xNwO6fPIDo81Bz8GNoai/01ESWFByT0AxbX
nxpyQxP/q6VOGI0+IHw6R41x17GczS9ASiaNmuQqFDq+QaOCQzBxWEG6bzbLI1h7VE798z1BBxAY
JZY/74nEfcWhh5zFtsSeK88kJisDvJXXYtO7sKbDwFF6X/GMDw4kA4s554NBYgJpOIhVmYC3xN3A
KjkkXFuvmb/TQbzzL1pHq/M2a2ipp/rgi2+X0lbyT/s/8G+2Qj7osbCUotlhPu/QDew2ZriqndFf
yrxU3Y8UxdbiQXe8Fj0X0n6voM/hqhb5FUPIYM7RUsRqZN6bYhd2Mq+kKblgLf5u/cm00Tl5BH/r
qHbI4F8MHHYBDQfDbQt2a2b4Pm0eqdktUsNnjgQEOBlfY0DicYKHRwSDjjmXRldyvXFpEr6j4/F4
PxuDOPp8q6Er9NRv9rcaPnPz2p3s0R3ineMwg8wjguc8zy9YWY15ZzXTMxBskY9K4n0m9sABrqf+
W1p0ctgpCmWs/VXbimha1kPQk7OWyExLKplTvEH2jR8sfG9ahqzajI4tdNrVUhvZh9+r1Ghmplrq
cdZ0uF3U1/wE6t2f3yH4B3INqVhcV5islGFTdVhrtEEaFwlVmg7zvBP9e9sHg1Zj4LYT9fWPN5E7
GZEX+/pJFHj9ysrN/Q3VFWZhA07hw3h9RvZB214saaTR73dmoTJsiGbrgInqF6sOLmh8xQsjMEsH
7+i9B2si8WzJHUYdwnNwthQqHOOnbmKeNT1Aiu3RnTJIyH67/1Udc5kiJeP24kHGUn1A69DTypp/
bnAeP07Jo5Je5hjri3njZ28q/ox/YiDTpfYP8K2RMNoeshmgfyORA51OQSGdtPZ8ewy616PB6pEc
dMH3rpG4LoVTeXlPJXPmFRMGRkzM23/OPcbnA4s802hAOML3/LnYehSyw/zY5BgjMd0uZYsaX2QS
QqfuAjoccDdnhZqh9MyPpGqGeocmaUd/IM/7ssWuayRXBrsP29QqafLv6qcO2PsqFe7p614auHUw
z3dyoP86S9XqQ1NJsINe4HjyDFPgPGmW4kpCQO1t4G/P1DtKjHqcd7EebRP+p1mu9H2SpvYrMVpR
Vk1K7YbMsDNEAuHsd9jEVwY2V9DhnMU9heCcEvf6rE4CkTETyvG8nTtZSYl2xa+XwTGzkpNU4K0J
JF6dTiMRiui9io+FBQqThdzcOGRIQFAZgqsyLcm+wGwjG0ClNdGk89QgA51l79vC4G2ZCXh5PEDm
zqFfsbx1pVTz02KaFfgaLgDX2jSWHKtxrI9FkeED3ClZUxtt0iOkRVold6IEXFj/QE7N7oZXnWX2
3VT7HW+o/esQprN0rFFzmW1pTkhEUaHRgiuABq+3n0Jw+fpok1mXpIDuaCtje1OGQ8GPNJDRUrNS
j7O/5/oZuDtQHUUinXpqi/7hC4IDIdZGkG8zuEg/blbH9OMq7rE9/YkbX8OzQ7GjYZ3OG7FAOtTY
vSEGByT99EN4eUFiKiAVlrlv0qovbrrq4LM3CDzBz6qGhMdF4QEm3iQ7EjNtbR5Uu88KVWEHOyzk
ACSC4zFpKAtCowmOcQsa/hBeugmf0rrYb9jLiKCiDUdH2BaH9GiJRy2N/GfFQHlUFosA3HnnCRhV
V9WCRB+TIq/+B/n3dy5jWIib+BSpYV8/mGuNldETZrVoAETX5z7CJ8duDCq6Pb5QGYGai7549Odg
wxh8njqEFrPHnin/+NnJdpQwpl5sCfKxl/SSc+wjxFkhUTAJS/h/AQzK+/tHUxsZMpmc1a/mQtCI
YlnkS3Id7+UN2q7RVlTATT8iiNnHpXEiGw4mgFQM94phjqFo9e+/mEWtFCKwnL0+AK0pgGvkLEKk
ZsbhfFSUf9OVPM9FJVIkdFgIIAHxwTWt9LJ4wbs2WbJvBjwKOnYXnvWPQmdmSzAHlwOIWrS/NYs7
zeP4PQUuTOlmUzDJPYqkvaXsObMg1f0MwAPuaHRll8JEU0f1qee3at3ZBIstyozVfYIvTnbyDcGq
3+eQMR8xyh7byOdfQnANSREtFXzsKjEAiVfpO6QYJ+Tlx3is20CU9B5F3Jg5A8xe9WBsQIVvfLYq
XAVOXTPT6F+y/4fWjqry4FaagnKqaSB5PKisWdX8gjkzbpLhIysOBwn21x9t57/KWUuUZDZ0XrZg
KRoYBmxEC3dvzP/G6UvCdJ0kUjxBLMGfivYi6X/MPe5CvGKknS1JiErdg7mJ64DXv09pfWsmaGKA
UGHnAgY1PuKEjXcFUfTK6h76E095bJnxs+hdO7EIHYoPFYbXpH1glHlXp86w1wz774qOmydwfAcC
HGi0mIvw488rpuxz4L5RKlv4kHkCh8YNXil6cFrGJRvyoXlu6woKmR/X3Dkuw6cI9Lk7whGT9RrE
4T7r3GoooG85889yJg69C+VGCe9EtbmfV5o6DQHeeCdGtjcY5hF8XfZp0H/5q+7+vkbRXf60439q
gFuNlXbUT1cZhitnYLQssDPmjQ+aLMJtl7a52vzWT49DU91UfAbFrE8TVm9X99nklx1Zwci05z5D
refLZMWInQLU3RZQ55MTycULhb4gOwt1uM5XuKUXYermaH+bzvMp1AQEdyEb2bkbow4IZct18AN6
BMmwVTJnyjsZIAFg9iy5vES9qSRP+HGYeBQ6R8H6jWYx/2mRYUJt28aMCguX4Hv6vh76styZTDoV
HWR3yo3kAj580jtCEqk8HFrvuvHJlJf4ifazdX4Tgh9anOb7aDo8l6mGiVeYXAFvqgaqKkyiow8Z
Thg4bDmBxN4EJnXk0VrpLK1PW79rpdnYkh7oDWMoNqsB15SMj0Ch1ICDyz+JZzsvELZNLMjdCEgj
dk2Qd4Y5UqSEnVztwRAUWeL2mACTN1TDc5xrGaIsBY6X6x2LJz0HMIjErex/Eqsl1SzhIIhQuiJS
ZXKEk5g1EevRZexUGw9hmLC2m6CJ6zxTQ5WIEWqEPe1e9iD2FlL/X8BaEmALpDEzCYa1l96wlBTu
VeBPkh3+ScdDmUrO8bcsqutvQ9VUtGnpRP0WtzM3ITeuMqsBV778mSyXPBWa9TZl2GQ/iAD2fuUO
v9me6rbm1GPMYqK7BSB0CqWdYcmJ4/IfntPGGJPOYiuiyKO4cuAYAwfysSAiaxc+ciVJLJfkBVgY
Hkktn35Cnxa+JsLcXfK1SpOtzJExEetWvBtw/i8Wpt+BAXnJoYMy2OdimgwjMRctcjYLT5hIUwU7
UGrTXE5IRTI8TvXYFSBPNcfP3dwceidYui9Ch8JeBvHJqlleQn8IypUkwxj+VDelaDKJwoUVLOwG
iYsSCbVbeQutnnA6glbBTpUjqIPZ/BMth8tap1G4bx42Xvh9okF7svZH6UMComOaMeuE6mGAuprs
F/UEmmhqvQy3udz4M/VkPCHmLmkhjpxraRYOgs9f8DXY9un8VYeTmib4naAV9VLq0+i8xeYWAt2x
CJMCSHyx6qF1w8By9/Vv9B8igK416HRLT5Pl1Ztwia93ruqv0wyGO9S4OFImVv8AccS0HYQkNYF8
rMqqNfRUlzdK2XkuoVwYMssxJsG2JoCTEbWoL3sM286V4FDVXao+LE57QnL6wgqzxm0nuCzg7VWx
la85hAFxQwmkmp2ro96xz1aXnoAi3HBDYNmED87cxiBFMLc/1qJD9mrDeIFQ3aRynrToOKvJOpzx
78i2vNBd49yUEoJUTAPszP28BWBvIdD61HRwdlk5s/NjvlKYpfqdL60FvTFxgD5yynpHCm0sHCki
W5oFxbAwm0x3iI2B75hl0KiNND6n789i6/Zdv+XQ5Q86xaqXKObUL467Rh6qk2vFY2ggfLKoXY5x
RSRVufRzs6Dh+FvRDFXSRRN4V5EfYWY9/9F0IzoPidMCdSipWHBGxyJ7CJ/LYCmozJLsY2CshHd/
pmDqHuk0XZitlPqmXFqVt2Yyq9o5cJgm8TkijE0jX4mbYR2kBdDYsFzaCuDu1CGFz+64zJuD6zIR
0CjGkXGwZp/b/ag/1fk/u6q6IZZpRn5L7Q0urOSCweWbPwlDCPGI7KrsapBZ+DIvuuVg0cuBD2fM
8pcdKGqH3wQ+292vYwp8DHjH0JpXIHIVx3FXJ0TYJYi7pKOXmj3NoEquTL5ejW3uwVwHqXOP3Rf3
WHZZBoBYbLXXPOYI39OlL5sccnx8c6pkk6ui0mMpA4rw9AqCIfNT58OhUd8gwv6kVtODKWMFOyI5
at8qPeIG02Oo/MwI3GqiP/RhcnV+NnEhe7FVFZBuWS3KkcyCd5K4Bq5ASqnINs0WJCMiA3xuAnD/
H8OWDt/RRQFxp6IfTqo/fIBDHO16iGkv35FbLSVmG6lXrfAmAVgSGretFo1ECPTgfjxs9R7Z2CVr
+4FYZ1yVL+4zZBWsEi/rtJg2/FEwxlZ8YIx+kTwJ0t+BMURI8HiS/OFQieXfuig/ZzZwdhKRX3dI
u/xXwL35kpJo68oUB5OMVDv1/cwDk/SKoQI2A3Om8BJbgUzDzm908qKAmZ1YlFWT/5uOtpJMcN9Q
HlCTuVMy9xwhQaICyMmJHHTENctuOb7CQiv8tfDfpfQkjjEBslCofXT3ob5mUQB/V2VpRwMUfh2e
qZUmH/dB67JLvHO27DKVFuCJFg+9vMtAJSan3ixK2G0JCqxmsycqM7m/x8ygx9+GzCMLoiDgz9Tx
eveIEw1VmI67lCUmNqPHqrRHWzWgJgmDTSGyrxhuIL5cPzBx3Ud8+RzsN21MKaCxovx65zrSw5hA
kee2wu/eAwvFUnkK2koEDeJjzYcqU6666pCnwgBbPBQbMLb/wzR7nOGfUJQ5FXUymaeF3UgP8Gab
RKGW2L2k4igCHKLciA7G/R4XsY+EwDuQwsbLlFwEbSoVTEpAg9HeMW5olV0etfWWgxDXTf4APcMJ
ATubAwBsJZ58A9+NjTt0MOlym5k4TUFkCPf0lYy3xxerfXjwOh7a1zLAVx/RULqybivoMXCZVDS1
0iwqOsSRkLyHhag1/gVPRpY8cmdnjEzFje3bRc1w5dYy4ZIsrZm+xC3ol3F4mX1cpXplkWyWx3G+
WjqdVCD6vk5Huxm+P1sX5T+RbfGhgmj6dQEmqBBIdhMkAeFq8X0VVoqtimo/E97CvyH05aN3iti3
rBJdqUIAcr1Gom1qAztRWxGmC8zjKoww6cjuuiL1wBUhVO3559u+YdbuOWRp9PONmnA6gd9y5FYu
LsNhpRKlyskuKGrGQKBz6voKa2PARSsYVbMLCljRDsgUe9UYqfpPfT2pqSNHpWHPiKLnrDKx4kQT
benrcWv04RYbQMKJnkBqmhJcqCiGeKImVW+E8rZWRuP0U2zQQfLrVTyOwVJFF/EuMRxdX4koKPs5
lwqUTRuqBIhTYSFb2w895tqBQCxDifCf795AEaeVgC3YpUkGco1Dp/AppJEyeyeQXGssbS/Qz+RQ
gWeoLHgns2KdlVFbC8G91/pJaeyfrgJltUJTpuOdDZ98AGVWmPtHoyq8jwxP/RyT0PFW7fHStR9F
JgDwTact9y/y0kMn933LMNcLpycwIF22geK1cZiHwrjkJcazLTUdOh/CWWfzk9gsTkGG8VfawWA4
RtiQCQdzr1+fXAuE2lRgSUCEaxKtT95I2QvCxY8i1CRdEryv5Zue87ekg2y+Ok6AOEw1L+ZMIJKP
VK0TyaglLUKREbK00m4PMwG+8vIrG2/rQBDC82aXxI7/7+nGLtkcGf7YtwRR0prqagUHH0Ut6gHN
k9xL8IbSGz5H/fRlPz41B7fJGp07TcQ4brTlIYXAX66jOev7l6QUVolnCzfOb7UdfsnAPs+18rCK
KFAN/z2KnIGDc6gng3hXm+zk+LYAt4eCeZ4Ab0DvVpiRVKsNDqLxdYhCj+hod18lwHnMz65nZDTS
3xoQe4mC2JEmisNKphdCcyrMgQVYlfYcWvfYFRwc+3Aube/TKfpISbIxSTv+3jB1y2lHmBJsHqHx
Qb3xOHdw4O2pqEFWzdUJDZvbQBBHPxGwOOU3XP2/PuDiIiR2wIV7KOXNxStact/n53OrOYD42jNM
kTElHW9lRNEZqFEwLr9JR4vOf3/fIlB3hkEZ5bXBlH9V5lgJ8MGoNu+lJo2rX3tDEEEFAZrEFzd7
/mHHi8fKtJJwwrz47DWxZR9LOUsmuUtnTtHWVinWdjkFnGiKOjwVqYV8k14qwolLgwC+MKhcMw64
Pghgy8kFALibEkBaK3peGLFaagx3Bhyndfv8TrOdPJ75dXa/+8yF3vhw835mQi5Dq4oERTufo/iJ
ZoqFyTjgUMz7ZY8P1YnZmiAo++NrkPJu74gLUH9gAGFdK5oZeP3Ar+RZz3dWcOCbvBPldtqlweHg
GI8+LtM5AFKsGLCgqh2X56Wn+HSxbQxk6wllGpie/lM6g8pYBCCHEffLk9xUv8HxHsfauWgyusOw
7LFD8tSboHVRatX/Ofw12N5o3p/G8PKFKrW1EJFRhisgZCqpCMi4Q+njMbBltSyzqLs0ml1ll0lu
6SsvFCOLQ8qiK/+EXukcfJuF6C9+cZPbbpBEmwOLClMMWl+nVbGHuA8roQtKo1bw6Wle7K34w1dy
xxoWCcXDExQUJC/IbJIZc7iButL/XV3Qh6H1QeScY+QYmAjfhufR4tWW8utVXNYxSt7PmuAeANXX
1Ska2wXG5SmNKNuaWqqspuQY32QcLpyyMClkYw0G7uuj93OT9evcz9aH4BOjgEQsO4r0zj16PKLk
rvdh5Em4jfFTbrW8aK2aNm1p3gp/MNTufxSORfBXPMZOKBR8ZC14+9Xd/wCg0IqswjZuFWpYX3Z4
qLZqJ8V2AiCBMhMEZ8NQIn5DyV9SyltI0kYDxLDtRG9/IixZgWD3G2qXPiulNXmy97YaVjBJYY/c
4BqgRjvjt5FXf1zTDjv6WvLXp+Z1BkCs7hILehdf7++7lMaBwE9AymF9ghcqDwe5lzIwgYbMm/eS
ie0IQ9E3PV7Ha3FXbQC/P/A4TotVcY7JLoenAh92UNoNA2w7laUR6VMN2BLAx78OUv++uQq+v53b
Vo1cMCHVFSEYh4o6pb3df2JP+hQ014ZwzuOgfdstdn3QXeVCIaqgupiZgkK5bLlBndGif7liXLGv
EgnG+KW0K/1p2V2p0ZAqIJRueFik4BaIF0xkZMbxSIxzwPVVm1b69s1KwFCZuHC2NBAmGwyiDNfz
P2sbvNzlZ0vzfB1bsc7dnBYqMy6x7V/9tEn9oQFl5jUQp6Mz8exbrJjDwmxvTl4neC0lR/bpY4dj
Ol5NGNg56Vww8l8ojxJgKDJgEDG80GJIyeEyBKbGr1Nd3JSHjGLf5ibLW5nse4DkS+zOGg0ek2qL
uLnZ64QXBOSPxoxSmrfG4+T5iwyFE3SMXBYGGRV/j5tRfbXkeYdPOjnOM25aPgsEeZlE9F2qxYX6
JT6Q3clUh4QlQFtKkbZBluaDuGBQxRDs2DxmOgfErzlyx3QNhH4hvilJcCbxwgKJSxA3edlwCjE8
Dxvcd+dXzf6yIrOT47ozbcf8y206iQGA3VikD8GNDcjdp2nLEtmHK/7LE/aC9ZxR5v3xNgdvtXzj
kIuGLpqXgK/lahNM47bjhwDC0Ok77Lso91lUqu1jSCBeUQrADXye6EGM+sMSz2cdXFQ7wMhXMxLC
9NQRG20rD9TeJmJnPMb7i3trvnj2eDjHbFYT1ZGc8FooxuK9IH1MXoFR5s1dPhbC7R5DJIY3xS2V
e/6BJ7OMJfICqZqxh5H7uvKmQO/ycoKZvl3lvxE7u3vZXR585E7mC+jTrHnGpoaFueRvMZluRNuV
oAQEFC0Azcr9lA/nu9XcehnmZgLRS8MCB1sg7LfugRnrDS4JdyjPaqCTX8ivmsvg6/ySYgJLr1fS
jdsGYk2khLCpAyerDGZlpOvvg2iqrgT8vL2clufCbN4LfdYFP9GbqigBHJDdMtemT5AiwBh/M1Q/
acB7m92dn8/2BZd690yqxe8SjyASW9ED+eAFIVFqJYG0eadj8gHQXQB+wmIsaOLnpOUHnB5/A7HQ
GfXVtemr2mECopI3sE/BgsAsfdhjttAVDrb+SjzJ+KRmzl/LfoXgr/G3N7BID/U6AkpuAsemPYqx
xCKB6O/jO9UbWeLfwJ7gkGqwD2S3ZZUE4JWLH8GYGE4L5Ts1E0qIIcxjIiW/t/IrYUitFh4sp+xI
RZnXDdn53pIMsXRzCCT9oY9NdbdZuMTO6UK3MMyUZBYoD0YGxAkDFm4BQKavZ+1fqh0ax5ezKzQ7
o60agUcsuJojw5jgCEUtkgNGar47Lpn47aGhuVxH6A1I4b/QIpibVjBX9vHlYzoUElSGN2EP8ejU
Ak1Ba+Dryir9YoeQLeAxma5DnKbe7q/9i7T48Rm32bBQOnMfmDC/W8O3fSmNVxR1OQFcaZumOs+5
vivJ9m5CrknOANWXxiLW9sLBodcAAfQHCNaFSWGlrKU2ZchJolOFs8JDa/WwZPx9v9QxbC0kqg45
Vq0BlZ/RLYOZeYJHGALzGu7dIH4YztOog9q5P7VmozC+nG5UNFMBQEk3LRHYMgKd5JUmP+jsYNSr
ak4BpfrDsMdXaLl9yUxhB2w18dk7f0b7kTG4ZuAX8uE7Dr6mMcxqtIyGLqB8ptj3iz1RojAWSC+D
R2Sd25NJlu6Vgno+UUZUOrA1zN6TMd25R+U3AZEhYReIsQPEGILn7BtxKa3nKw72sP41KigFdv3m
86mxhqedZRjvskt4MKZnqqoBQos31evwfKkB75/scplpOvB0TV8Sgp5izb6xKFz4lU4vhmR/wUJQ
Grz3U0sAs7JdVskwrggXOEgPAl2zjV+oHxwe69yigDv9oVM1Be7mN2Xws6X4pQnLCEwP0wJpFNvV
iSfCB467bYdpss7Hoj7VCgHg0esBuVcLmaX/RtLikEHTck2lyxym1p8XoPKRTWpAgk/tzOXsAkt6
Nh/FhdD+lOkHuKj78c4wwpe1+PweVwu0XR/q+t/TxC1rx9qFXIikjCteDZa4UMMqcASwa5EKMNNb
x6xqmZX3/hlf186bWXewhHQodJ/VvCJ98INwzhlYvu4k5yuxhFLluPVHnt9yRvlU2gOvQa37FYYe
iZ3AKSI0hM7ESUILtWxPgwamVk6D+Pinvieg7leKD5mL6qe/MDPWxrKkLkZsHuuefAAxTR61A3cx
PxPafrXscT0vq8mZJjtNutum6AEkleXRzEh5nZVwX8697aMvOyAh77UY3VQnrbMebfHn10uLOS/s
HrZLaLw04yAKT8TGR6tbR8iOQIqA7zZ4J88UuZRlKd+SY33UczdySlLlT3lKLzecHiS2wXO9Ma+N
1c/SuSFhmo3sW0tQMdPm7LRN2zZDsREYD5grPXUGwedgKyoVCtU7/Cjl5HAC6gAK1Zq+rr0jYh8+
/mDcWca8e8Yjl+HnnbKs1Hd3NA7YfpJCBZtt9WHfLxmqVfk7hHzAxzivkVDRrkPryd2CaJBb7CAi
gnTahC7sYPhC0LatFX/S5HDc+vyroD2gVL3+jy9URFAUWjwVV/Rm1aG5uIvPTyEn65v+rAWSGUg7
73uZ3GPhwW7XZH8KEZXVnlDuGJ3cqW2Hn0muSC08gXH2jSPeOuq1jsv5mrapp6M5T2P3Chx0Q9zp
FiKgGWvUCwa0xShKe3CWB1Yvvm7HcroWpAKyJphUQdX4RIP7WOXs0Gv5h63J4AmgLOn8VayG9UhJ
m2XnPhHlYTWV70Kl3qlAksE1+cE1WrpnBKt+X/cpBFL6sYZWRDIDmhzKPdc8LEFBPzebsbTK13En
w8a8VGNJvG/6QofRG6UREqhxn4xwL9b1wE9k/cgXh9irAraFLCdkwzesFkCUgBqL8GlOTsbENhmN
lQGZM0yLvcCR/OmKz/JUUcDl4fpwI67dlVq1GAyIQMRGcZGzP5HyXNtmeWXMhRIq0axd1gO6ivog
rbSSj9rzPAJ3p8xaM+tPZY+492uAc3t4RFGbOvylvB3kHmIcY/L655uoifVL4N0/bXBavuQevojh
4FRw5CBnwDdvijxYbasf2H/BQ9tTj8ndN9cCk/2yFqzb4II7RR5zIbP/EHXDit70BTlsZYmnhVrm
BDnp0TWX5Umw4uK++JyBaAoX2zICk+5qacXg0EK1PPmuVISngZvBOjj/k+p2azzw7APfB1q1L39k
GiSuQjCWI4jgDnl7V6078fmegb8Hg5lIrLWr8VCZEQLUY2JgWVKrrdSO2L8gEI/eRT4QAuzqBGpm
PonhCRc4zgRkh8aJxJ7vENvs3iBIGiMh9MvDSWHw+tPU6LTvL1DOT2y3MumIEieByKzrUiJdPwuR
2e2pUxAnAXcM8TGHBDYtHQM0dUqK8K4V/WKMUPkBObnANJdkci63XDRW0bsK4a7a+fsC62pHEiNM
MStafauRm5R4CarD9afl/9oQDLnO+HrCZKK2EMYqQ88k4hhMrk6+sR9ly6GWuRolQ6h4oE3zgLGH
LXVGvNvKBUPXVTw9qmq5CzqGCIcdBuczV3L/cj3lUJlX1I1A2lKrsTFx6BchcwyNR8i9C+lFyLe4
7hFW9io7LPGkBQghBLk4d427PFAbm1Vjtgra5ic9hhpe10rgiQ9RH7xouJhxC6flKuDWHMA4zh1E
Ec4uGn3xHHPr72gL33QA//1mluJsjpl3FXRIwRCCmRjMN9F3qCsW6YvhG3MuZhWbk2rJYR5McvFx
rlU943rcIHPxux4m8kZkxDTOxmaSP6CRLxflxQ+mmkWLdhqLGSnYvJbAR7Zzc7hU34pmiMLFm/xk
gqY7zlZpE9KA0NFUHHcNqbwCXCs7r3d/cf3T/kpkhiVe0f3zgOnjNyBHy+dN0CsTUCYVlZCF5yDJ
cGw2KDjcfFGl665THhAQfnZyqZEFWW8UFSkRF5xDPlzie8TBonPFVWBXUAn2yC6wazmM+N9HGLtb
Sa+RBcbE9PbJf3lokmc/TQJJaMeX6wJWqJT8DWG7+JcXzk6uOLrPwFbnqPwxo7Sgs6znMKCIP725
2Mglm4yJUjXuHgZmmxBM5NhwHbsmTskrYn3PyfzwjS4QkYWvVlD4InuWLm33saiA1RLON0Yw/D1Z
qc/xgwXF8jzVAlrfsPzYMaYJo6P+lfn1kBLrepv8eDLMzWG1P6n6++NYlazJZP8M1n8eUE1gsIP0
TCh+OqWoGLl9v7JED1dssZHQoO69uBSPCpf9RW7yyH+qDVHMa5tst0ZMVAu36Xysxf8Yv+tZ7g2N
H91NogTM2T+yFPUAjVCCLeXwQJXFiBfWt9pZtbQ9OHZ0qBFovGwC9da0zZmqdWdqv03azR5R0QWL
AGkIF6bk54eAi/AtkusvYnbqT+PoOSZ+7j2suMv8y+Q2vnxJnPuRDlgZByoxsxbqKMIYIe6rWpVc
VF/jNjMDEv+DSAsOrcIqax9SnrgA3hZ/MQpn3kVX5HZ7Z0WEbE0yWNXmcW1z9Se8OlRqQ4AnGzoJ
jPN1ZtOS8dpeqSvXtm8oQVwPlOHeDSWV7uTeBYbYw4UllW1E7H38w9qhIDRNbeVbuR+O8otkrdTB
ZPnwsPJNvFRhmx7KYX/3pTbBfCqI2ScLgCN060+dzo77b0BwO3WtHg+OR8BhKZkqOiDdeFlsZkhy
cbcMSiUKUu+J4csn6HGjcYp1vuopJSVniEsh4G91uKzMju3PftrGwOaWx3gvwK4K0IO+AnVEVSfu
WpQ9i+tISC9X5EA7HOLEHEr4PmqnabowssQWfo0rFA0lgF8XIFXCr4DQcdI4aKqo3fn1FjAeARa8
1gA7diUDkXAlZPsKci5KsXmwPfuiLviuQCptoDZdUvvInScJHWqUpkMR2kmK8AgRULQYuZd7ydiw
sX2sCgQTAsMpDRwJNgdJkr6g5TZMW5+Nr0B9U777DyGVXfwzIJCRdBvqSsUSxxv8i05rw5gDWguK
CuxbDAaTQMLgKFdnkZZAE9DL6PXTvH72oAXICZNd15bE1OS98gcZE6nAkPHgtBMiN4OCRU0COSdu
gPSM7qApbKUvW+rP4+8hYdIBf3rCZvJx7fzW9CgIpRf9grkuzUkT0KFG9ignu3tpT/p+vYMoR1fF
hAoFJGbQhX+kVyrbfXcsOAbjCWF5VxCuBZfy43G/0uOZr83yW5xWojuaalQtow+T8WIXPc0aW6Ij
UI7Oo8u4auorrM4KPvml2S70cLY8TPROoCgsXKRjS4PgBnmKhzy3sP55lAg7JhJHSS1FHP07dUp0
x2cG1d5U4IJg9F8P4rJUqWX8ph8+yebEfBb2KZnHuN6w5/gMoQiPcRxSPND9TcjIRKMGIMTyPeZo
OTnAmb+RVlOAsuNfVohZwEcpfKL9od0OXjVIrVr7QsIC/vr34OSSws8j0KtuRDzXeKL26lVbS1do
TQQoQWi7qIeex2zhpP3dU6udzu1wYNi+zVmdjsrTIDLa3Zw4bbv/tfbCo9EHeEQ5bqJPTWZRXpx4
UiSJclHIeTpXxM2QKwl3bbACArT1x00HOy2GiqrNNKHCkcZolGpjMOWxMl2/istfkma0bRWjb9Rt
+Lfh/ls8+pUJ4dgeWae/DSTthHFjMfsxBP8k4m1M/bs86mxkiNNB8Kv7z5VrwaeD66+evlR1kCiu
53/h2PxT4K0hqCs3cFvGTL8pj2k3wNdNMBtohFyt9IsunL0dP018KT5aHTFBjeStZAstElKVVj3E
mbEXL3lbVcos37JTKHVQ3SSYM/Pp3Ldxuo2XncQlL22YvR1Spy0wf+tBv1LXnbQyykxzp6x9Scrt
QF8raanlXPkhZhGRheQZNIpQvIZeNWyhu8MZkC3WuG4Zc/kwgKd9ay7CsxjEqD9QzIU2gVZX90vd
vc5ejo1VoAPeFEPQev4NtJcWIUMzBEm2z9IfhEM5ifNPkt/CWn8kp3r8St8Len+Infjl9yaI/3iD
APmDhGsiYm3Ezh1MqileKf2bRbh6/F9LNd9ogS5aXgSpBBC44mznvAB+l0tAEbk0e3EO7sQSrV4Z
FBMe5ZzO30FDd8kYRJdlsaMuheDDb8BcQVbs7CbP3r1O47WzmyPJUDFWAmE4CUkodOjTIiABRAMC
cBH2utBN96W4p4BXOfmtr/6CfsH7dW7YeqmXXJi8t3l4oOpZjt6DxYCdG2LL4hLynZxOTnYzFi8B
lymYtHPCSKBB4y+mWkdgfUlCttdyfsf4vyIjtcmpOVapnFlHpfxdz657G+ruXzOP1JnQpwxJ6yK/
Sc48topK/PRlMJsCVjobBQ/5H5oicqkZWlwirQr32A+lrvOPATn3WRVnuDEhorrvoofIuH9jyemz
SQW/f7J/mIKMiuGgIIYLckSgHx5qO263jIu+YpXxyG98bMxn5w5gbZHowI+VhWPK8OZPlRH6Lyx7
W2A74ksbi9adrXOJ452QbL0UAjjdQ7qdY6/DUXdIARwCQnBDHE6tjuUAhN90UPamsZaatID67Li3
9AzSfdy6Jw/5gu0tt40yxyPnGvCXVdKtrCNqUsnhGvtjWhfBELwuf+WJhPp5/943ElBGKjxIsoT6
E9gKKYJ2ZyjhG23flU6H9coBg7wytBxYVLIsT1ISRfl7G69BhG6OAZDSLN4ikXUqJE5zsS5DgjmG
f7ja1APyc5zqBeKrqOPhRPyBAdW02i4O6w8dyxB5BKNUKb/zIYEDTX1e4qWtsPWB9cSufgmh3f5K
5p+EAO3nk6mZ+YiDtcjy3P9fGVpbInFLnOuTp49XCaRyuzUNEqp7UrdJzYMavB0WIfGDEw3W0cAN
lZRJJo23CdIn69dGrA/DluAmAGCLqLh/9zpfm9TKk/8uSiI62785ap3dNCgSSGbHDjF7BwuRc9Go
rO7NPZ5gxjlA9dHEw9Onkj07affmNPLD/f24I2KpiSClImRVSMcK4VSouVNmGWB7CCx8okPK/mNq
j1Ssm1sCC0sxGnSnttv2sFlklNMyqhD2Xpb6ZkTCLDoL+L3Jzr5c/Au082uZ0U2FcWgV4JSphHku
lNtvXq6ErGWRISxJjfXbQofBDYxZX3aT7SwFrRKeTeKNRipjj1YwaMKXFOQIB57SbBbIU7tvJhBg
h9p7TiG5EX7CZY5DhJDmBn+aOPakfAHbmGA1Oru8cLTkFLm/89XsXDiWe8x8lv0aZevm0Py/ObmZ
wmBUXLqhJx0zmAdwk1Lh7bLW6XFESJkTdz+78SNMHLZIZ+dteB/oMkonBSN5voTUSAcjvxQ2N3MY
o+jDxt4TJnf8uc8dhtRFBoggqk60XbV8MiFP6juw9SmYbgDNDuzljbD/iPdBdBWNhq3Y0rNZ0MVy
mETpWS9F7QiTEfQyaqXO/vAjdQYDZO5aTdZdaYlkukTUXl0eqRFoyKzU4Esu1IgbeSj405nXCtRn
tqIpHvnvC54BWGCVkQzE/feHw5hnardakzdcUSOf1qOPcbR6Fwciys9RyTGviOrRoeyBJkUEqK8h
pd8dwijdU5GtjHrkbA/hmdYQdVfHYVtGavahfXJ+oX2lSv4V4Z58HimcW2/68xMF7lmn2Hxn74Ja
hoJJFoHQByszq4Wjih8wGXRgOymPcOTdL/93gQoaDZZ5qq5rZubhO5jsjwp0eRDMPjBBRNBaL/Ie
mQTvSHhiFVD/9kOMcYlZU3+hbXFpYU/4+y0QYmp3dv+3BeFgAgN0LIS+rBJAXfp3nF4SQcmivNBM
m24jO2GFkSR6sPn06K8I8h15a70pMo0vNGrJDZNz/nfLs3ZXw0WiFnzyYE6gY6HKRjvGwhMopy41
89F3H1SFI9tLl1YfFpcMDyvDjxz4a2vvkYB3wq6SRp56t10x1It1aWcJL+E4dNYj4jxOa9qLq4bh
kxetTsaWwAyuhL5p53T5RQZFZdnTFIAC9ldzB/QjpcmuuOreLncHF4FcBTgKjqtPinr5sEhVE0e8
1LKe5xKS4H7xq1gPXikO1b+1QauCDgnIz+EfmKxdDS/jNq+7VG/zF30D4Cto1yddauS36HvZ/0aJ
rL2SK9zVRMagVKa0I+E6XyCYbKqrZ3RGhzKuTRMyu0Y7IfNkHUAltZGYRTaMvRDL1IT8m6iI7c80
uneloUjqrTmx8D1DIdc+IY7qn+esWtdYMRtMCAQPjqS2aQJ86ACKl3DzM580iQrrdairvb4rmycU
d41yLwZTApNGQ1Y7wDIJDnhP8QjKzyHrfdtzffl3Eu2J8LPGg1mXO9gkctxURU/4OXz1RpwCuwcS
TQNHPIgrt3Ke4h0WMIotyepvcH6J+uCH2hNOdNol4tt7glGWR+lo86klvsqQZu/ZqFyI3xk1xOaV
/CHkd6vLDhAg1839054lZBtBwdxUwESxcg8vmPl8noNRT7DBIkE2GauS/mkQqE4NPfEZiHcepjjP
CJdHl2vSxiapgotYEyFBJ3MX+BwOfJStfimqOukUyQpCdpFiGI+q0SkGeHIRFv2jxYHetWQabe/p
9j4nO3p7+gm5bxNAsjtGhpwH6BT7RGPePARzTVRVJi7MLlGPJE984PG0VGTWV2gN1eUELWv5tzIC
dBDWMkm3qNMQCZlo8WsGoNPU6Q1iE+5obTAJprcoWXfH2WfbHrrBvDtD1RKOOTdaT0/XNJKnwZEz
tGGNKDRp8ABrmQ5e35bJYtcLyU2xCQMlHaGmobo79rb8lxbX5qCtRehEcipJxXY1oukDgyzGomDX
6Ipid0QMiDWNFMUBHKLtCNoe1fqw5gnMzeYtUI02ywoiQvq9//M4+5VlKRwqOfC+PAIEZVpZDEIv
kMZ/hnNpIIJq2XKHkednaOr11pz/r40dAqIsiG94HP5ovMrRqe6uOsDv1pKRLsQbvg8pkU8beahZ
6Vi8kFa7WNL44SU3yXjWwgyWDFX4XYCdvjalMVujHL5Kzno3aJm3yAML22vWa5d0rUxk9Chc9lAg
9ey4DbTM3Vacr2ODGkPrk3VLbwoYUh5/UdRF2jJSBKFJCjclU9dxlEH+vw1jydjOd2LJzcYEU0QW
kIAdVMy69XLhgv1KpSMGv/nuM3wc7UbYiaTolx7Nev9zFQSLKbDePn0cSYO+a8G90dAxUKRyGhzp
iBL3zFktzhNN/wZ0dsSPZDQVrSn/BhAWxWuZu7oSSZCeL313Z5lPMDmLUaQsz++XFdbbfPERHP2l
WwU7Iv+9IAFevbyKtXi1DMIsspWs6eGkFrWhlfba9FZ6WdqjxdRuW7RTtOXA1kU1r56uEXG9Pw7J
/XnHwAAep5ErQkiESQzDTJDYrAioZ32YohnIIO51DqoZH5qgAdQ57GOMDrj3axGic5deEialVKVX
Yt9yle/q9/7AuzHkJpRyIaMnLFLkQPl3/2JwO5/9wJiwuiF6ebeGc+KjtFsXc/DHRi4u5DlDRZf8
kqG/5oo0k8hjcLEuouADOk889bQRrlU+KJtLfi7GpSJW6Tx0HFcBb5G1IEcxxBbZ13FwrZoNjVgE
pAh+XgsEQEEpzasKOnytyPU35AIL7hY3hgqdsIN3uG+A6dvtX0wBUd58xscZMcd6Q2simKFR5V3A
n1GYx1OFLyA1kPUxunCIyPWPU6AVWyIkHhc4KQJycISqvHKhagWlfWap6BWLqknbgnnkP/649Ry7
b1Tqv+OayG+iIkJTIFTAJ6xGz5vNaffVtLTei5VsxXfkp4QPKpUJHIXujRpcvb5RbW1RMMfqpK1U
rjDcLsX6DSQdfVQ38VHzTEzXwdE45wQvu/A0L8mj9V7xTvmAWiGy9lYBPphhyV+ZABegKXjNtKao
sKde2FfP0QiFL5+A985AWppvG8wYN6/iZv7I9Zw4DSeVszlghDHk8Nu4Hqz62gRbET9eZXkfBKqu
99wuL/DFI61T54q3vR/4TWwxLfBf1I3HhBLnJnKU0ChnUMFxU2NhTlDOaLdOnRhKJzu/yztVI3NJ
SLQkNSiNxsDhCA8hxZry87Gv+noiVcWcw4tt796SCsAmYo0G+W1dSF6xpkba+Y572yIjO+FC+2R2
sIiQfuMy7FtuV92TbIRighgDBlPF5bk3wG2+4tFyPergekBJQYplWfkV8p9CvR4mhIdD8ZMG88dd
K70F64GiG7nf6syOhLGMevT4T9234kbwxCMwP4J0Jd1KRrkATuxlwP+nLWF9CLwP7J/CZCDqL+Gy
q9IoF9fK/xRdJq0xAj5yTd8jlzh8c/0GHqK6U4AMkYBrawNdB2qxBUcjw/aGW81eKE21CJ8Wyf80
2X+lPcdcW00l47MjhF1dU/saLwUWnXCqACen/1DR0jJkBUIa4fuaWIkT2YQJ5pIx40rB7uexS/ao
Bai0tvWARehVGTo0Otuwz7eFW/Qi0EnPbI2kuECLFx8AjH0wP3TYRd1OTt5DTnWRwoFWsRSNEcx8
WKr5tX4clY8J7bpQ/ALnvaxvpbhcbXIqavVUj2w//Dn1+MWWPjSNqG4D0gtsFlFz9isY/9YntyNE
VX0BuBjQ7C6+EIiOQFBe/fMUzse0Aff8FP57WjNhQYUpO380/Ok2EQuD9nMPjW7Pb6vSxAKkp8ee
SBJOWLloQcblE3ZYRMXAif4I1v6X5dIo+Xk+sfaF7rOrDFt842SbfT6dUiTZcroQZ/95+WBXwJOE
gTWXa7c3RHK+cNoFcFD6CSnBezj2looQ+Uw5lq3yFqAbmbAaoEXod0gQlFpPMwHmPqUyPc/c9MwB
F/M0J/wME8mWEyjt5v799cmIvp2sYRdwPYIedqOTFPD3B4JubHMsfo5/0L+FOb5eklhemOeeU5bR
wbvJ5fieujn7hJWnjpbdvamfDYWjfdEkHSCK/6V0CjglM3Gekv01NIWSWrCPTLq/hZyOYrLixfIt
2I3sFgwuBZBeRyGlffP4vnBNNX84NKXMXh+e1qpKhgvXVej0WV7e3CDk53z4pYEnmxYVlSzrFZ/i
svhR+ZqmIQw8FJOo4kZ1+3FspfDEfeRDNXuXDz5ykMRBRHLaS7hIHHY2HMY80ICm+EcLdfXJZc5z
4lDME4fJlI+Sk659k2gHoT66Gn87Bu27UJgRx1+EmIh0ssXMQkVjRDWv9dCFYfHL6Pjwj3U5l3j9
CGMCrq1vQtdfRl1zYe26q6HmHzPwJerHwaw0TAXf0MwLLp5S/hRhpzuItl4aDVKMm2j31L1Gh2+p
uU0ZNtzZZRdoDRja/pbJvaviicG6IlBmr892MM3kELqbjpD/P1UoXparzHPjDn6mU93pWcSAitD9
rt3DQ8Y4NrUe0ebDxESFDc04alSShhS+TWDVDQCil6gY8eRu2HohZ2cxcpZjU5FqSVOYXi9bgRUD
l2kmxbWNnqmT0cbDmbA5nZKg3wzduAlSni3TMjpX9/lda04o72gtzvpmP2vVMP2UFZJxlwKNvxX9
bGeamY0FqGRE4sQ3L/kGkccLkA9PKsj6xi7VO+PckUVvRkoUYR31C5d8cNMlY4SU7YW0cMDrOiNB
aR6SPDEiSwvUwZ19dKN3pHhRJhzHsEQVvJTMHHORkMjMsp43fGNeh1SeKMu97KKhNf/BNACGGvL9
icikHKkpQn1DkqjbRrGKYM9N3W9kGejcqHkUEvDCVaSsN+gxBFdzaTCA11S7dzaYt+F/nWDlYTzz
DH2RRiyNrUttXq1OeHGnEzwmmd2p2f6HmJKPpFOIArmFl5Q2klelF1Xd89SzCI+gtq/gyu7k7XJH
BeT/m5eZIU3HNvkEzoNxN9wA9eqeJmeJ2F0pn+UIQllI98L+mnkjX7gf80OrHEq7o2QQNd/5eohn
7kog5rXEiYrmX9WL6l4LjymksBrf0PXKGsZR3IdUue2OI2wMKiiICikbCEIBS+Dfsms2xzL+LuXn
LtwfkGzr0NdCcgVnGds/G2Nn87TolCFKtykfY8qgjEQeWVbh8iZFaLp3aZtcI/VHuKJ32MIRuUOi
Ydb+0PNbeYy8tzCwtVC5yoyB+LBx4yUEJKFlbvBJ/sVTCzMYcE7Dk61iQShRsrhXm7c1DqYin89o
iGMJVP/byHX7d0GIW+puKajFymJGsUO/dQ3jUr28DHsv9yRtZ2wLK/cHuhBIHtd4CvYZGcYLNukk
GhR91Yr/Kt8WyiOeMo4CXYys0yEowQ/qulJl0sFvMq7wbTTwwSXyFWXzwPBu5tbuTauUzQqFMJX1
Eq5828IC3Sz5yoRJs5rJTW75MagkaIvdIu5D0gqtf7RQpFRBD9ybVgJ0Jpz5Y8LCUuYR9nrzCSYv
f4rIkiG4TIYj6M9S8Zr9RtyjEeefiY36o0+iB4N6E9MHFvCgW0C6EjckXVwagz9SxraSqiSyy7p0
O3lmLvfI8MqfNyi+4QIa4lh5ItguK7ryIfTG7d8Z0fj7jzDb3ayKizQfBa1FqnUqV38lTFhzxjse
Bw8pTPQiPdhfeMZakAY0fmv7KHcmgx7gB7GOQCzkohlCsJkABl3q+vCm6dFR6WL3dkkiZcwKTNd8
T4zjNTnIX2gaSVWCyaKjt2kkK55LsupEbflP6284MV7yggUP6wL/BE50tBaCcHEPj5OmJnieS+gs
z0Tq4MeneKXTc76FHZctw5EbYLC6x/rtfElfiYmQuLf1NitnBehts8KlV2Sb/C/wfCXeQacOOFjV
Pc6k4T+gSD0qDa0FGGS+1IpY6PF5NIJ6lGY41o8hFcg26fWiT0eXWDNOx51LspI+/uDpr70Tmta+
vJd2bmGNW3qVYcE8ihP0FYrv+sMECSuy64KwizMtqItaRsIHkrnqM+Yf4atsY5NHTyExff8C+Uh4
yCivc7xDzsyyWugxv4s79yoRtoDgGrPTDjWOT2Av27EYQftrR1MfgB4jG+OFPuUpTDD4YOVlaYM3
rWpvjevOIs+K8004YL70A7XExbZtnHPRbD9XtkDQXx1SLVte/snQbfkYjR3Gz7rMMlWySUQYDdfn
UmRdffz8Gvo23Rac3PQgJyZtJSv/8d8OcbRsNiar5R7Fhl+eDuPPVkF82nSw4gsmOjqtFIXTkbSf
aYwELq41Uz4RjboLHbqFZS5fbsHpIkydSO6m5F+hYcYdgkE893ReSkO93/0uLJMpc647EXljbnKe
PYxRDc1Uc8I+humycg5LxXmKh4NDNe9pVLX8kz+zYwd6RkSk8wR86VgKH+sFsN4c7w2GLWRuFqUd
VEnMe+OdiKYpo9VBKa2URHgmUu7LL04OuAUeFG3Ahk27mz3FfadmqVRYjKDYJm7GC5hsIaenoAED
Vx8uuN7jaA+fnNRV7wnYCrmPB/Fd9CLaHUWm52y4y3HsR6DdSu2uNHa1WW5ttDqjRkc4aui7JeoI
WwRb9ZVMx3iHJfDNzhzbNt0VSZhO0mBYiQptEMCZh2cjlGuKa3jyrRUZTaIGiIP1LNXVDkuYstjr
5LR/i4RsZOciBrjBFpLuuwW8EVw8lREFEWLFjVmwkizcI2LELkxabfPG1K13q+v0AjLa3rDY/ppG
xlVNbsz7pPlugAkvbIvDstKzaOlNvYo7X3E3yOTUGEMCYRZg1iH011pBL2t//95/ycRQ+Tima2Q0
yVm5jMk0bj8xT05f9suhwSin1XhBRXJJLZyezL1FjfWvU+oOnahbt3xF6Va/hUcKZpBgvXJi4+S+
3O0MSIfyERS9ZyaSKngJfPRvKNaBdlPLJzppyAStdOyQAZfVLjjb0PakkFc/zdsQHvs++5l77hgS
Ahto4Ykn3cxpf9eJf6opSg9qkKv7DPXX8mPycb4gdObf+85UGPQ5aPcSKZ+FD/yap/5g0CU4DrFy
CwK8FaLsiNh3qjR5HpSHNJfRCzJpdFXkY0BW02Se5VtSe81NQ4ZjJ5dlojmp9GgEHKFOd4Rqngsl
qeYV9arUU4WnJA9tfx7sVMn+8dadkQZqkDn9icVhLHmKxyuNlRay+jJlmedHCbKcsgu3EL7laVuc
AJvhbDr0TdOoxyVC/Zra8tbP84cytZy8ygvOYwIgtarXhDT+tjhCNBmbpQ3Y70nLEod/36bUrw2Z
vkY1TQsMd27ZW6+OwUohcPvs/BL7z5ZMOFtIfO4ELDqdDqWr6RuVF0XKDmF5zzE3qEs5r0UEoutm
FpnlzUlFtvR05AMyRX1lmegnV/NIAebw/pf4IgWYnJj82eAb4taO8QtxBIRZ6HBKt7dhP4z4fXWp
qKNkr7otyOij9nrm33JwEP3ATqnKnGBEN9bZw+1vROztzo8+IJwPBrT8XDChcnZRbwXAWLiIwcJK
wiKciSDzgkwThUZQM7zudfIQ1aQKt9boN0KHB4fPMQXeXxqiPRKz5Dk4XV1kvIIiCeOdjbc1nU7G
4AAN+c79i4KgD2JZTYSsrgJQ/Jh8JjO7os+OsrgPXartqQGQtLldw+pBgdHfKrA37wGE5PC7b7BU
Fv6KvmEiSBVJ9bPBgPVDrgV222NebG+8c+YPo4KByWI6J8jQIhsJ9bjYk5Ju5Ba670VQOcSE3/EF
hmFnUuZG8roNgn/3cx0xNeU2pxch+OyWBolCdTMcsVX50hrcVWK/GFz1V+p8u8g9GEjmrYp0WoWF
+4lBAv13K0YPomoXzbQSngh6y6JvDwSbRTLBY+rBJUGLGa1tCCurz+q46NqhvJ4RnT6ewYnmATdd
yOiyGW3iA/tM5oQh+aBfEwXa3ApZrXoJ7N6nzNhFNjgfF6VUd7nPO2bD6L5YjjujeQCBKHPWXfIu
bmygKjFXPSm11fNfTeBKmL2CXeFlIbKnNsj9b/F7aFYtdzjypjmSpteAX3xOuCynqxn2IxAVVW23
6er9SH7cXSJ2sH2gsDfLAxPp9kJvgxSXY0MbcwKI86WifmvvCUy0eyztEka2JPbId58AtZ4Z15Yu
ZgRB8XVjFT4Vy05ZSlNWduYalqHi20ysLJ3uop7vFW1mv02kY5xmL3rOZbD3iGX2BEDmgYmVlTQj
t6QgEwbPNBJ4W1piiMYymkr90PWVsrWcFfivhwc7yRMc3T7uRf6RpRhc3Ig07b1Hdu7AG6UClus0
tCSUijLtuiPeMw+sbHQ/9UZ1Ps34XiX1u+MCbJej+iT129NWtHFIcHFYTFxUWdHWycdSl1n6Cr2k
dTWx1RJNM/3Uk6Rq7wEzqff2ORjwGepCNk1ZxXvjU5uF91u84i6KDos+IlgdzErwn87I4pDlnO6F
TbptXzAXlJJrkwvwzeq1dgzJJYq//BnK3GG3NGtM2OizM2j4EuNQ6+LIE+Bv3sWxlF5w0xeL/y+H
gz62ImZxiCTWPGdtIq0ypXSwgCU3s13B7nXxbV0H5oyGTuo/yBesiK6ol2HiU59Gkm5dpdID6vCk
rC50t7f5ydPx7R2fO71W8qKd6miBgiGr30vsQLZkR2d3TqCXm1JdGblSIqMTA+BunJvgsFZqU625
hR+9uKCLwQZpvyfI3FfS5WtZECl8wAHCyGkqyVOCkotA5RHlR7yJnDTA8MMM6y3MAh7dGcfgk4Bl
SZJlpBDo8V/l9VMiwvCYVvjewJrPqXNfB8R+FSq5L19cYRUwUoNPdNXbGOzApUYqIaYcN+JqQwOI
SLFNc5NJunwFwHBIqJqglxoqZdMGHdNw533jT99O5Xoq491QDNlyfABNQdbwh9avbTmcgrcmTODl
b7fGG2zIt/q3p6PYDEpMz05SkDuzjb6cQ9o945CL6yLT2QdkL74hER0aH8DFY+CKOwEtZL+xmmlQ
U7WErKYsUh2A2m7t30q31hP70a9KtEAGIv2Wn5fPRdErbtKEtx2tZnR9wQ3TWMuQCdnQId+J58bE
7whG5EW8fUXlewh7Y5SRU+nPcQWM8zDdV0g0pOo4k558f+Ns6xEylsL13i+8jdJj77nmO+d5tyRK
tlo6RUhdv3/sqg+MzgFg1o6DT/e+iLU2UHMMbTdbi5I2im2EiKheRMXu0hvWwY9CaWN++r5jaLUb
5SIPIV6zLEfLGfuIT39BHu2zCQAZxBaJSf5lfoPc4jwWK9dD7hdTFBCLjBPEWJNUYy4ecq6OTPbW
BIrxA7raSU+oZXQBE2VakwJzyxdzW4G+lnJMyHm14AzCJ7RWcYtF58Z1nMU8zwgAS47Xuc+EzeDi
UPzd909ruApu7bOkiVUPJV6r8GlOA+mfZHbJPg8ubTrp7+1ukdjM9UeiqeVouC/5Mg9NJvYW59Oe
ENpYBMKDIwmnoaSwTeMkSYu6AnpSOF27fL7oEFSj+3ni4wFDpvGYo3jwJYZ1LftNqKGoZVvQVoq0
qG4S2cL7ToJ+i5PquCsiPa2punz2vb7EYcc4v28q+syegRUVjAOiP+qHmZ2EmWoCLT6pva/LMvMV
lfUhAnoH+XY7QzA3nIfuC1sq9Nv2yNsExmy78f0LtRrBYWiBm3piD/x8Sqf5QZqBDzUD7Eic9xj7
lfiyS+JV5Os7JQ0EtzYKn4MzLCqLG5XzQCf8dNPtc3NzJY2iGCwkyDn1spQ3ZN1hmL/jrymfgqKv
RCCTiqthl9FEjAfXQ+6toO4xAfMUMqgQDby8Kbk86NPOn8PZZb+GhE/ZbuKdClILpM7hyO8UPATX
RiQ74RvybKzvQiyYKfPu5dpx0LfWU7vXjRpDc1bE0pIbwULH3edN5MvxQ4t5FMTgiSrqA6P3JV0Y
ZjquOpO8NoEk3W8n5BVIQM4hZQSP+CW4S52BsMOMZaFI7dHTe2xMHIXddMiUOTIOgcB2jF6krT24
8XCTsRoBOwN9dO3u0APM1hUT+YQfUv0PbEm+gnfSZAvm9/8Ox6iyG392YQXPQ6sDA0S6u2GhK2mi
z4fDDEUc4MNeq5Z3Fb78nfB4SVMLDhby2kuPg68mLYM/kRXsbKZJjL6k62+J4vCTR/3O9n79gK5d
abmVKBzpaTpCzLAAu1s39kQdrr+A8Qc8/KZvKrSkJivsjUZpp0Z73mn8RtTj/oP+Gp0wtVGC2ABE
C0x3G9eN7p5x2zG7qMQWEO6nQfzRaJiGgmyhKU6RWEDI/PEMKs9AgP2om7+DE3/vJ/IF2/0c9bfY
Spi49eoNjiV6x/DieRgDgU0pzQFWVdZpXuIG7v3kw49U8dNT3vAfMhILsL3MT7i3Qp/Mo9SUACAS
9cV8jGgYq4YjWQUvZylLoWqCpGp9CZLL2YQSxHICrICYLWgG4ISlWBJxxQlSgA237D6C9JO7/xyp
S3Nwb4bD1hrB+paHUu5ew/MBjhVe3yVgt+cm3RcWKtkr1vG/Oq1Zxu/oSWa+risb9+oozPzI2RXQ
7Kn9OywnE1UTLnz7m6d43lhKa9VqGw39tlt7AA6zkaRGxqjOj7D7v+DpkghenQi/YZypRC+xWYom
wZermUK+neJcFy91t6XnclW8G5EuVtqShSdJYs6uDuE+6GKLjjz+t0XrHJ9LOhXZmQNMvyx+tx/g
f3WsuTt8pvkoqU3PcSfOL/EQx9lYn3kpWNcw13TEvSoRsAQyRxX4roeqXbONVCQ8v3dBzewNG12B
aONn3BK3kVeZdBkpSKi4mi8MJV4yqp6OyNLS3xqeTJ3boQSRMeOipJnixPOvQhM1qkhxl3Px0/lY
DogYprfQYF1dRlt0rMABYY5ZEW9CYqrN8GlL/lrUkSKiWHFXu7wwimtGTwXWOIXrE+wZOJKhIB/b
5g1TCfdi6LOkiXHYdMk2IVmJS4oEgDSa7+tsCqiHQECc9iuffeP0aQgMraJZ0ohZYMcd61m8p0Ol
LDfg3OB/TgXffZ/tcCH+hOcdpi5o49+LpMNNsQiivqySCFb707//U7dCLQdnI1yHgdOP37PDTq4e
I1wj40xzAPkq8vHWXxELA8yfRkdrBogAYZcYrtfVzqoAgXcBUPX8EXXk6b0wUgCCtgurVHGHKHAO
mm/JOdzFIlOua6YBWKBCph19RHg4Ho3xCfw4PSy69LE43RQUlsPoUwTcu1U2gKyoJ2qU4IDrFswj
4vYBzN0xypm9Dn5iXtptWbcCwCANrrs4veqWMV/zlN1B2DGVz//SNd74e/HO8aNHcSWPT7dF3EUU
AUj9Hlf6RcFeEjXH2ExVeiDQs5tacu6GlO1VA4sZsD4CmdKEMAXlGMak0l719YNjmZe1P7WPTRqZ
icG40bdivPm+UdikNMU1DPmY/jmlGqP5kDW3igaO4FN+E7pyo5bG4iwlf3zexZXjWYvkB7T5+xD6
Oqr9F3Znnr7uo7vraoMVnkkN7aXVQc4qOps536z2UAwW0jIW9zdraBXs/GcR0pBUJ3DoV5wSsOB+
w3YnByFZYnqW2AV/zbVOSs+CaaAh+m2aI32G/1yrem8U6BY/USHCXYnEvuH+rAg5Qtox9GNLXe4H
ey2rxsRywsVfnKwFkN8SL4oaaCxlIvB7v2JJPzMxR+aMrsg5N3fqnj98k9Pr+l8WqJdGZlmsMnIl
eMtFku3jcplMVtuOyFwmZhs2LqWqI6y92bnp7LYjv+BWbIGmbcCAJTk5W8y7u2sz4oJaqiV/8v50
dec733SG3tZ6h85Z2/Jj1cyrYqi3ah5LCRK746qw20rswILswUkL8rvwN0m8h3XUEGo7wkcFyZtK
8lXoqaVeZzi1laj7Rbx089n6xL8CwXVxOy/VzkWlC0Y3MLhsskIY12wlqrUUjzYI5QtLSGK4g2PG
qG2kPVvxx/e9nK1DZXTZXMaZOkqBVixzg+ZvfhkLlwJYD/XulIGOXIUqXqxEWkXkvJopKazKgEi4
88lvc4DhH68YKE2MQ3Y8Rkn53nCY/dHfXGEFGnVQ9U+8ozo9PtIgJpnbkMhZhtN8Pucbr2EOm9YJ
z8yOHsUruxo3PWLMKe3CXm/htEkiNXvaz11XkNjVBdTGWLLveV358IUWmKbX8NVQ+u5mhnTTf03n
8p8UwSUWGxGzsiRggJbuQKmk+KRVD+H7dfhisS3snmhfThaI+49+q1aCXtcX0htt6jLXSfPzrIiB
S/bSWPF3XAsYuKQ89+HtPRkAzKScVIJjrraBQzR/wQZSh69F5/Q/KQC0K6ylqFVpUCwnDlLjK9rQ
ifB/zNILTEE809MhtW3HiEa9qQpE2h3zgIqlQQ5vxthIolG3R7bMdPZHkPymfybAFeT+jeHm/Dob
x9Vb6NqQRe5dtKwJHwwmz2TLM1elgTC2lutsE2Cqj8WiB81zBPEa+WTodl+wyYC04+mWQkQBAWGR
CvID3nx0/4tSvhRj2q4Rq6F1IdExDP6C7FL8KRZyYRyUmLepAL8ZVOvH4NJftRcJNDKwO2Mp9JlE
trbF3dfM/+QTBh4pUxnGppl2wsvmFCNHwRlkxJEgqQMWFZvRS3As1KJryVlu7JJ4/pSvgUnWlXQQ
lVGTrPzRn19IZr6ZOtx+2y4PJesieWPzwXhzlOdW/yxCkeGEoL0JCaRSTPhd6pBxqu0xqttPzXU3
0gubdlIHXF1NpLCfQAH7L1IUooVnE4Lkqed7HcBQS5++jD3hvbpgw9FQeFAtGKlcxyt1kc1YqBxB
PobNO8zpjv7BxjelBmiGWNxHLDWl48iCI/SDXOy17VFMKjBPrc/AcfayItTvSOfRWsL2G3BAs3p5
Wh5rhNbNDmHRdiD045tdQIr6qCg7kqYQrSsKWJyRrWpvvfQRCYAC1ZY7Y8Nr4TQVAMoJfhv5W4Fy
heRPruMln6v8yZcM4YIjOg++mLQxYq5g0ovEGSssxMh9eCpic30Q6EYJqXsp6BoH5Ne+D6yJ4Zhd
56ccSt/yLwOT0/255BwaA7np8jmEGgz2z99ejbac8+VpTx6GrXmtlPj1UzCFf+OVMP+OEtLrwxTw
121eTviwRRZI3RZydXCV0BGkJsFgZb3s805hlN8PFt8QQ/CeeFPv74NK9jXPnLsCTNF3dyHn+F/F
PufoIDMjRMLy+6SriOF1rn1ERBxHYDJwoG5yJ2fA9tPAHgT5+v4ag1nMe7XAxcoQANIOHQt1UIyC
8vBAQgMs2Zniq6VwIclQnUj0SlNHFo15xHVcDrToIJh+0noLwPp0DYRSkNMsrJxX51oZ+9sTpTlC
8Bxj0pJK4F+6CZuklNLFG23MFwUf0/q6zrC972Jh4MckJZo/QRjChtW2cP+rbwk4nQrbDBDOZeQa
Bk6sqBoO7ru3KJujQ249nzfd4bXTH0KXjiaRzTwRvUiaiN6bLGiJIodpwj1CH/6g4ioJB5Er3DWO
mlrzgkjC26OQw7SgKFDGRlge3YMM4Wm8r8G+63ZJaDNdMY+Z9RtWV8CTi4mlKwr8A6oRyQmLBwfk
xDm/TaoCH14r2OV7Qk1tl3TrtW+yJHtsaDws18hmF/DYR1lP/K8aQ4Mj78YnJ4ch58F29x4s5rzt
GqYY6x5mk9FIGAVBEpr0FClMWNR5BrCBLWV3ci+o0ve2Kk6qZ8Hmm3XbLXVKSSbOoly3cNdd8rN5
sVDPDkyahjGKfrpBRPK2VuWWpmZzZnI5gQlUwD7LPzKE+HNHCVPblyxBG12GztVy7dlij6ajxmyY
UUbfhIhYFpuEsHic/gCc1uto8OgReWr1+OH/kvJ4bqj1cDEx+tzksBi5r3xR0XT5oEbhsKlS4au2
Ml6XZugHnOBdTXoGk81omqjN419SFZFNrllNVLXrHYfC7nQ8jfpMthHMqMKIecVwRzjMfsjbzNed
qRrhQIHauiFltGyC8lPdjPJUk47G+RgSJn5Nt/W3auTDwFXp3ZBWQIbIfx3/x2DwCcsABR18F93O
ConvBgwCTxFso48/seFSR6y4w+em7JTXEuC4uMc/tXE5/7us+FE1sZJpAmI8Y26gZOPEhj50yuq1
jjY1WCvUxe9Y4trD+mqGzHIidvCETMRTw0LmtpBm6yztbBy8wwN/yDGq3uDVXgjTEomL8v733U95
4Hq8U+E2/+4RzqqZt8vEA2kPI2CEy9UB59zSUos2uaw/ZRBU6PkaLd80F+A/4ltiOU9CdywvQk5A
xjil1IxWV1iTxe9ZSNR8Bw8azL9LySUS17RWcAqvzwxloexb+MZZm+3PL3CKq2SfHwhdPNLCc1DJ
ANlQGwQhz+OHCXuWC0oOGDSCqcQlYUozq5zyYI9UlTsHbagRhyQc4omawAM4TIqedA9xt001m6LR
j8tWD1FGraeGxOgYNcpwXBqjv4IQAOjjv/drfHzlj8m0lnMKwFdXK6UQvlBY9uibeWarQt38WkY7
bpHYmy1Rs4c8sVDZdEun9ONcZizZ3m6aJc/5QDU9EkPEV/pnCjdQW9iEcN/e0Rdi2xIczjMOWrPv
kGFPei7hMRL7hdrlyzwxjz6K3PuM7R1F1kviWI3Hh1K0ek6qTwOhUVv+6ZYECLd5BXIl/XSPn4+o
XAPY6PpCp5KI6kvaoE6/GDPG9ML25MuLMXhj882M5aegkj17Po0ELeXS2pDBm/Tlsi22J7YSxGyl
GWLKXyPa5WQUcYJkHMjM6q837xlQu0e5Ug2yrB3OkifodAhTPiY3FHg+VO9OzlmJY3LCJGJBtyie
AcaUGM9j6zIJu63gGr4kk2m+JDrZQbd5+4v9tVALf8c5cjkMida/vUskj8SaOJlhJwOiTpeorPVI
ZhDSV9+AD7SJR/viQwMJBRaQpTxn2PhM5e0N2Q9MwkZGrs+iU150Q+TmKob5IeU7P8MUhRiOyidV
4kh0AqPOir6Aonm1hbJrrjAvm610I2lUT5KTA6o8jpWOXiwtbtoQJSySnzV0G85t09EoUcPxhDQy
KSFC0jF6yLvywg/8HcMzDuKxGuMumUIEC130tpjy8I4YC0EOhUpKiKxjCNVySJcYaDcXF0ZD/pjU
p1LP4QmucMzMylDlzKPMUAHmPrjBETIfioVmYQ+XE14x1LKHjz60LOBVcO3LPqW67O9lOPkBO+Au
8yr32RyZD/WQ7E6f/GIqDiIILIpVen/NTsWxXqIJwM6SEjhGLc3/Gpvk63JwWRZm5B33bSSLLb2X
PZuAHjHTJq7pGUigL+5wIjifdkHL3qeM329DUr9KWik65sYAH9PwTN7yplOUiUFbCX83TWIhAU7A
znZttVkfdlaBukwr2BFwLVmgyGkSGShPabTPh/Erq62nuLcIECV36RhBwT5wUTos8AH6K8gv3JiK
5KH/+EdIPUMnVx8f/WIUyLPdccbh00hfcmmjhyyPRbzyvVnmz4yy8IGQ3yXtdn0ZeDeQvlPnheiv
Qd25v4FZrv3Q2ZbyQM2mmGprvlqP5f/DmbcWj0dpXNh+qJ2zfDeE9yE5ru7AzfBGM7zahAGB1Qsx
buHYP90N28pQ7k9MkbE5+qeR8VQTwAr0cs3QV//L5tADrmD+RkkeNgRHGHUNJhx1B7cFa4D5P3IS
tWDibSy9fPw/LVwgU/JvfkBzRSrWO+PbtF8ePU+LUoe6Ptpsy6yYlW4awhsjLVRCnk46ikYlCDc7
T3WumnT0c2tq3vnVPFccy0uAXYbim5JtnI8qF46/um/HnqjYE7ypItJBcbmSLLxyUHh6EyxF4HXg
3frj1bCaz5F2e3TQoSmV8c926QJkCMiZF2M/WJmNGXiXKiWtNnqMABE9GtlyflpC20Q2ZTnN8R5J
BlfhtPo/BRp/GNAaiFRo8LKaCJgn6kJrpYilAv8tn3x7KU/zRmliZF30z9mOCS12wsL/fL8f3u8x
Ut1HxI8Rt7dg4i7blXAy0ssDsIHj9jr6cRjDaxKBI38ln2cAz3hCrvptMCqrViIMgSdbczs3cL83
7aIRT0LKmAyYzKZJm/pj3YiyQxT45g0hPN6jY9nGfOQBqBoFM3zFB0qEED2g49LnJ2mRNa4zHeAP
yMx8w8WKWRDUMSuEOoh5eAQuOXmrSq/5544/0llX9aOjMn1SgnKyyZCCMYmZpZqAClEr2m4tZzCV
FdABh2w4LYHKCiJRNhaDYcHb7b44Q7tnJ5g90Ka3JKhBFMd891XbhCZD9Rux7Iu/okm/0E8p+0gp
RIuW1gkfovUHQ1ZEDZ1tony4RdCxxbx1Bf+hkqS/ut+NO9ymOJ2tmDm9D5dOO9V9sxMC9l1Aq4E3
wAIdj0Di2vav21PxVdHDxiMIoMzbvsbkPxNClFJ4EsxXaTRo4yQct5RP54RTf/KeHTDul51bHSuL
LkHYTVcozd+XRyf7Wte6v2oqdIJ+dgj9q74nLKPjKHigFsefgN/8vfHaeV8gQHt0612uvqUu5OiU
+hLs4EZAUsDFC12+M7f04BmYOcUrjo8kORpdfCSH2R+BStUw2anGgMrS7ds4Ba4O0cEVWpph9kll
S1joK6jTfEtjnfXruJvactuBL115nhizIcwuFUGEolptvpgVciqAeZZNGl+t3hBcqzZTrl8udAB5
EdCLCvlEGqPtt1qR+izWgvaKpqKodGh7UG2vD6doVmjxLY3XtHztS+xjqAWtv4MkPD20K5Trx+zW
XT9tcAMzDARPRgCBV7btE5Ta+RkMp0WPTKrKbGDJ8rM6iL8JklExDL1n5DSV+wCzXCmA68pCtJ85
m40hrHJo/x6r32tduE3gPJMptD4Hl+0yxFTJqzMWxFUPUPXuQNVCJsmF9BDdHGcH5pfovYZH1WYG
iSGM0vT+sAezNRiJjhFe2Ebq1VYAShkeW7zpL8bnFpE08m7Z4xfh9E1KMLz/ec41GDwYBBN2i3+N
AKfbWwi/i2H2ZQpNGUAPXHxgqUJQP0ND7TFkBuADEh9wYLFwqzd2mwB10N+R0JfmrNeLc2wAPUFS
4fJ9WIXMHgyLqY0BGpqgDqwxhVYj2ZL9tRVnoWnHlt8eZ4ywFrRAYlrGK54AxCexmXxvTWgJYSTf
jUKTe2Zn1fdkU6hJmU6hDOM/bvamiN9yncek0Vuhy8nGgGkGw77hRz7dHT1T8FIRFV/v9X7e0n6H
El+u/oPogKIWfMcxpbFEsShRIl8XjbCP39SoFyIR+8FURxhSPJcYssrOGLR4gHOu1SPbpFao6DO9
v1VKTkEphMUWYExyxiU2JVzQfVWTfWXQEJtO95xl4sWa/bHlheS9/0DbLXgKyFhsF4CxXVuwuJab
Vl26mhBfJw82Sl+oSp5sVt+1P4fQPvw1l6xdeEardzOLrA1dXyJMYBGFcwXcKcCGg0/LI/UoG6O1
cGefpu2osjCD/5PS4W/ysmraS0dMYXTOCy8AmzgYG489RXA0qlJC1KNC0IA/GC/ockOSsICO4lgt
JexurM+Kq9z+WNLx8iKqILYu7rcBfg6m4a76s4aDADEypLncZSlUMjg6zLU1uVlTiV9Rp+ZAvcqh
zlyK/7hQ88q6tiEtiWof85T0xz2SAgkJ5/ZeackMjtFGYyjLeu07Ij04GMHQQJQfYrVB4Jv6tHD8
afVCdgg25Iky54HvTk/CrO9yILbdJit4VjXJ7907yxJTSkCpz8HCEIFKfzXGMErsik50AtBmqyYF
W+sgwIS7ewIDcIf8pbi3XUrPeyx4+kApkC+e0MkvA0xWjF55wIvJDNDe6jjEJqHoFsP64meyT+FB
7msZXO4FCv6ixXu1v90NLmO0oe4vggaPM9T+yBXp+AzBew6rk8bWLEHONPqhWd8VMeWGs8uipKVf
w0LeSjrxOpWdrCl7vgNorfb+c91IF63vzqLTTik1x34ix8an8Bcax4I7OlWyY3xb2oHeTWtkXR/u
f2HcYsGnGNKB8TTf4sv1J+ol8KEq+5gB06c2gfH94pZhr7zDmdEP6MBwEKi8PVIi2rxy8oT7hdSU
6snMWbdv/Xq2fxtUy0xIvlRrWGLEX3df1uhI/P14PPe6ZbtA7jofEjWBGfoTPm+5LziaClQk0bwY
CTTc45DvPPcESgR24wqoX8ghKMVb5rPXxqJVL5o9c5RUhJO/HoY2VKXF3J4uvg1mWwyOqLG6OILa
VaZxRYDAY5NLQ98xBrFuPI/xfCiwLBaOMtbMuUMtrBLkTJSlgUwv6vIAfWWDUNkaXq3CX00zMFyj
obNqgADp/948I15Jp+VhDykJUDVm/MwX7/Ncx7XECVzieO7AUj9+ORHZyG0NJP/i6Woy5erftSKN
7C+WGamPdP3TXz8Y6mGlU2xA5J1fEdnHKIu2JfK4WoKHxA9mE3vNFTuvkSFnjW8cpzAvQCS9HJHa
i0Ihg7ChpjmRlj6AQzSAfHC8HyogyegbGW/HQ9uWzoFfrcEXihkCwyYwYTvNKamRX9Y9ixNCAHce
WYT03MiVuhhjxZJBvJvokRqySIioQOzrhXGih6TcX9Wh/zSqLefxcNb4SGvqmlQ2aWp2b788NtiJ
Dqy7Etf44Oi/y3RhC/gi+8RqG7DywvC2TzTSyJAlD9N7dNL0KWGSE6WI0rYDkY7EHS5iHWR4tn3x
78RCsASt7Ia7LneHJwm2Blbe9OTF2+cEvkC/CKkWIu6iWdYDVDawNoCzYU757ckCbnvLne3BLW1q
OpDKCE7xnkLoCpwUtffPho/Kgq29MQpJwfWXydClu53e8xLJrFddET082QfxohHxjN+482FS1Jw4
p78gyh8aAF5ssnFRWaaaaynqx5kS7R7N347fMY+2bGI+a6C8+FgGfjV0OcIKHd+i0GMAIFpuTHvH
XGJPu4MNBSMUOpN58WRezD8I2+98YY7XAsOQgz8MUwr/aWhCBDVj7xVIYjbl3jOcInN6CdMrFagA
114IjCKwz7xAAAPp1xt/st5NAcTLd1Z+o1DIDqx/PeP275Yl5p4uAG8mU3LU+eynTqiKuWiKb/tU
q433eo94YhKH6cW3RCuIz3XuoOBbATOUEzZ3zYlhEIWms0C1axdUNp3qfrwXYODyZosqq3hm/Crx
piKKLDX76EbHw7KHm5F3CB44IZ4Iq62z4fnZHp4es4wxXPN/QZYw11GVqVduXeBH047gdqs+RYgZ
8SZ85rAvG94wxHneh3tDjvs801FN56iUYBAgS4Y7gw2Ajjdl/CZG8CNde1X4WQLo9gEK93z4GIxb
FDGDNfC8G7ga6u2Ec+SHz0vJXpTvXGJGBnSVgJQqpU1zvYWL6LP6sQayAp/vkT6BJ+h6fSmMIHBc
G6en5d7bzWGW30qwn+6bv/gqOKPOBrnQrakLI7qVN1OARG/ObfyCIhmaYG+Md96z5Ie6Gg2EegmL
CtNLjFgdgX022tqo3mZuR0xe27WQecpSVljy6Uy9DotvnEUQ/nZifqBXimdEEhknGF/rozEje+BL
9Q4yjwNcCACbt/tVuSMSwrVPbQdqqQwNx+mSXSPYBjUjfQvhthgRy+Yda4YtcVYq5T93+1rVt4el
Pa1RphDidj+5SN1/sSPWxGJnK/MkGrGCnpb3FFxo+Gd55L7cIt2vjhLVqsx4Kd0OuO715YdLn0LM
9pDWI15uIdDJWq+49dUA/4XfBHaBrErE5wm2qeMOqB/5swVnwg/DNmKB6HNHOBRlshsvopwPsQeo
K2AxtdERJRe2sdaLyf8lDdqjE1sSqTVtWQMP2/w0LY0PceRBklfyKROk2BGHm93wkRQN1oQnRos0
ub30rHI+5gTynU69HxGj7OUYyCppYpHxIeeocStGSLiHDqNGyoOdEwdFqOWJ/l1O1rjBi6bRFKwg
VtH4dT+hJNjUn8dFo2q0v8v5jTk7LaQl6r+76XmTzfv+AZjVl51LDOCrlbXhrSJSFvM8Yk3h1pwm
GIaf5ZuygrvPzmzbJdAZ/IZfzW3h0/SlJ+KSsjDmzrGtN0Q+9+EpLHZyp9sZf64wAUbRvvBUi+Hu
6w5JFB4Oty+IbndI377zM5/aI4cSuoyZVqy9yX/WngEyM3eT2OWlVkuAx2LPU/0ejTSgWjWiHdJ6
0MD8eEGDwLB3T5jz3RdNfp2mSd2HPSnFaFYZBIR+RG+pZhllJvB15lJsOXh71mw2UE7tsw/eRPFI
x7N9sLXskfdp9BKTPXpcA3glu4OLMKUqtA8Xr4hbhw+YuROFT1uXHQuM7YNFxfGiaorF2Hk77BLa
m8/ju0GJ8UgX44QckXiCj9fOet7qx4jf9lpV3KICvOUUOCg0zpfOoozWSmc4X8twY3+Vqdf38xf4
QbN2AMfynG8lFCLQ6IaHM4wrC2B2IMRqMtVRypEDqd0Foy5JhEN6tPDvXwIf9Cj4EB+Bvo5YyyJI
HvIqm/g02rVMDN0bGKnq2pCaFarMN7r2cGffJRNKpHOZuNWq2dArPRVH7slNrtyzf16YKfT7HIV5
Dmik7eE2ZzAYwKK0/fAhLZup4c0jDNfEdQi96Jmf7JMOBSiRAdHhHX+Ktz2fH7txcazzOzD3sDtI
hEyD56kAmaaZCc7L71ECxdRSZPg83Czc+T9jz7KVkgwj4n+P52MZticXeDrxTfqOXJWxJXLdDUqu
BymIIBhGUCEg+eZAiLIYoDK3LN7OR1Go3N/vvqFgAcoeioBYq+Zcc58rU7LK05zhAYO/QRIHPYf0
S+BIBSBk1KWFRvCxUX3UDk+zFC+0l2Dp/LIF1LS4Li40jj1Q/T99H6vuqW1J9RXPX+Hr+POMdowa
jYQh/Ng/AXKNdNGevI9RErSg6BolWtL97OLpUb/Rl2iNsNVpG7IPz2xo7WCcPHnsgRwSz1VomOyJ
PHpPekdQYhztAW5aVEAYFzOmBxevupR7LR9ieoh1ALl8OvMEcUhXuCbX4xwosBQAoHN7XP8Syhnj
oD2JvLyoia86gvoU2qJ7JdwtJtMrfcJkXxZJmWwoxjHkfAtJPK3L7O+2wZo7gMv1lJwzkF1jPsAt
6iWG6q8xDzDuhsSc+3d8MLVuA92CGjB2A2ei6lvoqgQhoa+JV1PtNiyVwJJSiUVNjbbV+DaCX1Zw
VsBIsL4YhHQrvNLz8llNeYbo4gB0Y6Y966JjvJ24UE6XmN4iqzRaATDIsUOm4k6ABkdPaZW4oXUG
7xEjFrGeP1SMGZpHaWJeoJVONiy3C/RC/4TFjtIkdUGEivEaYgRe4+oMiD86N82uqBUs1J9spxXP
XGLYSO3Rc7JpxfaviDhiDmZAJl6U4+XSRjcpi74zppg/mqAIJKDkPkALYhTfrr1olwT/H8j/mZRh
shQW2PyOXVZ/6KsH3yu2nM2djEt7jbjpBdPM1AU/L76PKHgnOG56LgYU0jpGzgvvXC+SihiwHvKV
PVtvGJw+mTi1cc1+hQFjRMBYU1K57Ba/12rSKAXA1sBd0n9Z/zC0j49yTNlcHS8+SlwXnApiT4iN
5Vc9Gn/+2ypR7bfFxFt0Lp56wjBUJgiHF2+WVOcV342pHfvsWQvxEsdG6cGqG4L64u6qn9A2LhJO
FFOjn3lS8qJEKkDzGSjrD2cvkxTPUHYSvlcaV/ER38hAswYrSIb/hxSDXTkuRywS7tuxXpIMs1iz
PLcV/XZEenw3QmHG2MyOVM+hqT0LjYqw1bcsDFbQzgZ0U3vKmRuxIRNWerPt74/PqoVISBE5hH0l
UjnhNjB/3aasfKJeAbVxEEpGDMctqIMcO1n5LMbjUt2yHZRpMb+IghzAtUVBXJVeDvI3fiZnDXYH
5NmY9g2u6DcCrMgcbJJPCwKETO7q3z17xkz4+dCGis/TVImnaWdVLO64CmRpJUL9CWf5GH3ut/Q0
8LvePdkqYMVptP+x2QREfGoG52i9IRrDV1oLRnHUqwHgD5EiJZGGT2buloti10XX0atPzU8xU/wR
L3J1RkzIbfFVlp5OQsY0knRGhBNzYkkIZn4x8fOshMf115cwoeh7vphNCNoHwuGXGMyUPZPmZ2Hj
K7uTC9RNELd7Iciap+Fj7PEJJZX7dv7TVqaQ+a7otlE1+DRkQLmc/1n4OvxG7Wn4qn8PMp6bmzsH
Jy59/OIBHq/IAc9+NnhMFnBKqI0ZKj+NkTV4eZ7VNucgOAJaW8uJ3iyVjFPhsDB7eRMtLaG7JmAt
m9lQFBCCz8rX1UwGKdA2H5cfJ5QKymd0meCo3qDeZFJgvdhOxJIDR7gFW24P+BOy5xGqmdpUvL3J
t/eLspJfawtvxBLf9PaV/CGL5oFkByJigl9+aBt5MDoxnJw6k4erE5UiZmh7KdiiF92Dg773fWgc
CbX70BmEcBbWHQBHGE5bnc7d5YGZhjnM+qD6m0/kP1OBYaPpnhazgOHD6aUC/FZphQDsF6g0nS0Z
0cJ2RecRiyKkK1ZHMBD/RncVoWAZG0rw2VjfX7zgI6EgfRLaXOBlS55fl4H4FQKLVNEygcIhZ2t4
JLOsxO8v0ZLW2kkpJn3kMdkgtCTsI7Vqtu9nYJe+E/ILXN4FjO+Ou5o9RxLtRo2RQhQOoong8Wv7
PmxchahdaHXevv2SwqLRxgJSH2M5pHlAV3gRm8w6eEOL4JbVyT0nVurbxwRKmSvTENiYy9GD/a7/
P3/koHkUhQrDMvEJ0HBkIeQ4clncrKfdynONrMvxmPLWfgMcJ8HjI+lkHj+0MTLeJAxfggMeVQue
knju4STMPw17uulBOHL72YnVSpHJ1Bp4HTbspLTwU/Th7iwU/jRtMvedYx3yB9HDryT/lU66baRq
vLAVFGCmOKt5O2rlDXBzHqtrkpqHUYVy7lZ0CeLHYq4yeZPxFclb1lgZGK1ckcjZJYlJVlOHdtMQ
M17YKFbkNFgBCA1C3u+xqDtcMRM/1mgOwBvxY1ABNBvEhHsjG9StAO5HXd/Wrg5VA8IBc3BYc+vu
lRcSrkhU6MhQU+tGM01Lgw7Tu5UVhan6H8Q/UIraUFyteal2JWZxiyrnvg9T9yt1mV1aOz/82Ys2
bP1GKbsASj9dKQPvjmPcCmKtsBbbzkxwG59Du6tF524HxuwZ177d8y1beVJ7/wZfNCNnn1sY5zov
apfece6dq4VsK4MEKBZGquEGjD4Ue+fMSgvIBnC4q9WW+0zL+6t80liBo3EoQ6x1RbB1r2u1p8QA
MeZS7qlaIVDfmIeyvXh6e5Xr8kBgt5xplb1PQyV+cgHuw+mKQ/nJOgO/+IknrbVDhAEUFuUN0low
KXMX9hxTMA4R8v0S2GZWWIxrG5nzrikkbg3DqxV/AdwcWvntUvIRpq88mRseGllNsuNi0vdx/b3v
PDAa7GfQTQh4HBtu2NanhlfepwO5aq5x9SQjmp3lztRfq01IMKChRxO7kzxDtSxDGhjsAyhc9FXg
WVsC1EMZDFe7zaxogkdWoMP39NTWk3DMQXraU8WyDHlZV3DXcDZjigfIRyrJ9LcBhtEr+gIhhDym
xAF6IEiTPSy/sj/LU7I7EAd3zLKVKcBWvHD6d0aJp5excfRhQ+xo5y9liyyu6uanU8zmfYL1jdxo
0CHhJ6UPeL6NPFKDI8tYptzQOgintVwO3Pq4oXor5o19YbeF9dDCcK7amxjygBLXcJyfSN8w7a4s
CohGJVPkDGoDY+ywP4uJVu+ILeALq69+zGyiNHqAuZQC+GyDgmw+Xb1IhaCBYVrREDhUkFfyeDVa
n8GNUQSF+/jbFnBlydLpV4mxs5edE0+xxss8f3EhE0t3/LNcDQwAJQLpDkCazCzd5jJYyipd2DSY
jPz3DhKMR7GzXafcKTTDU5KUgeDdKgEwcwVoE0se6YSd55sWNJAT1z8ADrddfzwTEihcsQuU8gIS
P/Gu3+yu57esJn9qBQzbY02d+s7tsWaXkwZ+yGhz+afF0SJ+zMEQHisxpZlC/kDSYWgNl7H7kGH+
+HnP4fUvcbak9UytyGBK1IyG2i5WbJF4XNVuj1dDkkLf2/R/OkeBrHAzJqZ3kJugIc9ByfcxYhEe
3rCvRYBnAmtBofF49kgi5KxZ3FlQBttdCOJAwX5JvUbIYMDs51FV04I7bxkVuGJcd8oHA+W5Nwbq
3sF/poCpHHC5uMZZBxnbkX1oTVu7rC29X+IXK58532XuTdhIP8syQXdK1GEd9FcUVc+6cgs5fWsu
Y9z0Hrxi4Z9SUogbfQR4U1ryL5aFZ0CnW4ldz9nrtHSUlyTJzVOuC3CA6V/JlMYoyurNfCl0MTWh
uielHD5rrAoI55WeY91njF+VjIDP2bhaHbDVU63t8+74V64Coh3mn8yKpN1stbNua/NRH9c6ujZm
4CLSsj6wlFAvYYX67e9T/RF2I9eMvv0bK7+w2qCEk95XG/CJWlIikeORwpeSDN7U6mKS7pT5Fuo+
UmuqApifhhKgfVkUZ8QHf1tmH/2NF0D7JfO5A/Tx8nEXDmWgZU1EJNqOoN/0HwRn6FF0jbIxe3bs
iLDsPQWxPXKDInKa2Eq2XTJfgOKqg+o5DJIBuv+0Iujjykm2cjS+pfTBOQ0SnWt0KQgZHGWoC6hJ
68jyyn1FfkGscV1qdNvpJ3adIecamU0orOPViI1dznN0LlYu6Savs0iZgJwt3Y0aXJVD7OOZgHvq
/zyDbgiGo0C+eQ2FgQ5n+PQdrRh1v1OrRkltbPNX//HCFBZgAqVgEKenLnp9YedyvTSOE/Kd4F5J
EUMayN0AaiUXnyNRf/gn/NJ2+maRNe7X1uj8qowpW9yV+2M41wxsSRwBPE+9u72GqBl4J4tT4Axf
8e0dzx9Rrtsv0DCcOjLUXMtpFuLwtmNqyvgw6q60HS4QpKrVk3hQdX+HHNScc+qoWc1wq40IOdBT
Tue+GFQ3v2SMDOijQ09k3nx7e3L9Bc0Z7jvTOfURY3AddJToEjHL9PxAR3lmF3nfM/LMrS11mWMO
6K8mnqM0Q61nO/0Cnful2eRyRQjub3+narLrWkqjVL/tPNtoHO8M2xzPhZwk+Z78bCK6gngMUSR6
Bw+Hej0qeCiB+xQqQAh99qEcbOHR2/cdUEr4uqaJ6pmg9andtpfE0V8CbYfbrR+EP2h5MrVOUFPu
6gU2Sqhtf4CYObswbPiQcQEJp9FsLnYBfXFUzxq/82rf1EDfsdaDJLlrWURxvTP9YjK2j20akFGW
a0wmEgTn5t7Pbs8aj942QAEDBShroArAFk7dcpNj5cynnWZqRj+A9bPkUXSPFqzAD6qeQzf3cDsi
FtcBozGjfRy9RwveDlNf/8qxCjXWIyfclnmSieyrj0pemSwufMrUUJmXitDo1sYXHrmZZP5Nh6Te
oRtlzy9cW6oAG1P9w+oeyeknt3spmIwV2FLoyE6OsoJ7qMNdwg7GnNh27dekWnG196BiKhptf+Px
ifsimWH6DqKCwt3GpoerrDXJHYfLBBp1WQneNtsxkKCc4b6wBkovnqD7U92k7/LyarVF77G6ey5r
gGssveaJimBF7WwQsVlbojVRUJH7b/jeRBw5piCSFqo3FAY3p9quko1AM3VKsGBFbc+V/WV0x7yF
0UWQTovleWfU1J9MzUgTsdYUse6EaPEJeCnKDMoxHcZWwzZ1EloEuAw/VwvQC/hdIWej9XhZL/LR
kupkd/JdnlCGUtobkErxGfQRLl11TokWwI5MMcxiWyNhmA+NkSB5mwoqYfOdvTrOGMOP/YnLpy/j
SboGmIjkrNc1lxxkoxH5zDfIYKCXOcubnx9Ub3kRED0VVgIPQisrGzGvfBQhaDWWinYDC1VV1Auy
cgO0ov934U24ESWPnf+slpqdXFnOW/MH6jqTVOQE1GaIaKR+rmrsdAyw0E4z70xBpvMXxzk/qlnm
lOZ2hszsfm8ZQqnCyICJl2v+9P6tKQcOctyEA1Q9DrbLsnVLQjY9Tv2BZaA7AtQG33e00FT4PSdu
oNcHd1X8WpwjD4hnjzegme0YDyzlinocGcHJsUITk9afxMWpNz26ft0/iwjyXLDHuMJ8i3ByZb71
L9cLf0APR/AqffCn1Lo66ULQiYrNY1RYb/+eCrMEWd8ISvUqLWhi4WhOXa4Vtn9ibEJVjllIQlyg
dbp2L/ULKn5NY8J+NEYckVhzV5xSTK876QPZ32a01VfsENRTuacZcCONH9G16qq1OFSMpm8lRd0a
xtJEVc6kAsFiOG56jYX51TyHjMpL/ucLqX2biJbo1UxMAc9u4s1P/kdPNEeWK29TScIE5g5FHi7b
cxWIonPTfdZfPjXjQQeabJ9g7nh0KrUtyzGgwDwirdaFNWA99hM4EsNumLfXLTTfj9dBb/C8ZIbj
6buSZFkHA676E8R9U/1JFlBwzHjyy/tYBV17ZORNaqUQCUTcookpRsoWn6CAIXUtWkwFVx2/+zle
kqx+N13eVZsW5wf8iPWkL1lqZXZN0wcpteJ/NnfVm6rnZfYBHaKN0S8OT6HcnQzTY8wfcakvQw9x
JqK3Y2rmzSY2n4Q1MfTe+51IW2CXsqX/zzL41vPDvx7cLuYJUGoM9sJwj3jnh27tdzIelJuNn2bX
ZfRw3K5Zlq+h1auKVMXCm2j3XH+B5onfyGszupMWsrUOvq36puALjvLQTORSK5mEMHg0RjIhD0qo
f96C81XM5wIM/IAHJIx2q+8Bl3rFdBiDP/NVJ+8+aT6QL/S4QtEnUNxaA9gPJ10zuNXW4X5wLpUj
jkGF6DRPWxecZ87cMYSdd7JH6tWCp7SJzQhq5bQ8xc8UesCswAMvQJepKo21FMTUa7tps5inBv8Q
R1bUSB61AZNbRFUgIchbMXevBVIUgbXaMjGsnY8nh7OQF6N82rXNqKY2CI+bq5qaAPSQSS1FfB5s
oqxPsdUpTyD3mcgPVC9RqZcQdJL47idYwvxw6hTTCCbv7fclbp1DE6xvXGJFQJiaHINZ+8l3g14N
RolBPWvuY9OTZVVQT6RsxCr4UB9eauKQIuH3+Et49TVDKHQzKQQkwL+0ATOcwQf937RFgYaMAb6E
0YWfZ5T0+aBzreYWImxIfUINW2CFv7e/4J/T3bxz6dZO7JO6L5/IwjTqth5/whT/b4LM0ksMLmxC
zUTfNGKTx8H1sBq89NPaTuuBfJ3rI0INIAKxKw6cMKV7pDVJLCTW1hl/dAyHzuxO5Ie2WEbdvgf3
QpqKYOPup0rYSV7L3sKYKJFTTAy/sCPkqfnRGS2snARooFp4qwkJmBucSwy4hQ4XzZBG3VSc6ABb
nS2B/swPMk/DM/2kk2/Sy9QkV1m0/brbNaHQVEOUv4bwfRiatcYbqXrtVFnUAZXzUFxnm3+f2dks
ndValf3v0B481LgTfOMFNuIk34HjbKZ6iy/CDZ5f+tgATEBh8BAJBCPhuMhfSt2WBuagOZGy3pi8
2M4RPmDr/Oo0z2lb1vc9RfYBfiLMxRFc51U4leGJSViL+1UK4MpVmzmgdoQXC5djunMjKFf2cV+4
YpaQUb32197+CSKvLk78RhWKW7fRV8fT4WtH2qdUEwS5MWnfyZ54+QqoiP0FQoM1ZuBYqywuMCYD
L0XbYUfmrcgwNrbuVakuZJYJHa9n97BvsymKt1MCuU7Da3r/yRzgADKthxIF3rZr4abWDQOMXvH0
o/o6BEKi4Wn6E112gGTrqP8ZIt9Tglnr259QTv0UZSFs/goRP9pqo2Lf6xbJh5xxehDQsHCsE9NM
aMDWhn+KU93WgnUdJK6jgeODtOSGx9x+so0XINmJWS+caDDQpfZLRRDOi2w5uTpZa6+aoqJuOyIU
Xv2StQzlz3Eycrho1LsNWIQFgc/lcRu1H+dFGShIKL2nVq7Dur61eby2bMchJ6trQOD89plRpvjw
SNqhVAjHZaELx63XSoUuOLe+KGUMwsKH34NJubokddXdBYzuwfkdDHs9ENvency+T9adysdapTJy
bvqvttdKsQPrA+lqZThx7MnO0NL0E+962G6Us4kUmcyHkhCswl6rikuELRAG7cJdCUpvMkhvCrKt
Y/e94ubxNBHSxFYDB3YWNYFYbGnU473oxb0JJOYf8ZetYuoBf9+iYL82esoDjws6uX4uJ/m0cjSs
SKNBZSReVJcua/UKeXPxLG/PcfChJq6Nzb+qCp+9+vJP6c0c8kx1Mq3djbrspkGhzVxzzs6MLw12
HIvO98TwRu9lI7F+P6WWi/ywcBhsAFV2G8hFe+xT1XWzymWAdHJWw+irCyRLSu4rfzA2zQFTI/t9
lZ33NbJEXVDcGoCq/yBUEt3ozhpYOoS/M8TWnQb/GQ8fqFo/ihZZZuBCTZY/B9/AOpwSCA+jUu4d
oNGmsEUst1wCjzmliIjt3QEL/dqDB6CFDVLnBLuXX85Ry7NL5M0jQhYwFjCGU5Cs8bm/PKyBN3hc
R/otM4Vyu+agDL5O+nciWiNqw82+PbD2h8xJFbOY3UVmnaaiNZJ+ni/GJ2JWF4ZMWHhCA+IxFPkX
+7QMkZWhbWCHUTmzqs3ZuxlJjaQqTbEhsP18pEkA5lViDQheB5YrnXRgD46TT1FfMp+6V8hMmGwj
0srkvvGh8NweMTNa+GEnG8wPNEeyxlmhhoh9wmQuIbwEI1jeh62csYlhqRBBDJMOYUmpXauj1lRE
Xe5tYhXXPs2rghHJAePv+rty5vvF6EsGyIW+6iZHdrcT7jkc+j3zIjLZccS7Djio5A8+rJX/8wyx
Wup8H2sU9X4Q/aZjk2G2OhB2JuL1TlEH9Dtf2g5pwuLVAdNIHMG7CX/hpROLZRrsy3gHy1UVCs3j
IclX58LDdF3SfuDx7D0AfwyNkprxFxRXQtzlr6G4/kQfWorv3MNf5DtycN39FaUvxdkJH+U+c5JN
pSd8/k7dj5Mq8mlW2Oy2rLK0X/b3KxBLMRK7CduuMMSmeFshL01zkuylLZpSojrFn8oehxfUViZo
YjZlTKCjS5leKAK55065xCl3V1Vf0oZlrftSwHnf3lkOUqCLvqgpzulSxcSwKyMWw1mYUHFyo9Nt
xODM2YSMv0GfSIIWx9kR6EGGKQyEz//4r4Emp0TFpPIxKSBhEdpbYraPpQVYJzsD4XWqF/3oyRqk
BdzhpcNAZdaR9Lp4i9eCBTehd6TEUuzHDKlOQDLdgjNhWg07BV7sLaupuwd1vysJLY4D/cztkGCY
oA6PBLruSvvAai4q8HIhYfXDDcFyjE5+rTnd8HjBoidoXtgF9J8sa9ur082Xwdy+UQOsV0CgEc99
IZhEQ4KJpHZvXpJ3en0pOYv6hI3V3O9ThECcetst0dTT3hCh7nZtOLCiF4sxK/uIOrHvfdK6PruM
D5OV88zxPV8Q0+qtL5p6no9owmukRgGNcy5iIYRHL3GXK8K+XsqoPEWDv8qHnu8J5KszdlJrfOL+
2cHW+rLbfkOA4QoOxiAOqNXyIo/bOejGaLBGsjoVqL1kyQVFAgpg8cq/4oD0VJt2UqmQMXLQV2zB
QXuAkA6mpkR1E3Hpq4zNwYo7CX4YUT/jgIrZyvWgBomo+Nvxg8OD4lKbVgi/yKgXuWFrnMEiJ7uP
Fuj08sL0a986SYObX8N/zJGNpYhr88nuB/gkcQ5y50LDhHjzISC+GTa3muSh/KFo+CDtw1rDsxj7
k8qWls0W8bnkNdHSIeQaVuQyJcm2bmviwDbxOvvfqd5T8E8YFNCWxhxOfugrU3GNdzm3Vzgep6cz
QxE2D5OLQzagNmFeWTdI9Ng5bLnG7Iy7p5nK4rr37EprUy0cmGsXamQ/nYGqGVGRAf3qKWuGzcSw
Uyg03lyIFQShGjEJNhLRp/1eXyV947DK8VsEC592KLp5LGuwsgJfY7PELp3BsQtucsW+cSxFOoWp
FqGRMe1IZIKE/ytp47d5FdcFNCbXkVfd/QxJcX6yz3e5B3BcCTLstkjkOQxn4TUYIDX9O8kkfgfM
AFveCbrwyQRcI2FVz0BTrad/qQ6xmd/XZ5cju06zFU2Dl44C4AH1aRSPHju4Dom82LLfZHOOi251
Og/kSQVmZsBCqupLDdIlMDDgHRy32XJUYm3OBeelVdpJKzBLOeBTsD1yDJG+n+0z6IuGuOPK8MK5
HUTSyJwGGQXmAiqyPVhSDGxosdS2B/LLtfh+ClqB4OwztvsEG8DUC7N9hiaY25k+tJHuI0RoJvAm
1quTJQFNXmPOX3yLawoI3mGGmZYQ7zj3jBuiQodC5k0fHKyiBIqkURPhYSjsqDK7eU3zbfuLlbVt
tAwTDoY4wFh5YkHC3JgTbJnU15s5pA8hM390dXXYJv6I3TCvHYGnxl6V9N5YAXDpsEo0Udt96Z4w
ZCDmWkyUtdbjAi0L/lWBE0PHkvXIhBIyU8XMOuyyiG8HRNCOWX5xskSDasrDPtqpNxIdiXN0b1Rz
DBkt7Y/e4PDopYVMn0IokEVzEP3gowNgBiOq50lnIWoZXxTDwF5aG0uyiAtBaFMNLd54qLopDzM/
CrYz77sZjRv3FKl8E/0mNHa7Wef6mL+XY2Am29HlVAjr2fRaXwQ0+ncmMnYdloBGBS5mw8+228K6
pacq1VLh0ZePPZ5/+Cn1vORRIbWsN+aHeLQGc+CEhOubnBK9Ov2HrxcDBmmQUfPaxW5pUc0P+rWO
JHZCEfFQdSdSZDGvSI3+FgeArjMB5qZs7NSBA/BYV6BewOGPv0ZnJ2zvHbEIYxjwxumYjiuzFUjS
0svpLbKlk48+KD50mP2vr2M51gVuPCCQY0XBpzy+y3HT/4KtTkgsNd1m91tUtW0BH43PR4FEhMpE
S0jURE5kCGuJLvKOpEMoI0JcaHtPdrJ11O3UdUNBRSBvTn2GbFX7V8LKURB4yVOaeLjigPVavJ82
C6Fxefl9C/LPVc1Racm8WpM5EH0Q1OIe+OLBWy6u21z/UTmCxnC9J2p9VXW27XKt15EHuJmvfXHP
vsBMc6puj1HnA94raAD+6E1iEFCbQ98mmOf/DD5htlzidon0sVLYAnaRjJ2g1IJo8sn4GBZhw5CQ
hzdgH8FY10d1n+O1mY/3pxHUXuKIQu3jneYbyl3ZoiUvjkgQKeRWE53Dgtmm50w75sYZE8QIH/fb
4VRQFH8DSRdjLrczDnKhUnM/SHMaZjGSoQNcZ1lQRaB1D1W1NoXKoNPEsqM7pZSQUNzEl5Lqxi38
v6GU6al9eru5zmgB+mU4MQxzKG/508+crLJgnFghMWJjel23Bci/ZXT6L3oKios7QWHBIz68z6xM
cSLTgipaClgnV0ysPvp3+xrYK6p4Axlr0VwF8uci7DPLZMk8901+qBeDM1nUdM6mGLvOag/MpYG6
wc473oPpg6I2/eWzsoZVagW+tkxHJA7kwd70LpvrVFyhgJeJRbttUIhK6eTC5/UqVx71ZCZfAMpn
SBgoXjzBOJvr/+RF/yw8y3jmxE1hTtd4GFy8y8RNuGUwAi+ktI+dNhPbpYsihGRaf8W/t7sZz0SD
cDv4K9vl0scLKeladOVoygVwI4Cwmyvuov4a57WuqTrnSQQKqw752meJ09QIZ6wKmUy/1d1G2Otc
EEnvkF+0dx8pi6wdRa4iF61nbZX1nKc9amakGRTu2kmX28upFA3ttcShduLKqCLJ2Nj7q20BkbM4
PqfGG4Kt8Aj5kK5lWk3tRBbVBY2zeY8ltbaUqz9tznB30EsuuKn90zskVl3JSoLOUvZrIkeBg7bF
GVD1EVI1ghwxc0MsTjZRckWJPRUZQwQEKwOPdZeGx/I8BjkEgD19VLY/RVYtJ6xnAa/axacZ/ne+
+vFwRpHiqpUcvUBrwTlDgxswtIBk8eATc5ZwSxKjjMMqefAA8A7bK5CVb21IUq0ihr+7nP5+QN4A
sxfIZ0zOiiZLI4UEoaWUz/CcISwEmhiiFVZv+9Fy2CQS0qbvTloQUzCd793ataKAIkn0YnCjERZU
XiGOZJHFYf6ZajnL208fEfDmROQbDyPd84rp+OQDgX5MKlJbADAIAVIUzu+AFpS5YRSDs7kriM1o
MDrzRQ+tSDJ0jR4yV0rWeQqmJVcRWSqgifMuyXaJXCd3w+zuQK4C6/5K2HVnGf6vbFh6OFf/pm/b
I1nyjxiD6JzTACMQAPMgPepLGMcJtX52QpSGj9XP2359gI3v/SA/Ejn1iX7ZpbKCnIUoJI8X29kh
DtS5J9tjp3/pPGU7H/Z/2emnWW+G9uHQgitdLNjb2k4lXLvI/rZ/mEgegZh3joVlWOTz0fSEG0g5
eXIq3vUIyt3I8j1X4IpJvUZTkhnmNuAwQTEaG8CJyki50I73esuh+LjrVZXIZcgEyyJrIWSKIdpW
T0CtRr4JCK0+6yQe3oZcfSpIeDa4ztrLAsAkobZGGoyTPDvU9bTqwgaN5I434O+LASf03K0CgjAr
zh/9uD4VTEvaS3LgJZiTmP0CgXtJpttzDtO2XJ+QukumLQgy7eI4s0pGLNXeCsF/9gLBUuAPsko2
WI8oXKaeNNuzpKT/TKuTeeJ1aBbsz1AXOc3IVI8Mszlg7ZpueCGS1q2TZelbwwH/FNHOOQtog4yS
ydjdWNiiQ8r2B2O9k4e9D/o7Sy+s6JV+PCWm899NZZWQreKznPXbrJZ0GK2f38FYDYl5oOGcniu1
oSbXfYftfLQIPlDYuQacbtSg9BEBdUagZxdo5RluVmHfS1st59CCyCgQmVbWWHM9KRqHn1SJtAg1
pqJOe/x/CDTP5pOg9ubMTle++kMp7jriOgIJ8zOMWiiL2G3RwwruZyguXjXAuDKHX1OHXpxGD5oO
7b1Dt9lxGFHeNsc9eV+AsMON/9YemNt7wFkbWdqWZ6xmOzFTSNgHPzKDxedbcqruK/+ml3+gF6CW
FwGlRl2tvbmlyX7mwqvSfF20uY45uv06Hk3Rs6OXRDoo5V+O9dZC1Pdj9oGYaI1692CzgvAN6OA+
fwZhtqwGYhKsSw7U9c47wtFi9Y/Rvb/EJ5efwPnA5L+NJ0Va2amrnSUtZEU5db8nZSGhBRiZ/zyz
2dvqJxqWLEzyysgDaoqOvB/W7EHlkcbxmx3lxiCGDUoEd5wU9HwkSxhWjVINyVfmfQxatxeXio3y
j7roO63yemDC0at86Hpc+HzCRtDpbpiVnVnWkduKHdQkAlzrWWT5pV1pIKQu0/37msQWrXU0FxAn
0im8THcO4WfEWsdZr4dFUsXFZQvgTTdrdahFSLjVysfp54/YjFqSfYMO4Un3y+o0wIOGS5Wfysky
0T+x7C0ltfBHUm01CkdoyiMEUJBQ9QZJO4z5g6jm91s5kD4eJFz2o/toohBLntkzviKcCH6t50/K
bLPv72zlP2lO4JUnunLcYFAxFYex39M+gBzRPm0ahIshGFzG9L6BNvCzlUdvxVaGxS9nshdKwsoX
1dF+Ggxg/OCgvsWCMj8v2oi7T6+rGbnGhv2BP5eeiP3ARRNrpBi3MniTV/Kl0o9N+fElXkqF9X/Y
A6B84AJYYg+lKTpsHOSP6k0bhDj5va7Ozws/6U3j7ADIsBlSNBUCsBraosUvDYPng3YrjRLU3iKX
UWoYVkBOGKAQwtafC6RgK7WCJjeuCzob/Pbyx9wh+hcUB8V63Mxxexmv02oPOXHOk1pDGDFS0ocB
xefywHpmqzASncdX4cRUju9BsbOW2vkj5Af8OkLILYNM91DSKZ/uF/CdOciPmlGxpX7XP7yiSN0/
J5gAOcaAMeA7z2qRcvm7IOKA+mGgSiRsZeZt4KfVTI3CZ69lH/nimED5quO6gM6crhPuWpfGBYJ3
9kEmMDrZEC5rs47RiHi7Fe05EMM/Z8F7rMtMnC5301cd4HIWnPU8SC0BhGDYnfj2MBt3sYsy0NNW
03zVorc/YLt4sfP9/yl0UB9jtOxbHFbo+3PmhPRwv/C+xT2VzcVgFdgY+m7jFddujZ6ocRl2pXlG
H+5Q19vERzUIO/QbIOKRV/dX9EL81XPQRg66p1QPlMuc9kAWciMOzvtHqEbgmrr5g+Nh5aTs6lV0
TMYIAWbm60UF1vABbNfczgYFcyZNVBF2Seiel1ZuDlZIwdqOVMOljymCojY1RhlYJOWBHNWK5DZd
sPOydR+/K/SaxT85Ad/vi8IPgS5ngRgphDAkexhTpU3BOVFzDfG50N5lEB9ZAbUHszgFWYVF6VfW
QeVp10ZsvChL/jhJvY0PnCvb6IX7hhUe7O/wb3DXOWpQXd+sSZb3x8lcPkQopuEGbsdiq0MHpdiD
f3ZmvD467zuFsm7P/yHIA0GisOKUPNxm9LW6sx7gsmlJSUGo1YJI02cUoU+oxCcF/GecyqjIldJc
CE4VQF/+bfLV0Ft453+zZgiEu1/eluClyhpRktCTHDUrr+C0zsQCRG4KPh2BoeFwgqNUdbUcwoUF
URuVQjDSxxQx0LJ0TxvATf9cBVgJxY7+sGg08u8E996TcuXIVdcxONoo8xUoXsiw/G16drsVexir
goToKt4VyboyiRPfc8xTE7rARIJbelVYF/GZMjqyV8Cp4E7QMoXLrYh1OhusVX54+mUQE4BmJWyw
RXxJYTqjF//tFOpvnyEdC8T9UNJ5qCI8pvdyGH9OTXYNHoLotM3rgeMz1oo8wrn9ImZ1Fq4nHb/i
hHJQXKJKVEMydV400id5Hewg7mkXqakE0pxLtyspcZJz5fJ505N6Coe7za3SUb3JzeFy7jIFXBIg
BgXJJFvPfeaxeBvDSEe0FToAw06pqzLwdIHZ3tAd0Wt5HLxjs55en6L4CCd/c3fRD+yKbz0ZFjDH
UGFQKpGdzoeQwCeBo2O3/rRC0x+edhNZu9bvWnqWNnaNKUv89YT/sqNntc9qalP8SMiYHNG4bsVE
CtRVG3tfQgoxtsstEzKcSTkitIRwxFMyUz4oMrNFOSI3V9QYM/aUw4/YNxr2c5FlZ73FUGiTr7VY
jKJejAxqQBFwrxhK86IOrW9wElKhN/6v8Cha+WJCXIlnyIllfPqKNDqdDtgcnn7NFcmfgnIHxuY0
9OoOMqLw5VFo2ZxbxPmYgeSwhJvR0PyUQV7O4WrEgmJ6tJhUd5vO4maVK7tn8TgBvDrBjK7PCKrr
eKhbMfODiptlvVqh2bhWSI753mXvG/itnc66UvX8dC8zfLE9Kpj/vNqTCxbC55NffCoV6T3fQD0C
UXvM1VKQesPuD6ooeLY0aMswOxkDI3a3JAjjBksPGS3GmNL0598X7Kia+gS5gjKmAGoX649cv+2V
EECAyR3Qw+CfodRufCpSQjPtyungylg5yLRELCseF4UVRHO4V8mybPOMumL9SDeF/pUkaGjJlYXQ
+LrnFzW7UE8nCNTxxxiiTOW0OBH/hiSYqDJIt75sKbM7uzVeD6cwzOTguELWezX0/pmXgBacZcCB
fdybZ+LJrrJgGVq39UX8+zBfP2XL6D3/IknSPf7iSqevVM9KVa3RNbfCDHlkXRZF5Is2y9qlXaQn
ctDJIQHTkWaaHRFII6KJCKgvUb9DSNqR+nVsu41U4w9+onm5mppkLGSHV7Bjpq46tMvBQx/waQoW
8H7SDRtd/vRGRp8m24xIuq+mW5zOUlZWdIDB19yiE9TlogCa13YM4HWUWuxhC6JCuIL6/4vuBrUh
Eu1BZ7aGY4LWIZ5XJrjrYA2/0fkjbyvlBBDtyaQROHlKg82BxHAlv6UjabiaUASH1fHFsIOIbjLB
bDhODAPeXjEOMUm75S2VHmjfYZLmk0ToSDFpqCcnReZhLURJ89rDNdofaCWOIeme1XiOpnTWADWe
3gCo3MWCBjtnlflJYRJHB8jnussB91ATUqjuFxJyPY+RR+tPkmEorzMxt4OSNDPnbOm0aX6NyOG4
hExfIox8f3jp5UlHy6aeHtSaks8yE8vU0gkoJHBA3pq2lD1KuHLO9zBh/cDDg9bIWQzfv4j7PfPA
MG0u7JJW9YXXqygq6n3/0BIL3DRP5qKgHOYpz32wthOJ8JeDv8CdyS+66y2ELQvrcPex1LnmyFAw
YsJNU05m41KC9FKmGq1Yy4E3P3ohXindupw2Vu95b7W0ZxqoJFCjlM9K6TWqWvi2j5Q4TiM3CLrv
BSnyhYUL5ICtV8WaKbGrRg9uea040iHlwKPZz9vr/KjbY31hTEa05hYg8hYTe0mBEcB5aWtjVVFW
rCL0bKSReQP62oaIzYV7RIYHJDAWNyIIp60I8BOWizGNzWMyN9A1v9YncRO1L1Yf+AZn99iBgJw1
iG0lJO1lh1hpxppPZYj/wPnQM2n7t6yh4lAJGH31D7oSTj2MtiDsJdwz+PmKRO3323L76fa8nmZd
E9BGTzTjbo3yojk+yFG/Pc5rlBsl9g1Q8iBXjyHsqW6BU9olLtS4IBnLEQLyi2kRHFvgbyQ8GYyf
RYill0KR7/VDtgB0QIRFdxOJoPsxaQR1XPpnNj1iRZ5oLKEROHRf6CRSdpUKBnyRS8dsR6lM4O8P
I+lOdwjLsys8aVF/kGglL0ocNRAem2IwtRd4q9PMTGGjCMyoSrAE7dxiiFgVPMNr/BO0xsgp2vqp
ae8AG4s5I3xwEGPrOtoVyv1kaUaYJ8y44WpeOVZoPXlKGxQs2D6Yw/0h/BY4MS8NyzZ41PHlsbL7
I0yN1ylR40zpC/qMZOR6uLjOG7w+dS2M85DRJE3zWDZNj4lzNPTn4B6f7zV6O4f97WtBwm3jFZpY
3ZZCCQtdDfvMwBq2jlZZJ0960WaM2U+1ASPEgcvSzWjJtQsF/m0C3qgt5jMMEah2jnyDo5cWms2J
1qSDrapvf7LH12uylMSrCqxHETpGFxtNdH1MLhMiqMeOYC6BGVxPTerwLIAqBPOwtEjJ1brxg+4j
RI6xo5KvKzPF4RGnCLcYBHQ1pLyvMNapXAqu6ZbzhV3ISjcvTYK2olvXWrDAw8Yx/3QOrGQ8EYaT
RCSDIWSdEiaQgns2qrMGGmE5axwpPFjny3m264walj3boHEPkmC9HtnvPmwyS5X2xZ3/ZLB4jvo/
mK4/9tbHLQeqpca8owY6LrMBfhQ5qEgqgnW+r5Ret9sAcbwHCbn7zFJpKGPVw2IBfDldfZyMiqxM
mH0/aYAjBh7nk6MwgjDYrwhFIZGn5PafN8iIIV5djE7Uwrw/NiFHw+gM+WhWWU4QrFdBDDeygh5T
BhHnVY1CeKkI3ab1FdWkSyMmm9YPwKaTirdzQoV06q5zjUPEA2qoJVbRx239dlO4HTyzUDCwOu+K
FMlJMkatQfKp0Bj34dAQKgVQauuKnOIFlBFOsNw6hzasCDQBHA8eEUrJfPDkb6A6diMlsH6HPrT/
Ha48yT1LlJYp7IURYFWs3JqaDpEySqTmsYu9cct+LWYR9dQ6TCcl1tlgcj1U5bAi56UWhXu3sXZ0
jBzrfV6yKLP2CrlqSMjXbFUyuCMyIy2UIUa3thsanyKwJZDCbuT/n4fbHJfn2gcKO7dhNOugVSU2
yyBYc/kMpG0R9Lbw1P6FUDKouLkdhXr6RrgK/F3MGnrtQnDOTxZQ0nZ25/vrYw4CQ0zDgPA22II+
BbX9GayCxipfd22f5VlL5NJO/xGxe8mQ/zSG6inUPpp+urg0GRGAsznG5uXynARruRErfes+spt8
2UrAPSG1W/ZrkzW2G2QmA/SP52O/j8KKos7QSZwVHykfp6OMIN6J8Z8GTnvBOfDcG1ea5fHh0NTS
pUjYnfqIDv9jkq+nbxUZXcOdj2UzcphSpqPKyho9RhUV/gJ2Ksmu3X6b4Q4WXOruVqT1xmOvl204
dsUacHPeesaTGPQHF1feubro6GQNi11QJ2lH5mQYPzteg67HXF54pEELW/wlzwXOM7FTAsdXbTcC
jOmDHJV1np+vQvkwxIkMx0mrPn/69wJJXte6K43zFZUi3DF0yuYbc/89Fz+WCfUbj+nkfSlS48uF
MIbbPSJXryyMI2fN5N90Pp5un1mQcjM5JAr8KYTUaE0aCMX/FrByWtFcu+oNK3yV2KOxiIVoWFhX
H5TIvleYaG8vvLtngorA+rVtaLZj2xE9rQ0xx2YLphRHF1MyPIlYzaUJ+YKingi2+9xLOxkV1wj8
d306OKqtJAbxdSrZKYmKxhRupkqrZnvCaiev5OgVTujWGeRs9kfyrL8HaeL331KCn7HhaTFaJskK
XJfDD+rQFCbbplXzl+tX5LcRlMkNu968U248eWEOb7zFlOhZ33cDd/HbAnZAgSEdlvor9OxWyRVJ
jFmULzWx8nbNvbpehpbsgmcwbVvAc5UBiYTzaB6D+oLoGpfP4KzsTU5vi/ZiQ2pm7XPwLNQe7NBv
6FSrT7uFUkPUq0GoD/iLE6TQ1P4sLnYHAqiAC+jfLF3l1WJZPdEeLP/SOFF6qGNfXGc1n/omKT1g
rkQurtEWUIBeJd8K8XPtFypzQRD39tsxLk5b61I8WYvpbwOvN30cXm9tmUIf6orfcMFTXfhLdZo4
0I73xf667wFLMFD5F9uFnmNsQMYZzx/seTKIkoZ2YWWqVr34R/eUOkN5Rxg62yQKQakeym/RHbqk
6sWycUL9bOfOLH4U1dKVrcsDR0bbKD8JckZRFgWzrv2Ks8KwfjdVl16IV8QkJyiVEQBZUeDwVt6n
Nl75bzjzPcKO1WBmj08FQg/50hZEbVQXPafN8os4E+52VcbgLfuP81ah7QcI2wQ5qS5BBjX64alY
akEt+biUsI5+yQPYijsn+tPB+HKJylxYYL7ntJiAHTZDuogL26+HO4OVKZaqWh2SQXGOfafOqC05
UPDBVCieY5Vzt9jdRu+j44IoJgo77IVQkrY6emaOEpAiJ2GzUgef+bqx/8WYVzlnxSOPRQdpjIIr
UpagR0WEHfGORGJLc1Ftx2kEJRFfatnarkYD/vHydKst9BZuXvPXY8qGuJmVlp3Qi2M5teXw+RZx
xclKZFSPKeDFej4X89Qf8unQoXjcgt842jFy87eruA0dA2mRWyH8t2P1rvNTk2bIpNCegPOz093Q
LyjjXI8cC/gb8XBfjbyrQowJ4jC0aChrvwUsDu0DBj1nqBmOxtDwJXjkGiNlseIdZ2HAXjQvukiB
qmPVc5IzwO7UMfGs9/qK4H6McViuY8fkJAZLn/irLawbBa554K7TB95td0Pc8oX+aweO0joGDPVW
6kCSOOOvwqT6/a8athRDmrVXN6L2SYBL/LMpgeXbcxN/iStGZl1rCYX5ZY51i+IKLFYgS1Sw9kQd
GSFjAtRUkB4kIfy46pwy1vgQAzzhqK0RWWtNJWNZ2JVCkf9UfQw40ZAukoV4h34XmJHkNJCKX/KI
L2nwJaZs9XahFclBF88NoD1sc4YcZp2BVIcTJZx+Xt02Iirq2C8nfifrdM+rselA00MyCFXXuXSl
zyc5IKNBTcPpZcVmhL2hwv5HOj3+0MUMS8xREZJcVQY5D45V//FD8CyNA2o9v9T7B4veqPe3O8XQ
UQsi4ZdnQS5NJ/xfEg8/LRN3a9UNy/5ovHkB0yL2DlCcHG3gT4pZT9NO9SR/y7iA81YUcX6y2ZTi
OBC5PbzDcc62en0QHfHqpqECj6LFQDW4lLBPwmT9+m+/CcbPIgyXWbgvbOHwKfiuiC3D8i4LSyj2
shbSk1zvTfrOV8oJPomUirB6wyOYfXWjW/1UfEqejY/LI8e0DA7L+UBiiLXvGKaRJt8OPa6+OElM
ebmb3C2HEiVV7ckHJWsVQjSMn1a5OplM/CT6yqFX5932O4D4PEQX7pqhss9cBVURiq8B4k60Um6c
5u5eD2YtTLfwnm/1m/s8CAdfA5iNQopK/ZT581Z042NDOEyQZxaYQuKk6Y7j9+ATeKxZpZ1LYMYt
AQrHTvNxzJDFfcNdf011TV1Oj2PzrKfbBvSMUJLb25rc5rfsfUXfhQvIV+fFJNaToPiFLT3IvKhj
ixm+Lf0q2qOxPYeQwS57fq7XDlepuUUtEA/yE+bGsekoVtQXBttc8Z7syG72Rz5S7g1hraLrQzE0
f/PsunMHjxq2ikpgmQdQPOUdQH4tN8Tc6oNoyfA19fKnGsBQDVz8gBSuHJucwGzYULNsfgTy9ooQ
btcVYDR6eY0IShEVtSYS39Ta9h18B5JYcTnMlP6HBMOMWkvaa6WYLPI6L1Xp+txF9xvaS507YVJt
OUUGfXkMAlS7GSHxrfsbGFRR4NaUR7jyHEGA+rYx3tZw3aw8WNsSmeiLe3gQXsJS2zhfy/IBbJzn
n0s21OXqXDteKotMUXIWKiksLqoSZMVUw7easrFLiI5nKhnAGpn8G18DI+gREAURwYU/5qIFbd9Q
NQprSRSnI54p25cfXTju7NGUkfI5edZljSvT7z3FrCU8hv87XZFnW2HPp7YV2Bv3Kf7ce+xyzgZf
7EWc4o1WlW/oByla3ASmjtElHoTraCGo3cxHv4eAyZr0gXT9db6yEQf4IALXdkaqkwbWomsF1PbJ
sRNzIDIPg+0GRpO2+GqjZutSJhiVrXsUw8Ubxtako/2JKummzmgSMaFbfPcL6PIV6lSrfepMF5+e
wXMSHinl+BHSaqdTFYsy9VnqOa73rLNMWAQMvFLjc/i3ALczR1IEsF00NZuyBeePF5iGDd+XQIYj
J5scRPdcEwdZK01D9mjT/uTiM3JJKrYepfLOcvubtbxcg5C2GP5ENAbLyErh34bEjwxHYMXuQElj
YHTJ+o9+6bBfQdxNWBrL2WlXdCZzbVX8XKpgOdViXYcQmWTest+zNLomrg5u6g1eGEeTbKdr57UI
4XQC5w4KT4+CXu/2Q4WYXvFwAESYqjsM4WsGbTLEIiZ0XwwtyH3fVa58yFi6uRTRBdYNKf50poQG
fwuBkF2FhdB19kDSs9z8Ir016niRFFe8yFQ+H6RdAwZF4TA+7tFsbqyPprWS5Qk8SiXe6HH0znXc
TiV3jYeCpNHNpo7yFe3xeqgsf+n4YC9t9odEtOtovITgvy0ZmvqbKzeypIbTX5SzFQKgP06od9+q
VyqLCgcZplNtQqblehogzJkMcWDUxP/XuW3ByNppb6LF/Dha83rfNhqo8h4B1ssW3KJzCPqi61CU
Yx7ZwNeVSDLpBnC2G/8qafZPHchfbT99ajX/yIqBAfdRkELdqjeaQ184C6Z0bFDkYolIkmERaG++
Dqfl1KQ0qCeWE41tRj227GKkXBsf6CsTvONJ4/XTdLRCM6HhUQr2Kt62+Fzssvxxpqnx5nTqt8cg
fO/AKXFJVD8+kVGbeNZeF+yllyjmFZlivlSz/pj7SF7ZR6WwF6z85sfuPJwPZEzBl+zntcydaZpW
e/tAAQS7kgORAbETgNvYdakl+qGkocoZtNf6YPyDI5575ENffjEmojrTj5hu7y3J/syFrzDzBRcs
tRGuFIGy2KXBUFiEjnJfqMkZ3MzPVoPkSQ+YooUFVjSUyIYzvuMl91BamqjKVyb/Ju3UOnbvZib2
rXTIZD6oUy7YHJ5VWRSAbPnABAro6jUhdAsbA1e/PM0k9aGHuX+2dlPekRVNJWu2I//hWxbCG0Rh
kw+NiLEfOOFhqWA1HLc3orB8FuEgCuw8GD9/9V7isvrjMMfnNd+WnZzKYjJtV1YgSUiyotbllVWV
sJbHVc+/AdmkZshFMZ6v0g/cxfGPqhvDDsoTv4ZAI6qJR9WklPEnGQwXvP9owuSDQw2UPjzOmK1r
EwLxOXl8pDh268tKK+nh0u7nPicZL8wHl4wDfe/fcgq7UJO44WWAWU3dN8G/nsEIQjncckA3AXic
eYL8uheCUlDiesi7f3si2ro3sOPeartqOuepVf8X4slB6HDXuFBMNncDCPFQEtdJMYkWF8MZ3f10
yoXlm/uaSbetiWasaB0WdnJHjCgRjEtQBNgXAWw2pkaWPATgBouk2jszcwrMzhF2EdO9m4bze6vF
9AMQR/NUqTGh3OI5Q83x9r9J3CNjzj00nudzDCFMvqB9PGifV7QFNzo/WFRfGKoz4eK+B5EpTNN9
0S9o4Ah3ZLHB6lTE27S29LHD3rw1FQcl2EYnc9MMLD/AD8VYhMB2GkyeXMgsnfAD5YXraQk4Oidk
w+GFWR3io8R5wEj2R1VElj4LaaihTOJ/cJbbDj7NxSPJLHH7jgqbfX7rkLtHbqlHuLNdRYvGK2+r
cNQilyd82xY7//06w2Khl+oDt3MDLg6d4QXOav0BJq3P2TJrE13c7Mjhze7jJyOhmob9/ajj7hZT
tyvkDPrY4UEJi2Zih2yrjTlf8Qnh8MJaBvYTNOiDibY8cspzTTC6YRnnE8H5U08l/3XQhPZ49D8M
Kn0lDAs5mgQrcOS8Y7xCyl3H/pWsXhBQvC1LRDbuPF3olD1n4CDeQeK9WPv4EvFjxS0b6kGupgEg
0HrSrSfUZrIVHjlpluUiQWjWpVL+HCFMDf3AhoY0yIdx3GrLGZnGto1cvxd8hZSuiH31zQiaMxIx
UrSpuKCs4hkWZPc+fWU0D9HCQq46SMONTre6e+jk5YRZ+EmVEyj+6OB+OFrVdDA+urg9Xq8RwoJ2
7XY/uh1T+M1IIofFW8P2D825WKpFSrpfqOCeJ3UrTCH7DqyOU0+PPUV1eB+mDLe3eq8hI2FtdL6u
8Hdw1G/4I5zWUW6mKs3HKLuxJzr/EBhUb1ifL5NMo29sFYb6tCyCNs/xhrayMTCC8+7hA9FBcR4c
2AUdZ8Vkwdt5kG4yT/nvkYeUXzr9/Nz8FRKexxfNpQ+IfNZrnbQec4LjKwhDFcGbPK2jFQiQbpuz
JBPaeEbP3d2Kof69EhbuBQn274Ht6CWsbBJ7JeiIUXsGSkwakCaMzd5948wBcD9aFsGnK/icaCrJ
jGgZe2d80hUYxmEYHuexlnRL7bIENaO4s8XpdYkDGuP3tAhWq4Hn1CySOyCoCtY0sg/dadvivj7F
akKEFWLpYE+q06Ic9snTtytVNs5ZxrmmQQyqXQsvWWqU9wp41jJkLdasAEc5oFovAcW/9uCJRr4x
B0OX1vgE6kLUbZ4DSiN7luwNK1tKf4nGK1S1Hu0CpwuLxVWCtOsxdU0ti0IQb8f+jbwFej9gPsAp
2rYHnYXi3250ryH3h/QMF+NvyX6pyYS15IWxtSPkCIMDKzrvMNCBN6W389ndey/yqxV0NJbtOJcG
hq/c5Wrt6Hs4a/5uziLpzAETkrFYAwgIYicCZ11uYybEoiWo15nM9A2mKMkVC1Vg3yLCYCUVGlZI
Wupxp5uUqSUJ+zoiXekfSbTIIxN8DFXsTX7cv9CTRidwdrEPVu9xkLcODJHGOX9rx+VWrSmJAs/b
jrEP5J3xSPWt/FL/buzOV5SvBXOfipMJF5Syq5dC9hYTjNaC9hPB9P6jmqDZyMPrD1m2zB19YLQz
P/aQ765gi8tMiE5GKC/LhrU3afwO8N1M0b7YXiDNQdx9vfrQ8uKyEhA+WWtyAD1eYuh9P5zykxnH
gU+AVsSkjhnE5tZDK0S+YVn+Yc8TqqgjTp1HYnoqV9MlyVJELyeEV+xWhnGAvQqTm+rIg6b6g4P2
pGZaM+Gg+YOBvfM3n357BVxKm5OWbSX/e9wK8gooI/7OU8eras68KBzuBwXC2tEhAH3egaoolDzr
S5msc8f9q8JzXnzgnjfZilCzajoR6zN+dcuCNj0cWYajEKWFFpG2sKPEayFqSvbgkDtFNQXOCIFc
Nr+J4ICqPlUoJ1WtzI/jXHkONUOgiJJnyK6y3EWzRPUSixZTqhbneqjBdVMLVbHOykuh6zVm6QpZ
ZMzNlL8244wVfbf+pQFC/pA5StO5RXP1Zy375Ve4ok91Jd2qqSyQuxsL8Bh9h2R9u5BUmXuhaYj8
Emx952ZMcOMikNbIWJ4EtkV4H4nRGzjdB5pF/ZVxYd8AIKqL7XsV4A9YE9cbUV37FVPBOBYJ10jp
BWDcTmOyb/bAwNkGPWgp2XfyNBbZ27YvC6OzIpkAp1d/wv/p9YFD+1k8sRnnEX/GGDOdnYdpTNuL
W9a+EQ1B3g5NxELRJI6GaHy5aHF7v4PdiG0XOAo/YKGgtp/Xn/yQS52gre8R5zxSspRV0x4dvtof
JuXSpbuQaQArE+EBs3/T9D4Z0cLU7JbLDxmsD4EKbNC/m5ySoAhGu/ok9+TPt3oiYFPQtA9IAqcB
FQDyWqtAK8BQxNzOUuaES2cjE+fXYPC1c8uJ+vQX7aTt4MAyYQdfr6RW/br3Rt1QV+6lcR9XPOZI
XMCI+Ynl+kvBi/gXXfE7wr5d5r2R4prbUSistK/rBKN7nc4k/Iq/XJ33N7fRvYoUUrJ4TIdEEwN3
kMg4PY2bW1+SOGsZyskvnXrPp8nWpDPzXxxjiDoYCH828PqAUO5tTPEqVVXbPap953jxDHK0AxvC
s1NUL0tTtqzGiDkWxaqKsS+m9MWSmNs/zLmbtX9ll1mfQ9zYf9x0dqwYZoiHiujWYuLX3J18F+f7
jzpUviuWTbMpru3R9JZmnoc/JSywHycIO/L3KbUMM6hznsMCODmzTATRb53qUMFZsL5Xzx3CEjt/
Yg6lL9rv5b1QCQsRdw4deCFlkqfIE7T/n9FyP5iiWGeDwnJQjAJPs96wn45rCbz7HDx7ACupMVIG
goz0e8WAL8vCO9j2npYvr1rImqHQS9I4l2ULEX3GLL2VoLtN9wCUSYNLMpE/PhBvbAO4VCNod8HT
vV7/+UE8qLxiOXC3FIO83QN1EC8cGeeK23R9g1AubEU3pZYlzYH5LLWrbgAnM83fHhyLwSCBOci9
km3cQDiJpG906dp5hMq1Bl8I7/1hjsBXVD32LSBp5YA4JO63daRW3EtoIHlV8gGUYHzA3jCmh2jd
HM0C7kPhRDhLJHmDxhcKR1PNsg0qLliy3+1TN9pD0C/niD3Bv6HqgqFJ3NY0q6Trs+VHonMQjrNA
pTxCh0I3Yp8txCAGRNJz8noUqKd2+a+S0YbfH3zSpIHKj+MiwL5RkozHF4LMGDURuqLU2iILKNHA
juR4r6wZdVPXgvZbajMSgvEoA++gWmWWyrBRsiE/UrhIEpQ1nNBbQTxHtZqnZ9wiK9RNGesJBUpP
dIRxJfrumy33M4CjFahOn11OV57HXspbZdN40D+OC4lqoPYjPmEF8Fm9FV7VHlDSn6Qj0kvUpVrn
dFQcsWcCfoxUyc1KQqXrVOTNyhK/NZlNFu4jnsWaCUXtodSNkCE8MnOtmKQpG3ZAv+Lw8SMklrxh
4vf98p9J54709MFn4t6ollm1XrPDSMEaYD40g2FdCWxB+sxlyPsqST62zo3So8YjyE6kUtbQ+WGe
nRyxV3SMmW9bwwCUQg6m1eqL3J07zlFnERGB/NdMFEP/BqB3QIuwbwwqTCDG5+bufmlFCQ35wN84
mymu5GBiFOoo9Z9YBsGvTH3FRlKujG9JH6Zln5nCdhqTmM96unyDMXE5h5FW2xMQEXF4Tp7vJE1Q
EFLxt9QMTDaAq9CGnieJusYQNny3/YmlE4w/95xLcrbVm7VlhzSEMuYlkMbROxxS1KxwIsU00Bct
yhl7EYdlElg2kl0d069BSerGeyACZsjU03VlSKNp5oIQWhzMtjr0c61RYuSkp13GvOzGmapAn4dK
8DguqMDmTl1sa4wlW8WrTbyJa8IYljNmZdH/wIG/HcvPdAQ2cW9uQ37jj/MCkBQp2Wv9gxDBa2kj
XwblEJSJcuiEJ296HFmfeLWPumzsrwJuwHDVKY/05JYm+MsrqfOOIF86pyyKP+IXxqxUzJ7bPHRT
KnQsSN5/DfPunnX8xCFEBDGC34qItyQFO5q97pv/d0W705TI+j6YnYf8DvMs6yfSfvzWRWT5Kz7P
WB2W9V9aXEoL6sVoxuNXM+N1n3vVH+rA53tSsYxzGlwYg57Eai76BjLmHoulG5sTJ0w2r8zcsZHN
lzG+3ErYTY+XD1l6wKdo/4ss4mg6s14eGL59++Lg+eW5SCNbYkxqPDffGZ1ER696QFC0BCz+MNvV
xBxrKY2RD5UXkP0Yr8iZbH7+EAjWK6SuFn16VZJvO1cm/X89kD012HhMQK3CVtb/XJINagUQt1qF
0iCqtrjnz1utu8E9q08prU37LP2rrpZNj0oynWmT2S6ZuVubxZxvgvmDNKYs3cuDOO0PHpMeygYa
HtrUz6xqLPMXGSGVivffm07VLqPPqD7ngrFFNfDh07UKAdWtpdG+jZJe4PJCy4hnTkIq/996W8DE
oFuTXRPezE3nv3ZioaGB5kN0fMgVK6r4no2nspjmJqdST0zCTKW66Q294Kse+gMc/aZNbkak4gtd
40zSJq13st3UAyL4N2Q4tZfzhogCZcI1HvKt4xm5HoWwPYUzjwaWKs9z1mSiiyfhkn0Fy1V5joy9
gXu0D9CWsk6W+q0necUY1QoBVRp6WnpkO4uSORlzl164i62JlgZongAanng6pq2mM12JuRei6cDn
Mpzr+/uuSGo6n/lHgRNIPIuTGqxpj5vKO9JlJD8Y9pu1lQ+GLLov7vJCY0DCEtk6qeSzl6eNvkFQ
udCB4nyWvp4QmMFkIex4cAo5E3dLtFbDiRxUxMbLhxpcwobf0fYxYejuXsILJk3TYtA612aDpOKq
6f/zojCqSydvMD4MbEKiF+mTuoD5/hj0M5qt5SRoQaibkJF3YQ6lIRBErd8e23os7lBuOlPhR08q
i9HADPncfYRDUSL1CAtuwBiUaANZx7EdMvbZAdzqDXY360X/UL/9oihLuJ0pnIoIZfFvi9FBHGKc
uTvbuuhpJDDSauxwc+Zsu8clqcLXNfv7CjwuAyJmcne9KGaYBAyqcbaxwEEUomNVs8pt/6ORcfIf
u2qxK8+zmtoCddY+KeYQxtLdsVC5D7yZydfBSA+9e8nacp40rtq+OjW6CiNnYbKw7NMgku43gUuc
M9Ff5sT1YMvR3qLTzowD5NgZPNy0M1xqgkdWP49cFtUNpUNmoPJaZlBtJWgKTj5ilbQ9LY5t+Tob
QOS4efyfHC0F1axBwka1wk12CnZbKo/VtGRR6CoxztOv48HFpbct8xbfccE0w4i03bFl9xEGrgbG
WAY9dY4Y7IrLR2ivOz8nvr8NduET1gxmKBMYavQ4szymQixrYnLNKV92QDhnTCva95tf4JJvwA+g
iUnKg2ScCSlPXYlnktdEK4g1LjHwdw0JBBSlzIIvP7QTYqedWB115W0krqmdKvuP+xTajwG21g53
M7DdlmlbQZ/VrOEnOmHE/9FbYaaVdgYuBYHrv3uGs4n1Mz0rUtOuSechYzzbZSEp9vnNo0q+CWrZ
kCnWee6grfehYAPFBpbYktai205vGPoDNQTfuZLJqgiErogiUVRL8AJHjTptCs6R3l2w7SoDzpdp
O6VSzan2IWvHk0xXtPwKTuALyzJ0ZLiOzo+jnxaGRdsbYq0GPd19dIG0niiTaE3yIT0DAASOntGc
WTExQLT/QIJ+zH8eFGlKsAiWSAtQ9Yb9zMb3Xw7jpWYyOo5ZHpjLmEPoa8nnnOYEPaJv8+IC1/I/
CCXh8CjYaDx1Osl+I1Y8iTCR6noGkZt1ALxB8v5cNlU21ehDO3sj/WyfPNMvn7g1/PemqbCwsHdm
T5NumUjbGvdtZ8I1G7/nTbep6BFLm9updtcnzchUMOtx5S1Bnf8752Z0tcyGbCYiKv6Qv3dS9imT
gIkGXiqkirP2Zbw6QEQcE0dy90xBIwnJUNy9s4WI2yJlzyDGmFbMLelTpQON0Ev1bmfw+Ebboxa0
//ZeajQe+O1s/wMpSFy1JUz81/J9FH5117W+GRqeEmQF80qbzTQ6MQVjrsM8xQtxLBEEx3tveAfQ
FK5SD0nxvHrn2deI3FXOHzVmMi5tLUi+RVvsWhqTsIWrBclm55jQMqjwveL4ZmA50aljdvDbUe8s
hwvE3f4UiMsD+41SZoVI4JQ6xSKYB3yTci+KZ2Q/Y4vEOnO8zD2oask8mSd9Ug2LMdVQxneo/ove
46C1DnpiDYjqEXU1j5/ISX/WgcJ0b8H9k5paAwAGNBgIhMOOBnbJtA1nd+LcsR8+dpEGWKBlgtNb
WMd6MXNjgOe9DVieRQkTzZuhs/coS6BVGQg+GUWu0pJeGzkrbJ+HVjh2bBnPYetASQ44h8yTzW+s
jCBWQ0yz5UmtXg5EFnemsWmIc563VXgbd46vf1RUIlwZMNkJSlNkRWrfzdW3awxiMldLm266eVAO
E1JTcKQcUIpUU5zdg77aFudP1ICDUQcGFIVB2uJ+6z/0pK3OgW31pRFOUrBXdw9wGglVYxV1JHLd
wQaEyAm4+nD/Vlu4Ku9Vr1IHpJA+OdFHEJBP6+yTv5RoUvG30h+g4mSpLIR1zoZqvFAaUTra3B64
SFElM7ELHQfFufF9x+4uertfequQvIm0aXwjbtu6Ged5Y3jHpbShsRFHH0ORmHF36J7XheKUlP7P
LioEesOh5oc69rDEMcYlJrjOStANMMGHXtLI6r2Bj3ePYDJDcHRbb6J+jTk5wo3SN8M5KNYJ6iUh
sDMgaIqzVh1ZVF5lpgxZfQIanX05Jd6eyJWA2d5ysb0Z/wreO0XT5V1njxN+4dHc7/Oqi6qZeLcT
sUrOIomWvpa/R1Eg38Md0GNQMzzDjmK3nlefe+5/Umdb8tv+RCWj7hb7yk7Yi7yEh07vioGvkTQs
uj/BCHeOhmQseR92dd4QJd+iRNWRfi+pjbDKBVbB8xenovzS94dXhPHha04te7jGix76DRxhylnt
xq1Dzhl3QL4bAKs+dXvYNHctMZo8ALz7HTRuL0FNbOnjjlq3LWW8S8ctacd+sKC6k9FR33blUIE4
GplhlL+1QGg/OyBnv2b50rBo1hOwhB5WJ1M0NOXFi2VoYfA81z6BF8gqVXSONt+HJzT+R3lF5AUy
xGDK8Y6DPCMKs4mKx86BurHX0iFjic5t68aW8wx3zmtwh88WBtFMgVTVEvA59GB/mjU9DShRbkBL
1/ACov95lRqh518ABER5ZsNipk+chtgOVa/M/JqhWsRhJsP3YFWoEDdHT3K5auYH92v+ayFBsYXw
2H7v1aNVlzuwvV+XCQ5cbeN20tIA8kN2GqYk4/+A6wVKRy1332B7eQijCfSXwf3z5SqoIamkkxpD
JtkM4CnqEdkxmknzltVxju8W+X4hDH+pGsaRTqdqggiA3NoKQkkbPLvR5i+eqC8dGWLbxq+xzGa+
XwJhGHxdj4DAPH2ambU6oRTJEQgZnfuA3sPoYFbOOVL/9ER6kGJFSPbCYvAbML12BsYwJLWIgk2s
6fnL0n2SKmB2uxNRYOf4iXWlvLlAfbGwdIFnLTG9hC1CbhKIQoqX4V2QRIp7sNFyoq1aMJ73EP+p
ySgSm7AqaPdG0+ssfbB5yque3hLZyhRAjPpnFr+ru0+TiTMUDbbbeXXyzNlYHsG1AWGUgggleQTH
QVIAR2jAYwOh98JwNmyhGdKStY/ckQEJ5kzaxZHShhXNmHH7C4KQoVONZGG7H3IHYpRHxCph5a/y
wDMSc7khxxu5Vr0mkeH8pvgopqamq+nvTk8z7dsYrNUkDGrbTeiWCKZIgubkVSBfciNEFS4HqHPm
dLvVB9+D+lERCmu4cshYTPOyLkoGSEzttjqDrIzsTUYxhD8+cjOhkap5QGJCs6bNk1/bqsBcsTvn
c71UUXb2ZvjE7ptAl93zICiATsz6zRlsC0yMV/pG9YepR2rMQ/jimvWDEx+hczD8f7TBOD2mnCPZ
iSVgvjdTVlPfFFh0gzmWRb5bqCltw0kfGS0hzsCppe4lyFrKTg5cDSjt0S5R0I9WEqtk58Va7pj7
+s3DC+5gIdfpFKnitqMPgWzJhmU4jCnnKpk6glPOTR/OI0SoqUseBqGvsMTO+nbkZXR7BStCi/tC
Mb8V5arFaw/UgJSTUCiclw6n/KvNfLtmcNx8oFYIAiRjo6dNRyGczGHgx78g6lXlMXxzMWj9ORyw
eqCeFPkwZvv1nQt2NYGKn6vV9bJ6OeDCoIAac5de9G7yW70vLb57iJDy/5hA0fep5Zgb2xAbNqe6
T14iKXrE8jwrShjSL80qEC14a1aRdLwHajrK9d7RcEGVP2iRDCAqAqQAF+GpNfyAvAs0oxL0a7S3
BsFp3ixMPQpDfeZm9iJ/+2LNsgIadCnRvgyXATWoVrWo8ywQYsZukaglB3ujhw8s1/Q7Yv3/8zFH
ue7X76SfCtbpwW3b9S3hShMASGfvPxch2qFiA41cXTMeDW1fOp13IXfRCqtrqOsjutdIPpTpuYV1
7YimkUxaFNegOSORrXu85oHRn/sW6WAtNp1L1hD2JWy5O9t/cdvqlVXKvlVw4ImtqzC8XFMWvwH9
2aSAJiQJSQMtiSO7//BGyeBoEk49jOHeesghBaUhc7QHIjKKiPgGMgpAJ87zb3ly7op+wHf4twpC
1lsZY4QbFWaPTxhJfUm7aiBTutq1JZ6rClVd5Wh+fzpEb5SCUtbsl6dR/vJ8VaeGq5jUjmeirCrx
ERDCtBelZoYusjJoxXEn6g1cE2Syrv/b047slntv3WPAa57cQvdUt6nJ/FaH47bL2pdKC8CzSRYs
4DdyMsL1mkSwL5cyXYkF8K5cE/gWhEXKRU4ouB5ToPR4ZJ0JtpcaRh+rgbY63vBGoF6p+bzHXM22
iVsuKx6CeZY0b9A/BMCSTcYZDJaIXJ9tn9Bm7oDaOIPPhhxJGqfXlyMqpv6/fvbZ0UW2NlsGxCVO
HCO2VSZuxUNAE9nHXyQRvwhU4pTf6Qv9XC8UfQLCMoSjaadVCPxI6aE2UmTSZjeEDBFWBaHe4ErO
+XhbGingyPNT7/nORFk5XxDpxLLwNT6q8yY/z1ey0hrixBzobiUgAj1S8ZAMwV5OVbDk+beTV5iT
yCZiwfF0VQr/fcNJ/X04y1LANhJmkHyILyVCBfCZAQlZJN8AGZJ6HkXZX9yjDIden8j2bBgJKV9y
APugATgcvc5QH9PjJJ/Oaziznx3U6IMuhzRwUzpl6LS4P3Eqmomqe9MTiAQ3bRLXka1iEmCzfze2
DscENHMPi8tTsk5BtJhJ0VEN3O5nI3w6I/ATsSM3/9PPeC3f5XZKL3DPk4xRZJ5h8K+4Z/wXva6G
E5ggxW8988e+zsbAVrSQnMH7mdfcLqedh2YNTXonjOQl/EG4Ch6/KmX32Zc+loGwP556xRUrN3sv
5cbxHBAvw0J2z5zgh4uIHJyCPlXkvUIotQTExhkcEyQiBdLGRNmnx2XCTu1ZG13h/V+p+gyBl84F
FjCg0B/xUGIVbsBzNzR/QXbDuBchd1fCFpYTYWHiRU5FD1XJD4W9Yu3+6O0W/iVdQAIBQlX/5vVb
Ov40qf4YSqhsAHsp4R0zIlADsJRr4cdFfihsw4icp2wUIuyJXAwF4DpcKGH/2/NUKUOvC3DRga1H
0NO9oPYz3qZJzZQ9YgU5IhNVNmvSsVdubv2Ybtb8hySn9GFkRmUOWN8uHfQkW+uQ6i7+R8JbgWBS
jy4XNQ2c4sUhLW2/CwHSPoewo/jDiIaIIl5FHMyD66w5X/DEilZYPPY+35MvRxlhaz7srJL5s9fO
f8cbRSlkLsai7BeapfRqyOXyCOBWY+cqsQbPDWA+li4SCSvSLA6UBCYYI16fVqlzyEIXqBvJoCqm
xtg5q9uHSk+eQSTln+73cTlCADdCOJUKXQ6TiIXD3hJNSqeVZ+M6/XIkJGQzsyNT2FDa6YMj+d2c
0NgChacAaXhdzJsz+0jLVNEV7P1QqdYlpd4LxZ9A3pkYOXyyppjRlRkDRcsdk3LZ2dcWvRjV1YWK
9RjQB15tOo3fh8RfyoHuwlxKnEEBo1Zy/y7GSz/Bjik1av6r/k7jmnVC9hAVxmeZrxJmqHmEkiDK
LjsEaJwBreBzrOywHlIjUAlfLplWyvJnTCZcrt4lTyzxlhITx0hHfVVmrxfjzfLx2vpZpikUIAQX
yrtnov0pyWPpmjAhbYQVFdMw+EYrZo5NpeM1g888JZ1cqmzkuyFmRYb4jEQfOtJBWUUoBeFMXWC0
99hytP95Y8xrqc15gdQwUjbZVU6FI2bNKOti2YioZiHpBhgHRqiwIc3uYXB2pK0hIdRroTN3oPTG
BBoNCfTtliiA7DQKHIGuaMUuq9tj9o7sW5lGeXzVDKxfa5zYfO0KT3W+yv5d0x+y/yaBRN1vNbQ3
KULUl2PfVusweKVxXYuui+E2J6GJyQ/qNghtCK8GufdR4xCER+k6xU1jZAS2OOQat2UJ43TNlVv8
RXh8SZbYW0yMSKPmssb3m+NOz/LF//5Ep6EvFqcbFbMrRWVi9TaUECqUG0kA2W/vOyy2d/rJEUjR
/Q7RBPtP2endBRf1Z9LYg0CgfuBHeP8er1APqxKUr4cBWWKJzBA/AJbo/U/RgymqDXbuSRi8azEO
BdOQfb9BDHKoXiTprU2JgpKeN4oxUIWZRVU58adIkz9Rt6IN61ufdOwpsZtb1a08aSYUcqNUveQM
7TDEMHQCdCYSXiroUb9FK6iU3+xbDKhuzfY60npfErNROWY6r+fSUbU/eUmkAczGIHzqq1VOwPDK
IIEuYF6a4hJ1fay0FV9U+ztvEuOwlV0NaVsezotXP5D8N31iannwfUcfqNrJNSunf5tqDCT7imiB
QTHTsZPSL6beMfJAi6fAMMYe3h0zEMZJHI5iSZ+WSgGvztJrqL0dqP6ANQB+2cXNbH1QNvwVHF3N
u/DwAJbIlA8EqEKS3cc+JSaaLTxDFeZEQHMnRxJaKyeWCv0gY2MwkMgaemrBFkU+zNTkRgzJRDMI
nPF55QqSKLwSrRIabLISVRLk/iLcOlFvwkRrzks6j5TRQHCZ/xsZ4VGo5lL9Yt9K0dzyZqjMj/aS
XY9t4A5r5E/EhEPOQpJvgfG3gx18SxOxsZAojPAnDilnrfHMa8YJc/B01l027SUeVPA9gKITAKm9
WcnRwXXUCRV/9fu/56HHzt3CgrtPF5JgUwgDnWese1YHk60SMhisZnr7XeDOb8LWczvYV1HfWCMS
xfWK6cCPrWeP5IAgv38yFUQc5LGibzn+vxlQpdzP/LSKyQFR5LoGnyoV9ORlY+m+zHINo9WaOC7y
2K8thIhPJDra7M20Mhxa16SG3KF2/k/SFmNemaS22yEPgiQqxTVnt25a4rKH/NMB9x4XiHOeSiet
HcUmPt5o9WXNs1kJng7ZX8depEGA0NCeamKslHSGgmZvbr5zd6RDSbPXxuXueZuRdYYirq48Lnxo
tXFClM5+npDpgEPfq8ulUiZp9/coPHYA2/920HQJg0u0bUv6S3IQ1kjFywdhF1ISRfjVo1Ala9i+
iWlAzTVVfeUTrc6xTmTsX6e29dGuDAVKa/k6cAUlDGwfREDA3dkdj3eufsY5qquNm9igFM3z8oFx
glCIn2uIfRQcCiFTjmtDBoUgjGxkqPkl65vViDsjEQajNVvfHbTlSSt/FS5/xIqp346/HJKY2JIR
P5X4Om69wCVXYaUJpGdrhvVM4nEdBgXjHATZzpbZ9xTWtcaLktWSYqkOuiLJ6UpQgQ3b6Y9s40oO
zzVHLFH5nWnYegL8o12jjkzxq8/Bj75HGg23u1SA7wCudpG4l7iFFnXYui/UsFAUGU8L9pwFkhZ9
D5ZuO0iqXmnJ3nqvMPUDzLCIQcpiJaQ8bKPzIFQeA8E0kBB+pJAks6KB/TdDnzQpfKutbg78t4FR
Npr29R65TTtZ+eocTEcVaFbnIR+BNN4RUK1S+nQ7wJoFLgdd3qyRDk5xLXVv5ijtLpi0iuFQCW1H
gdxBbZSh5fhUNnix62OLpO6l7uzSG9c+JVKirZwOowLIqtYn3ynB75Rmp3hP357GhILzP5oHv8Eu
wLQzGbd+nezORfapz95Hs+VNRKZNYe6d3C25tSZj1PWFEtrHIRBm7xMRMlUtJKyGRsYCXNcZEzhY
hoFLGQG2pPrFO473qj29AL3c86L+lx2SJue9tgHw9emYPZPw7kL7IuTcL2f74q0HdOXX8Ig+FpSo
6XXOyl0r+MX5Py/zZfGOSezh8/r9SPyu7dFqJPyS2ypqh85QHe1GDLIk95qdmcL1TjnzxZPLwwD1
HWbI3QR6ZW82wXpH8reeFI5+cGYqPxmUewE7rb9xP4hnqtcUN9EaNhzjhwWQyYw+b9WLh477vfQ5
gyN0gh/QzN/HxZ/lrn8JqSzPuTK2tWcOKBIDEkk1UqsRZxTa/QzjAuxYEVsWLWHHRTsjJ0g4mwZo
ZjQhceJZgE6pBD3vtuuvmL/ECG0ZwwjBUQ2XDkNRv3fT6LIJJK0H6QFZOKs3X7YkkKJ5YXmHf8mw
VvQoeniFv+RmuDgQ8Q16QOn76VfOhnSmLaOWENjRYy0jElF8Epe1Ip0agaflxupF5hKGMseICwtd
R8MX6e/ZDVLzpn/n/AXjushIJxdsA3um65bnW/rjQiKbgPucdL50+OsjgLv/3fpsRFnVTGy8EBbp
FApYbSY2wfJ+FbToFDEH60GmB0IqKvVmfyFmFEOS37hf20zhqFSfdwoW8cDhk/rU2Gs5Be4akQd2
goXx4zgXWSPXUYb+kYu6fh8xnutpVR2qk9m9pVS0jemopsRled6IJ5Qzrkk2LqtbrngZ21MwKROK
p1orhc5D0ZnhUO+HXCmcnp7JtnHhhvhbuzoy9BOas+zztW7HK27mH+U2zw1hdgKUJrD2Ux1QfcmS
OtzCfNI+j80/00cjMyhSQr+db6xeW9OYgwY1r8yuPNjHIpOt0K++HkanWgOch7Pp9WXXYzTU0T/W
ROg6j0zT5GwU7BusZrRR1gn3vlQz5H+bkMr7WclMwdxwwwAVJUKC/xfTVjgjUZD0SdR6dLFkXX1j
CyYHT1IJE+KjTaBAzup+p4YPssGBJIJ0VAwPQTGM/BrHGHk2xsr6GVuFBJAKa6MIUWMzvmfe3L7Y
NIUMrFyprU8OdzTD+v1GOGvoadjH5xyUWQSJwzC7d1FTGFdBOcswj+9ozGb0eRd1MOmwJQYPgvEK
CyvJbUzSlNl2IkJPp4gV1QrSSn1KhVbTjcPJkUxZk574LdU45DUk+lDcztTJvBAw8Nfg6edjbL9F
+4sbxuvfomkbqrhrEb9tYcj0aU7k0F/jS3/rSlzA4/Tjo7h6hHXJLJdGwRFs8Z00VuE7zCVckmLT
a6oEkTNvRYGl9i7orCXZ7INLmUW6fPnXfc6Wnd5GZtWFR5iE06B1JA0jL1WDkTHnMrBbkJwN2dk3
rEPnrOFy1eUa0wW0+mwM+6KGeZEsDR2h+GJjT78GW3eSppITPhZjWztrJcyttabEjROexVvN0JHn
pNWQ5fKUNiY6veXJZyBxcP3NkJuUpjDWLyogK7VZhqtuEm4rdg9ay/3zEIL62Nsd1eL9IFtmVnkL
cXTBzevgSd528xNmRue9IJEjCKoAlhdX3iw7dOTVE14yiERedsPksgwSuE+WNLvxbGt8nu6qXOox
GRMrRO3nBPxu/4TF5x/obvyaR5iw+1qgNFNdnGnJ3raP2UJbZLst2BC2o0UZCMGO8OOdvJMCQS6u
ESKJWDKvB94CR7AgRbRrZNOzr+RcHBUvlOfw6dX1+G4o8EyPqTh3KaaOwgwGmMmjK5/3ez0fXzRE
JQzkOUA4+v+3WUEg69QRSFzkJLx4/+hsAOlH+31Hwy/77vuXvClFrgFGnMQ4xvkM66WQzGAFRzk0
f1DfkLkFIqLb1Ck0K73LQNKH0nYD5jELIcq04nOTMfzmPZTbImPaGy/eNSCizdd3uKE/jFc/fyUf
QBTjW1sEdsO3P08cffRH8TIhNjzIRZZvu0OIBQlwJTI+taWhJEgNpSzshslQ5aeROHpbPHAZ38sL
rfXdr6vUxjnVJmuvi8tnh+W8gkzX2jVh+HoaSpEOU5mrkSp1FWmBuy+hfYfP9uCxOFnzgAqKUTyt
gBqJc8Qa85S3i4tFF2tftzgjHzC1dh9tsxmWsda+o9EUSUEg6NNKqymqRAj9PA8FNtPjiEWE3uTM
IWwEQgprU7umbhjv8s7p1VT5845kFyPS8Ozl+BgJuKVMgJoYQ8Eh7nBScyaWniid5mFrUErxFrnz
HtdbQz9Qj4v7u7IBMdgvQh7avLyOlt8MdISJIQfVOMwz8BmFjVjCDH8TwNzLp3DBUpDAVbL54Qv9
/WdjI72gTXB+DIo1/jwxGnf7YX8I0ykJfP3RhW0axfx9XfFsKLU8kx3Pxla4/RaTHlhYbzo80xlW
Ff3xYv4Jmq6u7yqXeSQS55GOzx2E+9+Tqf4lOQDGgGrfJaHC++1xUecGQJo7Hsl9WCunb466WoUb
5EdzdvY3K608OAACunxb5CEuQhe6sITYRYo79GN29F01ybretcN877C+lyKZRGnjfeIPR/JZ0RiF
51nJDqJJ7dP7v0mrsBIASFIPEMpzOVcXGLXOSQZnCkKBTXdjCdx1T9bcUvL4849dacfxWDeo20ls
M/3TPcBGw7lGMrDwUhvEeJhApyJCrknOuSs3lie2L3cMUiA7hHLnOkPyVD4PtfGAa9/4GuhsldpE
egAOHEdJ8Wdm/U/x1ozvfwYTKZXUFz+Aew8A+C29dJfkCbYWLZLYErAfcPVq8FmHjiEwMoTH4iH8
yn0fWH3KAB0y6p14qCbSJ+8Ew3q/+f3Iem8n3Ive6hKQLhqnmWlsKyEXOqAVD6gnfg/n3fwFAcgx
/sCzXAqud8RqLoOxGo0jjXaVivaVyjMw0hWakFW58FTcbvhhPY6Gc/lsn8xw0P733wCdYBBJ8GB5
UScoibUmidWda2Fl7Wu0KxrHSwYKQuW9RwGwGBMZYPBBQcTEKOaoOsBD1k+nD+9hK8Gb6eAW/F9G
cguWXk0tF1bw1KMGcgYqqnLKZveVUxRM+zFu3VWweP2EgWUGGwUECa0HMXhhj18O6pK0nvaVbiRS
ziC0bqFi0kjok+SV2IPyrmah4UNRyaOATN/PNm0St9D93KISLs/uK5UYRzJPCRuS6HOkeeLOwoYY
zPHmPE/k1BDpkE44nqW3dCij0asiMGDAQP0vZOHBq6wIA9c/J9cxuePjuF5vgVHiz1wxCoG9GvRS
CvZvEimrfMJbpjg6VKbqss2A9dVBTkI+h+1YYxcyqgzfJCrP65n6uSiirllUBcfPBBz5QPcGiKFC
cccl7IaCebfQ8PqwiPGgpkv27Jf1gRD12AtZSCCEgOrNzAMeBq8bpwV3adw9SkQNo8nBsdLsQwOj
vaQOvMw1OnpPW4FBwueN/hHNCs0PLpymb5xakY6j5pjhMrOKOuilu7pMBsanhfOxow0sqcsUQpFH
LZqSUzkd9fakorYv40hfKw1a/eLYxSgLLULcUuSKM6EpDF0k6HjGExiOOqi2hieep76NH7yPFxGi
uVbzonXgzYJs+RD7kBK/iUbQ3TeofW1O2+SKugCOMV8TCG/YChy5VSKdIf9NYp7IZ1e1DDHffKHf
JPPukDCl3hE86NVGTI/xnz05k0RYDqSd5ZVT7qOMBkqQfUDJeJ8z//a4MVnEtud7F9zZgSa3GO7o
AJ/BbJtSDgYD+rTXVLJIpZ7WPYVInnsq+L0t8ZfCEXTUpK1VfLbIqjklhRFqV32cT62Zs0uUBVOg
cf/E2BpaNormlNWrcDfTW0AVY0vs7UPP0zLVJO0b3qhRzlIen7LOH02+ktosHQXcotvWAmBwE8JC
M2xWsz97XxANn6h0hZSHnE0dmqxFpOd/W8ziMd1bJS92vrgTn8ZaRyhw2OoumnxDQ7OrHo4Jpi15
9TjcUkXdoYlbjA/EbIw2UyhL/mwt6Yoj+LGk4qoJHJBpS77WGDdwMkQXB4VrGE2TuSTV6pHzZiZo
MvJSia8kq4wUaRqfT1BfmGHVrxbLTzyPBL4JWlroWTUMlWCAr5+/plfcB/iDjjG6rXVv+x5zDSmZ
yVxRRJQF/irWu0sYOnYxQnkZmTmJZPjj79+jZC5nMGtUYVjYisggp9C8qLlqPyVo7LX1I9q0ZTUv
tpHQfK4vC1D2L6h6H0WUSBa7VAG9W/6SyokSNTJe7HdrP4QOL2aIAFVgoAjnANe9JEH4FCFtJksM
AMBR1iUim6iboHVTUkm9UTf7bQsOTjkZ22TcOnjAEKhmWnn6uuGiuXFJ3/jKG1XDM1AALxs0mN2P
O+BitGcrsIdYEW6TaWWHwWDZqlepnFVNLqHrksL9tvpaDulsA4rqbse8eYqpI/zqxXrApuWkIRri
S91JlmNZxwwgH79XKoG1xkOJRGUG7WkBswSCNmR+/M+MMwyp8Dxnnkp5g16CqM1C2RIAk+LRIYcG
UjN4Pt9qDLuNQgYFgg43E3TZMGbFiXQXf7l4lTg1iOLnyhUHbKUOHtfoAo1VrFpT7z5TFIE6QR/e
kBMD3mCpbCH9hzXXK57NqRzsdh9cFRnWUgD6oG174fzHnmzfBe+H+Y+c7eYUnjxeY6GBQef+SQ3i
/phigeQhKV69g03fkkGcoD20T8k71TeHnKApv8yjz73RpDvPFKpvMfqawmf/6IFpGcTf25Dny7UG
nvYsV0PqPpLdG421ED3Wb6DIhvZ2L7kr0838Q+ZL70PAK3a4/W/fD+iVqGxQv+L4GlttuX0846co
tkj6Oxxe0Pw3XWpQ1Bciids8It46QhYGPIUdoGxP/1oIQUB1ZcVvxIi4rL+B/nYIPOqpuXY7ubjo
+YixFFoc5rzh3vKJJsAk7z7ksFVXrRXXoWs9+l4JlGZ189DmulJoZxlQ+IdiTUbnKC/C2KbKeGUS
NpG/rs/3t8ce8/x6afVtVQSKi26XsR6p/BhjmC9KY3TO/TBdu4+qSNcYRTp7Ne+4HkjpFBVagbII
AEkCi545aKBw2pxVwG8J6v3FT1XtFWyopjXuln/Bq+nPTWblonNie5Y4yN9YWdIQTj7G9/N3B1lV
NXVZq1V5VVdpoho2YfArieujUZggJcjaq208mvojgOm3wEv2jmZnsr55fT+sSGqrzVY0ni4XIJ90
/+2aDzMmK1NcB71aeUmODD8XvZPR5BzUt3HAQy12V1SfZSVouQsjRgYUjLGAKB9oudclDfwF6k7O
IWAuWm/Be7e1iZffdpQnbYA2iN+Ootw+QGXaeI2U9JKoVVmbDczhYOvbTscF0K73bINKOlNxIfaP
5V43fe2Wm7Kmr8XKXFQpFvcvWRs9YQ7B7ppdrKd/fAFcmwYVAdGTiUByTj9DePijSUeOUGmAn7ot
KCy8VqhtP0CvqzsvMh0GZBryLA/1Q3wPFzDPzgEqt5pX2h/FA86ErF3fiMI09zTKuhLSaI/UNBzr
TFz9hK8pRm8JBq1pXbl9N+OvhnlNZhV9ReLzXK9l47QRAD5Za/m3Nq74P+a5V0HvfIkvWUBTXdQm
QXo4bkaXo9GXZjHCDQeFSsw6lCVty7/HtoCXI/c6fuTMmvrUsbEN+X2YCQcnyaiSCOBxuPI8IIvq
4wYPGSPkpvGSaihO0kscwh+0Qd0M00B+1sh5F0Ex+fgR7AG1Choqs8y4HIG+Vs5+6ib4fovA+Tdp
PTbZa+Trl+oZNR8s5wrwokRR/bN+q22jCbbFhNxSpx1LNXQkV4RK36O5vrr0g0KZbG4oMefJ4j9p
/xnnJ27PhK4W8NZ8hYn97Qg+NrdJr2ZydCypR9k9l1OmK924T53NiUz9fiHgXXOt7enYp7dN+rUO
sXPIV6bqN+eO6TU5kF9/pivjfkkFVdsIV5HRd26NrAZrUCWcZXAfbEMM6H4cuwIk8nQEWIMHtjbo
g05uDfZ9wAtSvP8mxDbPXOxGaKHuelikikdcCGtT0EcxIPkArox7WC505bon2ThjcR43RKCCXSSZ
yGEZJrNrTjDtoiRSNbudTrWQGrXb494wX6gYmXYaUmMrDPNOraGpllgNmxUUX7TlhcyfP+pYwEIT
nN563mIxazlu9LPjF05xHsnYNZTSC+YAp7bpTMG8U6xCDZu+hE7ZX2jJyiggDjyRdyzs0prfRFj2
BM5GV5OCua0cX6F9a2Inm8GCuLRo4/YIAR4Lej6QTVa0hs3HplYZeVNf2OSIuE6aG0lZoGvSOx64
C3BZu5mrFigX2IGh3mCqsmDvFhRBzVC8Cjp9CuuX5ox76l82dtMre+pz8MtcvfSLtpgpM3Qoaco/
NEbpvEdnpH6cHQzOsz2HVZoIaL3AVutOr+kcEC1uF0m/bzp37C/0hIVUxwApwIv1ilW/WI1D9OHI
KWOZP7TziFz4J3Enfqnhcwp3nLGv8a9y+MI7wUvIVzmZpkSz+A4z3/ZTx7vkCdiu+Nf7J/LGvFxU
QHIIpfGoXdm0X7H8rrTVKItYBTcHU6s7/SK8T4EZGsCvvtoCzIP7XaWyiK+y6Wx8vDHefUjtpE20
eL8UQZaR3q5oovjZ+WVi1PFYlmbzB2qMI+dMhAOHWMms2YG94g/X6Fo6kyPNZf69koBf15oLXaIU
CeC6LWQqEeSDEZxH3PnBhjyEow1RxBUK12/fMr3jPMmuo4LiEDXLH9vO6pM87MrTS+bBuuGt9RdN
tlxSD18zPtaMixVzhDlzKV4OZVhSL/6nS3AUD5XLPdEs04eTfYYTyy+oWrNSD90qbU4lgVzl6IXX
zoSSlQCEi6ICuee1VD/fzL+EF9Lyl3bfU7+n1kvX9KmJ0zVJ2X2iny9/hSkeQhGW/u4kmmu6w1mY
qOjlpgGWRMWiPqVs9U6fhBQC1Px746OgSnxg71yZD18PBiKRU3dCLLh3xjQM2Pj0ggCvhDP2T1I3
tT4WkrNMZD7WGGrClGxSjr9t49Y7MwN0eWjQY2rIgoXZSFr/gB1IAg5Rnx7HNA0/AMwqUxbsFzWz
LpNL6C+NHOFmpgepXlARMAE3EfOcUeN8+TrgY4T7s8u4dY8NRM7vMMS3VKFOEq5NeZzOmG+Ba/fC
ttzzoR5vVY4bd+9OTWUyYDZ54ULWt/lZsCGvqBSBRkkHEXT59j7ysxVFzlXCXMcU7gT2yYeA7xWj
Mp4QQZzgH5s21Rqdd1u7WWIkqJH0nhf1t0nJ/S+CeEGjKbtydL7DlFMJMpwcW1e6eWP1Zhh/wLF1
rzGcu0xtkfdQNaPrd0yRPBVWl4okCLDPUN30/Xwlh6AaGvds7qKsULPPnoBOa0nHd8itgCqsKOcq
fc0zwMo5ViHzcJ1IB9AP0SUkr7ry4P9S9UH5/N6N2fisRZlwnI64Xbi6egdjETbUxsusEtYgJ/g/
CFNfwzG0qU1jTLpBvxwQGsy3Ubzej4GbQNiVE7Zmb13og5lFuagTABPH6ikrNoxpYGnbLzR4eMGY
fJx97Tv5n2yi92MsA49VTDdTkZvrFfVbsVhD57ZSqjsfWbCj2JLK66NXx9hMA4ifVCTwQxjfNZhu
q2vc7JmKAt1fKfxdY1dlnxuvXlP/uiKs2oPB4cdXx1s00uz/zlGqDaAvknYalowzCPf9DRPOczRN
/dOnQF4CCLPdhhW8QV95RRRdbkJWWCVfKT+Yims1FXjVxB1jWemuxPuxgcuVwyRkV7mJZqzsO79e
yGdydlj5uA8rCtLHIiXjnudCyzaCf+xz/nqlJbRSJ0Wwn5heBVoEP/pJvqeGYOh7l6Se6g8OZSHT
3GdnyIp8Y1Vqv48hzmLK6t6/R28YJrg84zvbWGhy5WdmQ0sYg04S34O/jfRLc0DLsUU0faQBEkre
DTBYYwSIAH2F5J9habttq5w/kE4t7mem6PqfJ8ZCpKQYvUj9EewQoron86RwWUqFGxQkkLWz+Pd6
BrtzyVKw1tueaNjORgKcJyOA6ErL+3btNYyOAK2RH6qcQmb1q1jYYW4ERNJ70NROm33jK1AyMh0h
DM/KJhps6p90KzJmrGxxqM91DHeusq0cUugkeqkl0OJEr/Zcj4tixEOOSPYzLfw5J4QiIR2kKN1k
wp1vZEMSrUQZd6C9RY738GZWWVa01ra+6hxcRaA5wVAt+24lM6FwD18AlcIvcjX3wfNHUjj2OA53
NU/v3+c08w0E9+JglxCSgrnKQyNMdnqq9rmpN4JpV0S6gntjYFZUDAJv959cVmqClcIYsJ/ETKt4
PNA8dQoT9Covfu47oM+RIMhWRrcZn2FUkjUeWz1YAqRUf8MShdwjlY2eJJe5lhjkEWzVLgTH3+GR
B6yG0jAFWc2Jab4LZ6Syh8BsuIGUjc376iOYLS5F/wfqEKJCF8e6CSfJddHRO6Wo2vA5Nq6sQYsz
FjLAK9tBnaGHbMhKBXEuEQ7w9uWA0VxfRmQCCuoj0NhDRvJBqvu0kpbhJZ0ahkJrkOCnRkvCyhlm
33uzrv0KlsAyoacVZlN3bJfjFT4EL68Hr7gd14yUHuCllB45RUaudG/aTCCNcsUAK8S8p0Uf6gl+
09g2/k5uCM9ym23owSg75MchUZQDkjMK9iA2l0heaAiR4/3sXxvpr77lsTMZFd7l3rGIdDxYPzec
x83zDRC1j/cFBKNvxzdMMFhVSkGlQYFCL8VFb7vggl9nx9kVkAXx5gmXze631H6n+XgVm2Gg8fN6
npNvuI3eHrTCh8DMWyvnRabEjTVhCR3gdo7keM145maRv+3EPFbL5bXyCIJl8XGq66KQkD7TUr3a
/PGZS2zg3eGCtysDip0UGc5SB4CxcJI3TMw68eRn3VquasyZ2Lp7Slx3MMQveNuhn6gddT9HJGh8
krfJkKej7KzW+J25tSHLUGO3+PFcrSvxVi7blbHS4BujvdrxHp4HAWGlmcLh1x4IXuhcL2ksET5N
KYpiL8/iklZx/VYEJbRGyqIspISrYn2GjM/XA9i6+2tkBHaIr7sTMWi8Klh4a38FYDhXtQH3dty5
dnl/PTMkN06x/Jyle4cnIY0QsEOYwJ/MIHQ3xHJs4s5MtulzRKdTzgHkwFpVqr2Xx6rnKDhHlngb
5HnLq2M01coh5Bg9uujDMb7G8eD6XhUqegmrB/YIn7cZjjt90H7CCL9gO4xCgB7MYYElTdhquBSM
NAK6InlgfjdwZRjOKeGM++vMQ2KjM+k2Z1bJS4lXnnu1cugb1wSKEwPW05Yv0euWp0GSG9cNnfOV
lo2KkENIRmGzZdFJUI9i1wmu54/9iT2Xabj5GcvxS/xqZtfvRIc5l+XFwDzaSBXl29bjDf6emXai
1ATc6HcfCfZzErM5C/YOs1nrpcVgXAdGfY9cvSh6MO3YUF1Rl4X7z5VRBL22LNgf0IoVpKoeIG6m
nKi6JrrA59xz0uTyCQCcj7nySxNL0GziVx4T/XtJ4VK9mU+PtU3gYsyG81RlE1dOItWFKu3RwcwV
vNXqrOldELQJ5hP6PVzcTV1P0x5PQ3li7tzmFKJOc+jQLnnK0zuZ8l924P6hSSnrqxfZZC5kvPlw
+UHXnaXr4BPu5jutK0nhdAVEslY6tz1qWu+RqL13TEbnI8oEWhlwAkiwGLZ+ad/eMU2bebbnxyuN
Yv4AZh91u8F8bYVklT/qqp+lXfdGzuA/5M9ZBe7BoPyc+0UsbQikW6x7eqdDEIkym1BIEbh7bvY0
xeh+qVobTqLU+kNNug4yXl28RwYRbJgxUzEVZri13VIJ9fsjzr8K/w9cfvgUUs3B1suihj64kTDb
dxfKIKWK3bZv12fTrsKEddIOuzOJ8JMSjNgEaZzIsQpGsICy5vIr/WfkyMJE2vCwE75PGOGHjB8a
ZAuAj4xN/YigMBVXcr/izL9flIk/Ss5VqNtyR8lekvawEHYRc+DAn3BvoVN43/XtKrOUewv48Vdk
ncTA2xcamLtxyXem9Gxt5dLfhRqck43x1WIlLQEwXxMbpQkQhb00wuEUiWk8Uz/s302exLkvP5d8
+gzliy8wMj1RjePMiEg/ySTRtA7jjiteZLJ5+zcEmbRO88X87iVqzbW0qJ2NDN8OanFS/15Dp7UL
b4fRJoURXaslApHYqssZai3IXy010L66NNDWIH251nWomaiDS+wg4piTF1wTeFBeS6TQ7sPa7Yrt
g9bJG0vmCzsySVO//nOOMjcZwMeNxH0fuJ7oswLLJ1NSem7PBdo++XfhazeDCibt6y2EhT/g2lU3
kIqSm7Nbr6A2AN7ivXj2Zg8A8xmHD/QcAk+lfcK3LA+iFmUwNoBJkYNxRuzwRa8PiyvZANBfWmsK
DSFFGYSIWY9Rz1DAeCUYBc5/9v9QLxNdOdUIqkedhRrN+d5oZ2Rv8WGFipGAraVooAH59RmF5fxg
1Es3icBgFEi7UYF9AeBXfBJuQkOR4R8wjoxIj+GtxQVRGKaAzFaQ72ThQ0I690oKMryxvL6U+joR
RYEmcT3cOi7VvvFKGG/2ZzbFC++LaXK4RZ66267P7350X9gYCKX7HO3IAPn7YaT4PZRvejro5UjF
sM8N31thg5bz1IQpDRoeReXAyvYxvTt0Ayi2oFFmmliBU4x/kWyYH5HQp5AB0LKiY5XbC+f6EkRT
EoE8hx+zMSbSi2HCjKjKZnudKoaG3hQnLfUzc7ucbN4cv/PIS46SVhT6nHUrb42Z9ceR+rMvP0VJ
tavd3vUATNlKe6fqf83jv72dqr/rCZReLSiWc06yrzv9DCl0IIiEHYwrtw7FhTG5QJC35JepDNBk
bLNvJwmOAo7O6p22ccDIlM7znYJshC2z3P2ftutbFz5QooXoEBz+/IfYZn3Ro8FXNDoa+4y58q55
a+CdsAZMraQ2twR2DvyY70Sif+V8YPa+r3wjzRN1yH8XlpKoYVc82ayrXbEyIY2ie3vi1z9u/68I
hShzBqHvSXWCjbde93P8rnMHQxJQZSoYCWk/UYlRIEOFoUR0C3b4N2YtYB8cqE3ZoiVCxvbf569L
ly+jr6yEQg2Cy1TkCd6WOUrNp6xA0eV6WKdQTdOZczeG9WO8pg41lMqWriwKPf560u7EjrX6/OqR
9JNDbugbM32F1cp7+lfFLoAjsoaOm4TnPMQsIHcj9dut0XZ4nuRPDZLTl2WVHOCGXHql7JPYR9bU
vozfQq2s6mrPTdUx1YQWDlO8QFWt3G3vKtnhzjy7E+F0xr40FZ36Ef3+QmiXK1Ns8Ixeia+ZZnYu
kaoTeAtSNlEHwJ10b4p0uhoJbqbKpPu55nr2fYiTt1l4E/3p3xkMi+fhVB9ijbL61fqkWuX7mH14
omKvxpLeiWcGb8duI/SFiFZ9GMYy8SVAOzqO52+2PQw6m0952ie2iNEn359jHOWflBR9o/9mTYWg
QDpprf5ImudQJcLgTx9DiV8lQ85fnS+g5041anlzm0XF8hTZXaDMcGB/JTpNc3wj+f+WWP7gNoPm
VH1ynZysLGmwLkx4Ao4EI/xJf872C4TYucvM/cERCgUGJYs2e28nXKlmJNA236azQlU4VLI1vP2A
JMjz5ph/yR51sMk1ZcZH/8aJNlcE/YJam2yEVbPs1KEqvwglpPP33ICBSDyRFHxSWRqd/n9HkVH0
3VsZqJ2bsga0sTZkgpyKyX+JeC4zQvft4q8Qde1V7fvBJzkx35ui7mynfUyQMhUjTjLM036wg8sU
gmBH/ssvq+Yqs0Z9EapQyqDSspACvBEZCDhhYoAXv4IMenZF3qrZ08h6rCOLSku81tqzJwInqJ8d
8LXOe+5QJC0UVorEapKMuYg5WIyr1n11AuIGOitbiecsJJ0MaYVUDJVvJE+cfddkelkhO5ZOXdft
dKdhzdDSepyCTEb95VhWENMiwPF9OcKPhvx+NHlitIftNvFV0FSTZBFbdTPo/d7iZPRWeBXviWc9
DKjMaT7toU76Hj3FYtiMl2K2hCczlLMH4NS/ludtFcyxTsd81qbLCnemlz9LtbOBeT/wYUfNT2cp
rjaQBbeBoSCw9vGGGSRsxugXyi4IQZ3YAlS3J+8UMqyk7vfRqid3sesOf96a1aknREwMIp1tNUtX
v0yCdHw1rIolbCIpiotXg8By0TC5RtCykD9PFJ8sy52FlN5f7fcjvDia8Kv2xmc9uvOWKq2Bams7
vh2PwZJfS61eEMbzOP3/ruetVnGx9qJv04KfdywSamr7jSdfizw2JliGodfBoEWREuVKCioZaWE9
503uSEZXhMICiNcsK9kIJcAOMQAzm47vn32Cp9mMiSq+FqbutVUQBHocSccZ0SIkOTuJsduyRoar
SL1DtphaWzOhIzO373RT15/QxDvOcBg2Wfv8uWWqMdmlyOCoo0ADvvo8Wq5kODapeCqA9KrucZZo
TZblq026BYvojN0VW/fHOwLNQXFh004t5M9nCQtenS1di3+X08LHNprcAne2OdhPkIUUfYJHMyHG
ZsDpUA8jhcYsVvxF1NCIJyRfCYUqjKst5jILtH8S6E01bDqUAZ0kVQ86zdldKKY75Q1X3+aWs4RM
yUDkQK9cZy86cokYeRs2zN6ghwqSrGPyh2mQLbL7raPyvOvaqhekgQz9a3F1rirE0q9S4ek3h98p
strcuPUp3Ep4RmM3NpU51RZ0BU1g2yAMspcwQPbiEbxow+Q/unuD27JQmnLlntbfQ5v1NwaSu3OE
/HeUmkCB1Tri6wEIeUb+UD95YbBobbNysnAKk0xAY6bquQk+VYPLAip0j4w/j9RfvipHvqCFbRjz
Qsh2dPP9g80oLRBueDFUDDjj8NYYxAyZ1Um+60+NzN7OgcrpCQlifsfGfqZiiAwObd9KBGeWyEQV
YLwyZ4rQaCLBgGSr9n/pEWohsae3hZ23BAAwCosYFd3EkWrgE24FGAiN0P8Bv4rs5vaiecwTX/Ke
188zlxJV+GfKWAhre500GNB+QQmis+Jchx9LWP/wOvftjEO7RWhqQIA8xgXLCBopIWIAi9WVkjg5
bASdJ/WgWK8Rb6d+TWRELnl8m/H+L3AoGg+xv1QEWsYEgeiZt70/gH8Hub8L8Iy3GVfXlF16ogr9
6CZhN9eyIi8OROduFcRjExvcAVjkTzvASPzhU51v3Z5avn5Xo/Ds6Aa8CLDAQ7r0U9PtDLrQKiFp
gMV4xp8TRZYB+q7Bkbf7ssnMKRyWN7ExNXHNI07fp45dwEV25rONjucJmNz8o2w7XxpPmBiwDqdm
IHAe9Dgq6aPY62KKYqRUDEFJ7upsBKtsGtJMS7daGcLC8oFu1XkWIVeCzN+iy/3Cun7ooOAKXfvY
eEX8NWNZSRUgKlY+jD5hiotC++gb/2/O1wVJH5MP5FF996KJLRWd66SxJ+Nfp5z16fQbq7VVeOAR
PgHATOPZFmpMzBgRY8az+42lQ95y1jxKb6yOpLiIYk6+KN25nqUfz3g++1oNdvdpmkER1Cm+bQ5+
v3FH898RJZbL3fDxiKDoxVw3+v0kS6USkJoSdE2LzAZX/Lt0zthutrMS/oMJaV/yaugBPxP+bDW/
0Y3h3h7CAeIzyBZZK/epN8/3MHZNLatzENrYs/6jorJ6HEm9CnVgv4u3af910KTLXFN4mYmk/DQz
yr+4eSI/6ws+QMhTVZ/SFjADjjboyzQqLKqeMPe+ghzF4NKnJIzMknSFn7WFby7htr8vRKGjlh5/
BF3pBpEIQfW+XYLuNTs8Kz91XlRgYXDF1UE9fv5LyJENbnHYjwhwRBDHjKZM4WoHOeR3xXTehrNw
uhzrgVQ3t5S/dFrAVo/XaplWgG1rPHWy+ysHjXCZuhfLX5JExFA0d3W9xkRn2AHdqlpAar03SHYr
ZSgCNvD4/6zYQAB9haDH0vrm041E6CVb+tVwaQrU1XkK/MN8uLCHgWdoVhScVNPIaxA4h6dujXIE
aWfbqMym7oyBBB+5cVUMqNxPu7uqRhd0aeLICNToJWgoEWXWZ+wgE1mQwO7DyImMn/tgAqKOKJVU
zAkX+/HOnc2U+cMos7zYLDFaEvrM/zQH9iwUa+EBTYbIrhfCpBo8yyInD92q5yPqUMG+K7/BS1WH
Ird2wiX1z76bLd0/JXhdoBvWqoRwd2ImPl2OTioS1cQTcz+EMk+jf6l3ciudGN1Rl6WF3SeLxTyp
poNFGgiIFqOWQj0cS6P4IXlvwNb//YWYHCkSIztpvXPh2Hwhsaj/7c7fo/6qCEcZvsVDJGg16NDO
x+bJLjWFupniAqjjoUGcbzfiIPWlB8rukknnLABu4Wh07s3svUtS94wNik+tZOwWpAox+5Y4YaWw
NGo8Ew7PT2RqcxSzOTw8hEfsnffCmUMLnnzlx06nGM8LUsKQyovfk+ADjpDaL3o2eYASPbEk/bAW
OYix4/aWehqTpQYJvPHUPTXq4jDltubS9G7F4sVPNNwTeNn+0pKYCQHPtsYdg7dIopmxeZ5mkYQg
Z0gINQsQAiSiiE9ZyaYVQaaKr5fZmMle2OA/bzYGkk29Ps+QYBg2sDyK/8u0ug03jk/6+koBSioC
9oDmrIDhIG8Eb3+9ALnB4vdx7wlGOv9hM7VhYtfxezvlNDOHv5V6GNrGXZwbgyu0oz/AjkbGv1s/
TJPgNpsskTGsqsmtxkTbVKVjDXdI3NMz9229BkzlSr5+ihNof7ZmcT18Bm5pkPtVNKorJI256K6s
9IvZ6ID/yVfx83TST9dOETiTshhrpt5PTQoF8z4F25CTBYGzUJtk6H4rSlHrYvZ/zChoIbumiNXL
xkjnb5++QxD2a8796TDcdeZ6LKN1W7egfVukzN5KPWduj8Ctl/+MTav23p9JI4OFV19uYJ+m7Chp
LTHUZ0zh1YdgQ815T8GrRkDGUjmt02XJIf0uc12v3StpRRF4MAgBjHvirlAWYwJUFaBQy+cTKYjX
kBZgfAR1RHGDGwQyAEDSJGj3z/msHJ9PjLi5wV08C14K984Bshj/6ZrNxS+Gs04IXs+KodyCqfnj
5QWyvEI2OscWwg+RMq6qg0c1zTQO6sdrlFxElIx+m40hJhph/lE5mGA1rQIvQlCXRfJlmXNZfy1a
Jh2x6iFrZWmYJLgWwusCgD4qiihpOyZB2zZR2MCnpFETj0ekOEQLdTZnWycl5yptkLwt1eiDOnuJ
NQ2Ip8RmnSX334KzrY0Fd7xvOyNDNKivygUvk7bJydsUddQg6PPpNgQBek0oAzhvDR6A305P8UJ2
kHTxJKDo5nAM9MXdvsCELa/JDxd1Z0gCdyNWYRPKDZxrGs9y/krGbYI/IvQwIurqu1xfDUSDJrhX
wl8YbFr6pt1nyFaoQH6oMaiuVCe/TwiMrmH+CP31RhUQ9q5j2uULDuGLRSj6JqBwYzwfFX36/Jb3
tW91XlvxgNHTiRK1R4SrE8vlp3Ci3XOjq9k3hBBQRyYZ3D21zJTmPJ727XQsGas8BImB9Pi3kfTl
jAlcROxkOmvCzvIDYSB3o6HgHrSgAACaXYTdmxzqOSFkp/1ZfJCeYHO6wOfjGQ9woOU5h+wdiG7X
F9eCxQ6jba0ha4I4kfOJuYZw0bo/jJwk7z7lNSSQllqXa0jHEbFWDs983fkwGBa3OdBJ9TFDVaxE
k6ZMfeTsco4bBjyfRb3S2C6eAkMGFTyOXoZJPlJTYI8gmod/igkaxe0RU/LjGySc5+Z47eHv/fTv
dH94PIKZQ8pcAAmTDA7fLGxKqpua3J33o6+x7zfcCh1D2qTsNipwG9EiEyZZ6/jXvy/tnq/D3vXA
zZeZf+kpQ6q6JSpuNjreMtFrCRA0bxQPSRpQBm1Yi09GOFO+NeYWlnZsWeE9402S07voQqw95T/J
oKah/COBxUkidAwgTag6FK32jM79/JOZzSxZDiSZYkmyuohP2XpHcM1vLxQIJNYhXIOYVSgEjZPj
DEdWiM4PQclDQkJMdVOqABEI2aih31T5dAIf4pGOqtHa5KxcfDS5LFztjkiRPjLJcGAl+vpuDBuH
QSq+oaksboyGnQFnruQtBSfPggumnDyfjxzXcr6+qOC7KA4Grbe/+/x5ejCM/jobGH9+2Ar/hXlZ
k+hpEU9RPmso5LTXredzHpLjyreT/PPPBDdo/5BzST2Z2FVdYr4uNOdYeqUoxk0N+/UmJ1Y/rdsn
zWymMe5wB+FLN8qN33NdfX2yPqKDyqZW2/L2GFmvmoV34exb2HbwyhXXa2+qLOaRCuRJytcMW+Ih
sR7R+593tLDhDzeSfu2aI0jIwAx0QXSy2OU/ryjGdl4o4+IMq8Ir9flX/UyUCrPwWyWFoCq6lQ+Y
S7+Jk5njMNJepLQs6n7XobjQo/ylKy2xcxSciylv6y1mwV0H6cs7U+GtMwBqqfwtQRUSV01wOpX2
uaNlIw0jjC7zQ0pxYpBz0j07J9P27CwkOiC04QPyLWrLmdMXXQ0TDOjxUEa7SaYlaPCOLnBVsFCl
I/jJGKy+Nf6hsnfw8WLUNUfyw3194tiT9WcqjDaMGzYg75q4v9Tt+OO+Gl7RmDG2oEDwP3hdhgUU
Jct11oFabIHSXaUf2RoMTFQ9GNddD4BkxJ6uZODc6ctyxYKlHCyzKZH5F682ZOa+mPmBcC1ZGpQt
mqq7D+Go9OO8sQL3v11NRirpzWnJ0htjBvilL8Kgx1z7WvfkY7AuL8gHeURz+cOcDuism4fk/to7
/irfb87l52A1MgoQxlPasjAiZ0a5X2RetIWOmp9qRRpNA9LbNEoOr8TRoxPJwVLpnL1fpowtwTG5
3zvqnWkUWKfMji0W5JyfbTex0oP4JkPY3XzJZaFzh24e40FsYYsVuNirjdcPlctRCcOUx7RtKlMa
zJDffgkLR3AiFFwDm+8++cAhIOpsQRNiguYZkHSnNlgdY2/bnsGjl2eJLLQYdSEHd4E79/Ub6KJB
EZmzYFL+PRFejx1M/4lme5nDixz2x/FRmZ2qhsX/zkQ8vv1Q0GJb7uoSOOjQBgq5R6o9qfl2O3C/
7LFBmg/doMkrSNnjzN5j8OxoIjlvX4KD0wCRRPwF5YYmkRpQhOMt0fNeS4lPOVyL2g6xBnpoNCJm
0Kc8qKx8AGHB9F7EYgNF/lf2cPbVStorBII+YvAYlB2NCL1Ot7gDslwMGAGjbKS1NtdVBGvNx5cj
Zkv/gQ7eoVBSV5q757va8kv5qtWGsMBJrGvg+Jqjug/FqarqFayyS1SLRRJXZgXOe3b6uu18UneE
k/TyPRQvll6geZVnpI3mkBgTIZ5DUekP1kIDCpvaU4z8PBg2bVN5B7gEyDY0MCI+vbqfgL9Ysaaw
IOdgL1v7Hfjzb8XcMGCq28OpTjH/y+Yb05v7+VRX3mu6JXpQNMQm6rBn347PDupfg9YsVlUZUZIt
8+W3eZLokt8is0GVmef/nDd3PrduqHfAaXF5AmrKAUkddH/8BtQWTpZeNdffuazIn/xJ3OpwJ7Wq
jwoC4qlupLIDPKtC13GpX9kaGYDfeDvvaLMJQlWzzrtsdcumPzFpkaN+a1/Fjzzsr9f2X78g+hpW
RPp4ZvyGVxbQ20HcBMrtvKgx5AHB6w/vw9+3Bqt9Gzek37mvEUcBJqxR2OzYOtd3nGjau11/I1Sd
r0G7V4SAGrR3QpSk0VMX9or02vaE2j+9LFSHmrdOfjJVWWAmNJGT16R3Or8H8M80luawfwf0Gc0L
nAxZA625+Py3lZL90aQUO4DijJPTys7/qVO1SejJSmdO5jATLkj0zxqR1hrUSnT5OTPPjr4+HBo+
deX5xB+8rQxTT3a0+Pj5UwiKh+doVrtz67U7lk/Rz5CWxUsEqugewyzjzU6VKU9eI2fWSYoNdoLg
NbhHFosivmxDn1Ux+SJb5waf5Fieb1aLY2Tb70uYdcEOXxbzmXODftELktffdi5WT+dDrn/u5VG/
gaIhM8O5boe3q7TO7nTpJuEAJJcDyfodm7yoBIuMWGVZIHnBtbephQBgL04jZvxW/RrFoscvZ04T
Hnb1fQbYABjCJtFbSLhBxuJkOzVsMWzeNmd7/yVhU07MHuPzPAiBgJdoVP1zKdTE/eN+47epHLjK
sV4zmAYtxm4BDb6rOXmwd+iTDfzGUe6Qa/qRCxoaGjiMupSizgkMvE8/WhLlRGJGNTKRpyapi7Yw
Jw9yb8iCYOJG1YgNX5+2n/RSZoOP/J/SA+eALXz51r4FW2BGSJCwjdeKoyw9NKm6Ux+xbQk3yQX4
S1rf0aRQ3CZOIcvSH6Y8y6oN6nKInqc9TSXhnNYrPfnlB6SpDBItlJTLdPCRcSD8o8kQTpDHUNJg
SOLZPtxxsfMQpB70e6GPhBDfMhh1f4KGIVx1nAp5/bgZ1OXoojfbm2DOL9CSmsveZkzy9wjHpvLo
ySWSNDkMFrZoffY57ecJiK1UXUmftrrHNsqP9DDmy+gc6HIbsne+FKmL7ihDhJ3aDD/xai/djK3b
9eUP7th4dKcPFo32bj2slhWaxBrtE6SQG76sAWKrtmPqe/V1k+CGwABgbWnZeIL5Oh9nDBzsJWA9
wVYX6ZuVoalVH8IrmFpsjajI8vnZOD67N6DXPTLZODjNYbMG6slAh8PqJZe+6V4mxhNOZ/Baq/5b
4rYrC4GXqWJChRYlmTn1eXyRE8fLBjeM8ctoa3aZurimKvOpKIASna5+wZC3Vrh4HhinWmLoMBtJ
/8BNjVP+oG/cPxGIilTzn1YY2YXozQRIVSji9+VbLgpaBMI2Q//Xp41qcMzHLFDM85WgcLXOd6PJ
WeY6PTKyRNsz85d6aKEihKm+lUYqwoQ6kK7G5mSep342cuLnnFuyP1wLMBLpkoUYvOWyBnWkIVyy
Rs2VlMqqhiG7OxDNcZ/1ygxV2NStxOu8isTP2NhZsDZ2JySupvz3OXNc94lrbYzfYGX7mrNrZfrO
Z5Outp0OE0aOBCQ8on40wMM9G0RK1+5qCyQHv2dfjPYdK2iXm88+j6Bq8BzGRw7CwktjNngjN0u8
DiVEGWBNWg5W6t4x51XbMqJWWOSl6wvmfOm8R+G7AmMSs+0iYqLBQcaIXuwa+LtwtQoSxcedzNDu
LzKCQ48cn76fNemwDml7tJcapOC2ObaN0t1PtHS2OwjXbTLV1G94ptdlHWqoyyi4CGAT5EWBYwV8
6kPxsPSKqsA46w0NfQm01tUli7gK4CfUrIQcUCuyoaY+SLhJigi06RnFQp2vAYPUoVdwYtR9CGVV
CfLg3UQyg/2wIolploKC1aRIfOK8QmZJfeywNDFbIXNZnJRD+fsQsAqduN6xFY35fr34Z7ZSACty
H8BSVwlC6zmJTd5CcJo3AAYnDxFcJfkv+2AVWPik15As6883cNcCPa96V3vjGnb8iJ0ZCpoUr8dU
9b0DSvQMRFJQrk75ERpFvLQ4GTEZ9pSSh6HydIhxirna/gp2GiL2iY8Wc17VgKWlmeiZSvpg7VL2
Xd6DGSRvlYLO7OQDVTb/XlUQKgTPGcaQ4Fn5vXNFBib6P4KDXOsVQf2/d20UeAWQtyC/l7KKz3k0
e6RW1xoUugIGQlpAy8Wwg7KumxnwkXaAJO3mmvePyePNOrKoniCqpQnF/TBDSCheWcXfWC/6PRC1
HPaD5J7MTirYFoBoAjokxLaXCfMcAjNBOeqcAiirePH0KtXEqe9kUr9i1cu5Wy8Q1QyCroZi+iU4
pmwbUfLssiz5Uqx3trmzZE49NkBPIC1nrw1D4oqug1jrdW7MFju2VlSSYtazU4XpdtSv/v2sa6J0
Eq65+P3psH+Z0yPRywxKppm7enIZZYQn/XHVuzsvk/Sc5kO3awAu8TodwFtBS0IBMsi83f02ZAlA
E55D7cd4NNbdmwhRFT+FGFnfIoZTV8ElX5N4k5SWI5oNlsF/TkQxDZTX38CgIvI1x8VCqnp2pLLO
J9zbkxN8bIRiWN96DkY6hcoH3D7ozemybNQz+PoNClNSkAGtP9pMoTxyGzhu21Yi5f/F5G9tSRYl
qKIZfVulS7MEg87m4duNp1o8Eesw8U8zSPdgKQYBKQYHHOYiPzTCxuK6lumC5bN/tvqEg1Esi24b
ru0qHS1RVIg8zvNPMy85O2ao+Q21CaNz5TzVyqojKfZLbdkfa8BVeEgo9pOEbvI/inB0pFtAJTB3
1mXS2SfQvtA+u6kgaAI/oTqMGXn1sSKCkCHAQ5UhRSAkZ3N+jSb8l1TKlM+OMFxRbhQLYaPvA1HI
cWOyktERdJFw0n0+wtLx+d+BpCIgGdMsjae3yigzjK+10/JbkzShXGH/LdE4eFrtbaztuZUlKNWv
aiJ8T2nYXz5nPBeGhPmQ0zpxdqxPhoSoOqHrN1W7BCFqBHSgbf2gL2hJrxKD7NRdwwcootHw701K
1x+nKgtQpsynu3EN+FaDk0Dt/uAF3Iq4tsyO9TPLYb6jEA+KU039NrwFg0AtmBYyQhGaD5TWAkfj
WlS+Bs9tDnzr0waOMFHDISOrVRqNzZ5FoWLmAw403oyn4wkJSTNOCX0FelTaiAputO7mmE1AuSpr
a6rKPKYjzd/z4X+usnW0wUwgctUvZLMwHBWkXb80dp03pqaXXmxceVX9KeL4tYsQcE7NGr7vtvu6
hdPUfFB2masoxIka2W4w40yJ+JIptMJC6YBqGGHV3fhK2uYlhdbmaZRwTpB97H1yPxSXXicYfKv+
c4EQY25VFu5ZEzMGi5TctUMfrP2bhSDN5CMfSd52n3Axv+OXYSE+nE/cSbIbjZz/OpFwMabheSH3
BCYiSGUP2fMj+nzFIOGB+nO1P15TgF0Gn93gjAKVy+pGm6KOJoII3043pcDx+9mbl9yQTsEg/YUO
rl+JIR/BPbFlUFY0MCcnsl0sczeSXzlwLKcPATZaxMCTZWPn9paawvrtflAKczlfOsBnl82Xml8h
bcJ/icbpwhZscNf/nVQ+Clw2YKml/QeM/R5CcUnqutGZb9QDUsF4029HXDeStZgljCl71G+Z63Yl
u5BA4wEhZMIHIDlYGubTw9xHVOtMSpVvIq/DWvCsfyuN05rGsE1zuyhJCZuRuwHCGdd424iaxirR
7HY96FMtFE6YU7bK2wLjMwUApx0KrT6tXde3b1lyPkUJLfp+l+PRfPrJ+23l3K/AcvBlWeTJ7xPZ
U6qLnNqfXf9ndTTKmLokjk5jgoJIh67CajaE9rGpeFVdK+i/kMZgyHASITQYMP5REeTF6NVT1AFi
0BhQf4SGMCu+y86HVXnlvqz+CXjDEH++up6kWBBRQWwnrm+SMWPcsqfxyIX0buSDWd5lBROg3sy1
O1qNVIBw3qG/wOe4Gh81PT/VAhO4rFkf6FIZojvDBXNFHqzH07cV2m8bSbtWmUwBBxM/zlsfPyGF
m9d0W97DMPRq3YI0VFD90jv/S28rmQqrUbyUsU5I+v0gjEuJEo+Zcw8iW7/TlOXuuvkInaqeCw1t
5QP3e194A+vVF1ALLsRH8/S6ce3RIgPtn1PWBNApyL4UzfhE9izzxV4cNyzznZAuD+28bRMAvRsg
5nEW0vCkBsI8v2G6GsAQmVRbv0qgp7x/Gbg/b8Ghqvi9ajqR7ozyrRRUjGAF6SR3x1rdi0jTZDyo
yTbOQbyjQ4TBA5ybErpbunQhE3gfcRanF6c6LCKS+zlpO4TNMlgLowIaVaMnpAozayvG/xV8AVHZ
3MXauFsxFI7qEd5VX8jBkAtheau5sCX5NPLFvgm95DOv7Zvz5aaWtTPhnDq8PbqAeCejI1OG+xP9
zcouzryHlw1obVBrjBiARAbcxmetypatlRMQNW/c0ulHB1Uhw+49r9aUx/rdeRNye/FRnN6AFUol
z+pVs1P5cTEUp0UGHCfHwnP4H6RG1Yzuu9n2P6mSg7P+efuQujkMDQr4Mn2cFvLLC3LO7pNDJoZc
tYp3D0XMsbXPO3Ej+8X1Ot8i5Wcc7I/ikiY9QLvjk7JaEeIUq4+ZjE91+6KK/wgEZ4jr5QKRdtpR
qBN7eoHK/azJXom/bpj8X0SIssv1fOvr1WiOId5Nlz0X662kScIR4DHiyqOfD2meQAX+INUdN1EX
HJGxSvpAKgg2PRjmyT1Oh8uLB1G9Lx4A4V+HqQe+RT6w6YZaxcw8c3pAupURvT/NHqsXjxIEkL10
H68dQ5+Oa9SslbiK7VVEXnh3IlXfICU5XF12HVNAxvCUAFfskFrzyUoXCjHfYTK5DUwOhX/TZ4n7
WolH0AmFpGb7vIuBreu1Vt8KCce6zpAr6BYeTMuHBS2n7p6Aq6xp1Xt5jpZKBID0suNRwML/7bxC
lhjKZHH/BCmDyrGW1u/FjXKqWmLmp7En1FB2hQDSrH7vdKFJrKzAlrn0yJETFlxpFunixvSgslj0
qxdakadILyvYK/5qH7gXXVeBexbyjZWavL7HOFI7RBGAZNyG8Sb2rhDGoiqXA8PWN7e3ntUYfCL+
1QK7TQQCxpQqqmP/lroLiRm1h3vz/tTChKtwwMoR72HJOgLe7Rd8z7tDznsi5QVwyRttpQFqPzsk
Cfs2smOixCyBA1j85rdip7CLww2jckBrSs6yV1S4fqnpj2DqjVjJjrPMX8JfKydAtlJOY9y2pF7+
gIqi/wAoD1+KXL5Stz22MafFXA6ILuU1mxKd932hcQJ6/HLkIKW6koaZ1+YNs5HpEm9zDCiTEws6
97+vZr1eMyi5eO0Wxv3QpumSJ2XMJQVEcIrRmmvmqjDRD6qnJBeQXruQwM2Z3ESImxplmpWgWySg
IRcojcvdHyOalznSsB05DuG+hYhKJKQ0JcbWAMeuv0t82oj71b+SxBeYyfkkRjuqQ7S5AAj8KCdJ
eD64CTo2c2f/Ogs6ZaU1YHjrsLeQbBrlDzRaSGEjy50HNzEFpBhHK5/2DWJqY5T9TxJY6raiER7x
KUc0+2iSYDgqH/qhIDA5r9wmBq3mjZj30DY+xnQvDZbudt2r5Mq383oXXwnJKTw6UKTK/YaWA7HU
MA1k/kM4kQv7yfkK0aHOqG93ohbO0R7ZkqzWLN+IfnD7FWE4dqwpufNjYrklgpqjLR3xleyfX+5+
faZUTSbAdIrXCYyOp8t+lDUqx7h4IoZrPokOvo/CKl1hxKZnyNOvKYBMNktwcQErRDd+Px/KDvyc
ybWvnyFmbXxlIDlZR8r3FxwrWmA1btwXPG3Qk0LbsSxb9wpeWVyZiNTSLm1Ycym4qrySIE2RXW+Q
iJuWJsOiCWEfuknIB4N7T7drRmeYDYBNfKs53PaU7Pux/psQ512rPX7u5ic/7erbbGxEHe6L5lEE
FwBlQk1HfX2ElvH7cLEv3TaMnxEtDmy9M9uKqoh0z6kflf/o2SeozoHaRnBzRAB1e9WC66XkZzpE
agUtF6ylFGkEXqF6vkBiUKJUajdUplsSVCJshTupUpe4YMXEQq9SV+JdW2Lh2b/B302C4AeJpsaY
6c3HMof8QfiNjnofMLh5d7fjgNTKaJaeaVQLGuLIMZaVdZmBf/D8Sjfhi/jvd1h9jwIYDjCzTIfi
0fccZaAS9exqKXDXoZ/ns1QRBhnLFx6kV9chVDW+JkkEloTsr9uZmbqxEOSASEbP47ljhOvPtNS3
8nsIJM7zMO+saBg72GsVkrBvGN5GuNmXPfXhT5ZOg9QKq6q+SxDu9F5wR+4R9th4VmXg5vRWw3S/
/AQE4ub0mU/4PjTZuenflaE6EviUBpkb1tMT+seDjV6JoTVFcbLrH7r09MBQZ+6qpPBS/2Oj2+f9
NbvKHVHIkZ4bSzXYP8rC06PHkCgF0Z5L9EnvCcBahjodpd/vY8O2oyPf7GPo13f52cpiuS9r+shX
l3f/Oc8nJeI+k05CRrMqjSQnGWXJpQJY0+pNSVYDwpES13yID4hUYwl50kEmFfS3zfE+qeKNrq1A
jHlu6Uim55ASA4AfuZoelmSX0QD4LT8R5NLaOLH2RiGsm3SYrGx79vnTbYuJmnhZZaREfKndR5kA
SYqVp3Ur5jz8GSYGWa44ctZsp2n4RB1OGPAQO7dra2pcrU+o2S1rGNZ6SEYqiD9yp6Ajk4aUrmy+
+TzjsC0fX4E8CvcFAUBGZUvEmnZI/bShR1K2ih/nYWBEALc02BJE0M8i5O0nCZFG+tafpvnccLIz
5CFIpFXINSASGHJji2HwXi5xDABioxeoWDPiz0cq2UXy07+fQkjpSd7v3fsK70Y4NM8RsVPW6epK
qZSz5GBhjz6FYdmG4maAFCYMLscIcaY5Dw+i+4g+mWo9A2PIMktNFnXE9Avs1jgn/FLb09nM7iQl
Nnv41DIaDBXXSE6+7V9iwzDEKEbIKz21cF3TojtlaitmryELRdfi3RNuMOoOmwx8wWgG5J/6+cdF
Hh3vqQA+898SxMa2t7++Yhp/z5Nt6V2oa37XCDi57vqYXuF984VquxiDuvzTO8iVnwMksVcoFT0c
LKNOdvEmORNIYOImlaJME7YmEhwEJkO7liP5DDLFLttGd7j8HZ3GYAb+nvTy+BMhP7ljrD6Mmef2
sKtNz7Y7CbywkAXOuRaLCX7CmPspbxXf/Aqr5ZDJFQKss8PFLth8rGHOzQ0j3UqckN807yXvuNAh
KqS57jI346sYaK57eKEImAI5nGCCMF/b1gbk5okhgbFPoE7W7zd4KrEfu+8I/ZgH5h9lrps5uCYf
9+Kgrgjxnw2SDguoGpfCuB6ZqX7TLbwcs2LkSReiebmBpi57LLQGoIh/oSoj9V9PdCN/qOnTXHrx
wRpz40OofD6To4v+AdMuzWDP8dylpnFoZgWI6o6OvAxa5eC74R0AOOYebAOHPjS9mvlMac8/KE3y
tgG1ILLqWoJYwelZ3SzIMU0VjNbfCn8YjU9sWVgOaX+VkkPzbrJqgd/M7VMBYdmHRCuCdmRz9KzL
TVgPHWAICdAV5Q9sRrDkBaq6+7hvb9uAuRBgNDeNyI2ZhuSR04dfznASzbKlX0tu6pd9BgVLsWWp
eiXixNWyRBjpu3v48ptKWzwMH/l47xra6QvUbUbLpihKfBr6T8aVsuC2SUw1iFZTcf1VXSyUJ1BH
bqeGx+Tkgj8faf3pdXlKNjJ+OFX/mg4MugKw+0dW3T6PXe7HSiqfpwPRdGqwoESDsHizEAVWJnXP
zapA7DOl2NDAMEsYj15flCjXEBeHnDDueToBuPy6i99VN/fhOS2qZ++lBNSNWMuuFXiywn9WaKz+
VJRTtDBVZNaVaXWcd1croW/zWYl7w9QgnkQUs/nMyhiaoM6UBrQ+U9J5x+2waf87+NFC7xkXvmwP
64ytG55WUqGCZ7UKuavuAfb8wq3sUJtoZl18gQTDRPzys+aQPrT22GvvWCEbcTklJKI4edkYN1ES
fyG83wlIx3vkgdGW1BUS8K9sOgC5V8kYNieGHhyqicuhcGUp+h+DON+oiwqJMEeOwm7IhZjFVt+u
e3VHQoYNohK4vw4Z+4aIeC01fMY8ww4pOnE5YktOKXzp5w5G0Ysd3BXklE8kYbsKwjpo1qoavGUZ
znTpZKsC43x3j9g+GoHmak4BLz95kCI5TK5i23mzgLyLbcYFfZfRt2PEQ01y9iAcYQ+7vX3B5dhs
Xu2T+Wcq4OSfs27BTFgY3X/9c8EbQGNuYv43TkOejM8JOMToGUEyY4hxPyciDSpwh2t5pSRdDx8s
KXebjCuIvLjr81aRXcGBTe3IlJWBV9vnMlapd2XyrCggJWbcgySler7gfATWs9VHmsPaX0JqKl5N
C9oCWPthsWe6iSzWv8/Dz1YdXk/fjsU++wstiQ2g/rep620/D/FLRScFY0uQD0qDwdBxqyTcN/27
4lqgJlTkXyGuI5Wy0h5nSToUR3pC0Al3bMiIBnOf+z64Pe6yAJ6St9BQVw22Bh6O/I9cGYOcSCy4
9iEFHq0sNZO0Y1cgpOjh8msU7XOOlrDiCAmfWv7LTusLjiE2yBPcW6VU8jANGkpAj/we3TR4bV0q
V/3/+KqrCFTYHvPDkHkX+8gURi4RWv/+YYXMw513HsUoVAq1gFw0WEEksY7Sx8EXxcIBtIYk2d9P
DjjQ2QGhrSjBSvcPudsjINF7jYUSF9EwTaHB44c7QzsZzTjZjON2UDDgfMNVs9OWXw5sGHnPWnPx
lyML0a4MIMqauzuU2WausOGXbQtpH3lJHelSjPxppW0s0WbXxP5HhU5cdGIU2qvX/pmFQnoG71Yn
25oJRnBu7nREt20Zrv6z6W7Ajd/aFn6xWfRVyJYzdlt1zBwUDjI8fed/K3xrkkC+nLxpiY2Y6MRm
6lFhjBzZyfFt/pDLsWsQWBtCkw49na/j1hoE/y+AkxN8pDVEEJB2srDavyn162vgXCyy018tAmKr
rwR27lfgsv2T9jzO0gM5QCVPjHfET0yyZ+O4ylbgDFZs1Cy0tZ5+d/zAIJVbSvaD+wAaN32pZhuK
9vDnDrZvXXoEALy6CcLsD6Q1j2Zkf3N6PlzAvktqB06w0ev2vteNJkzegGk7Frh3rYde/wV2oSUX
3L8TYubo4IMjFwPvKusYf/BmRgyuhxbIujE973V6ikZFEJRsFIGjWJp74KV5Sj/xlxPsEqajvesz
5AHQhOv8CtIOQ7Ad6TB0qLaGghOsxuuc/cU3zFnC+UNjHHYNEVrzE6z5rq3VDuPtWtpm8r6k3Go4
Ntm5igu2TJWsHU45qQb8dNioc0GgBnY/Ib70L3TsJxqJNLNKNHEh3robViQ0Ny2yF238maRZNU9O
TrFi5Hk9H3N4enhgQEysLuhZyQ5okKenYbRW+HFsqokVF9isjm16muRO1X/lpHvIrMP+J6wEFJXK
ImwsGtv5edmq0yw0hNeihcxsT7S2IZDdF3BilnBeOjcatyJOZdB6fnkI1LWaPDnOg80g09waTH4/
qDaqIKPtclKzb3YA23iaRY5ar9qn0kWIe3HBAoc92u/m9E8Mp9iecyvQWhCW73uP4J4AIT9CWh57
2OmgshSLJtMnoavzIaTlcntYEiQdZIhyJ0CSKDJ7Yx/ucGXq8TALdIWWsxILV/cIEbkgs6MGP2If
hIQDNMcmUsh/N/YMPvNbfgGnaIGrbG58vKBv4SyZ3TCL9arec0GsJ91ABYTJegl6O/GmF04OiJJz
YptX5CySFXsSMj39CvR66Zoi0MX3laBv8eAV9tl9CjZHF/HXpSC+AW2y5gDi1T3AaOKPysMg590X
IkeD6m+ZORFjktGZeU9qSTqVRiqg/0IoscAcPdiuoiJ53n0BAodDEzoUl7E5gvx/nAq2j+xsWlOV
wxP8fMSHjWuf1u795+nJMk7eUQ/eAfGXvOXuQM0tIBt/dfLeHZqN4znfM1FMAMK799XQHgcxISf7
Zk5GYtqq7r/MzDioZi6Ey/jUdFpRl1iLASevj/rZdh85Buk/CyhM88HTuMqJYgFwF03adWjXu7VZ
reJWlOljHBOg5J7H7sPNmw7qauTIhDr+xrjf6ZY4jBQSAhJ7i6Fqgpbq6tbKW0WFe23CwOD22ER1
y4lFw4qp3g33utWxoUx9XjOGB8PaQzAMUPeZUfg6cOYcnxPv6bYZcaiC28W+Xf3hkk++zysu6icu
JG4QEPHCtdUkA6mJjWYYAGtqgqWF/Bwj2tA55o29Ch9tA1icfDjNbANTnXPtajJerVne1NBf4rYO
dfyVDHgFqYzzfXtnM8XeUMycGOQLVfoAZFgdeA0QETQhQXzxuFEJymSN1ElcGocahuojkfktbg91
z9Hj01YVnk8YMhhV72DyhwNGaKjzSLy9aT+4ZVO9h3zt3RAkLPoXINvxrysqp5d2OKTTPDe6Wi14
6L1VsBmb1CwwaTClW5nCFFN2VS+fbsx8AMnNLMJNXD8YvUf1wrCGFOe75sGkcf5J8MYVPsjHJ7Lh
uOXUUsXL6PxptYfXtmCp7k+dyM0DIh4LP40r2xroNeclTDP38xX8IS1+kwm2gVq2OSWPeT7bd9cM
jfc348kK4tMJDecVe73RXG/gGUv8W67WxsFRXXFd/3OK6h0lo2O90SPxpiFe7NUy8k55zYfDxQeH
hnoEMXA6Y+r4ewsORzH89kYyDYSvihxfnqMucmZ78Ka1fgLe2PUqJRZL0dEsedxftAR0Y/x6tNJT
L+spN7Bybiz+3jPP/1M3C+jMZvAdCiTEOlGIjwEyOVCZ0wYsqZmr7RBUKAQhm63Q2JwGcYdCKNv+
JymdFvMSngJFVdmMRpT5wutjQV59/7KaylJ4IFo6/jXpfI4us+4Qksn/l4TD66bYVFda0IiuNaRX
9LZekkL/2TnpqjsH/KIvm+R41IzKJely6PXeZQprG4nHyh8WgNssP3CxW1QRWhJDMwPggtJsv03E
GJLivCkdTHQmJMN4iq3IJa74kiFGis/9I2dm65crfnCLVQLtnCH3IIiPL0a1VF9TzQVX9xnJnZyD
P7hA8o+nO8aIxI4CEwsvGN3b/cjuW+/kaNXe9VVnQvEalu0DtJrX3BOg7ZbVUnfBntpSB2AyUzIv
ueS7rh4WMZHqiy51MKer+tePgiov2JH2T/NKXNwUmU+gXXsVYxoyo3gWsUwMmgGpOH7YBAcUFLif
My9JduAGJj8vI39i5IZH7mqY5+Uq1QrAiguwrf16a7W1xojvTjTqvB5kqT7Yfo1I0ppNOpwSqgkW
sJNwJ7fIc+Wqc/6IHAV8cFgcL5dGuOc2LNQdH6sqkCKvJSIFg804wOlvZZ8pxKxVRIb8kA5auO2x
DW8WsDODT7m4YV8b/z3IK6qt5tUDRFlIoc3+fij6+wX2QVWra9VhT8LQo735Igc2pS7HUM2GL6W7
picZI3M7q+PUT9pPNThzeFEDdmKtOOulE2DfsC5FJeKhOg95gdhq0CRSVeBeoQOdn3hNYs2KapT/
tUJsUNDDgP9MNFwGR56hC3ztHtmV0ats4+tgUkLHHkqQq1tlvoP87cjnXtLLCBzF738im7jzkQ7q
0wpxh4+tCRguFgXSA9wYeFF8aIfoWDdH3NWFO7RGuIEDBVlkgVnl1v/n3EfYW9xJHfpFjD4a5pVs
Nag9jKLTMZMutlLSad67nbHLqszljAxdNGwRbLkU2om2BmnVCPFyHvmw6oRIpBGHkCEcZTS/esYL
56GTH2V770T7vR8cYbiXI580CpHrqvfyoiqnZTi9NEUsREEtfsWhwNdokjDah1KssNsmt8HObFjD
fAHKXzLWf2caDxFi64B/uGtDeEHyly2Cl5XDjeUbSFA/QXA8FPhVhgaxEylE8oh7Fq0WXyfkYRl4
bGRzxzmo2XfKDTN52yBDdkw7rY/OuzabXd95M9iKrmfYCAoCikm2KK0GbsT2NTZSgmm++v8LXc3m
7ztYm9amKO3MbWvQ/PM/4+MmOnXKGtuJP9BDlO1rOiRaTogx4dxhomBW9jvkhG5xBK+aMJspgWz4
gNuqU/xRfZnii5xcAa2M45Ys3R6CmbQ7Gbt6/66lNL/VJLBs0drlmonoyLmSWNPKsAA2iScizVdB
Ka7cTbxBEs/kI8n6vIWaTI41wbsy2A1rIVPNVmZfcytC+u9dLn09PAuDObzumCG19e13/N3XbpTt
Fxj+petjY7Y+ttdxNdGSPl3w/HkY9T7xKPkXrb37jWOwiTP/pUxJrC/uwCRG6y1eXlmeTOlt+/vk
P13Ta42asDQ8K4Ow9R472cgnoxE9TtwvRLBXrBXp7QtN7CLH9D5zS3h297RCaiNp+CXw5MIrUTmT
W3YAskezVPB7nSqmXICuT8dYoZ0kAaDZow0fIRktOUSba/GqInpBdt9jRC5bTpIuscY44H7Vx6dP
BtwggPEaLLwhtaG1qiCwMV05FKWsxPUpMQXJsEUU2QgkcOpdPWpnRRLrp0Rd9IZP692XQse+2vym
CrR36nqZw0m05U7AiLCeNE9txgoAPeFOgpZLvxAS1JNVALMcqPHxp/wMN+cQPvOVUXRaF4Vuokci
tM+dHv+UuQZiHQO9Wi+bLERvA/siu1MgZVDzeIhxNd0N2LqibyEydx71/i/ps2J/L3VQxLjQmbT0
JlhJsoXyuKqP8kjGIIMw4Sv3wwcBaL3XxMnv5snvo7OOFu0cC5Ys/mMOSkbWvDaASdpWXlGXSR8q
dl0cCTumAIPtdVA55UqjP4B5JT5pNK2jgmWRVI+oXuevrkz1i+xF1Y14lKuw9UtWlYU3eDCY5cXr
hNulJHxjQZrgPGz8WP4DCCb7iq4HIXMh2UA2O3cede6tsMAphjAIGDgfER2JztNS2MvxKWbtcggu
bxo/eyoodP/ZeaDSaXAxS1p3W5a+XRWOVx6lX4SP1KD1m5NqAf9wzwHZ4M+f3it10E0ild3Ci0sL
qM/dcM2bbnAukc1TnmA3zQQgCFU0oTjL5RE38t0Q6q2SYnNlp6j3ZSLTKSXlqytsmETP6E/1zmTx
92mYtyOAZ3DPgmOk15VyuKf3d6sgGb5dMQDqxVlVgeyUsxRKYuIcqQRPtgVZfF7cxwEjrmpyX/ET
d9uYkL6fywAQjFDtwp5FMDgPiHl+u8WcQwlUyZd93jaHQ85FgrolsGf2devSsoqozpH5PGxoLb0m
c7Epkm/QoJUZgq8+LCEmSrtrrJt8pvzh8/fQQGDTF/QvT5E2bFtnOgLlPLvG7jGZMxEduNa6RF7J
FsyBnfRpfgYL/WMfQuwFd+DOqmxlczuWY7AXnogbj4aHsQFDgVt0g1cUO/4vPN6Jj1pFdlLxaHUd
6JBGaS6dBSo/EEzD/1YXjIPtvGfc4ee/HPIpHulIc0VOAiCa0gt/GWc7CK68klil7bFvLyBl4mjf
njDy8ObpV+8oG8xQKyxkdav1ZHfJO9YVykhyPA4U8Nb7Ynz6xlhz64WSLodQA8uZIpg4HrWyl0e7
3+jkJNeIw+s6ajf+l4X/F/3IofveFGBuWBdQc5vyzdy69mN8rsnioldrykhDEeyXGG2AbpJukwTE
m/CwhzGbzHfte74UQMjynS9usi5Zszq+ZpuD67chqo7ZMxGhJQDsL7F6/YlpRR7c4W8/5+sDKR0t
BzkYL8oaFWDLNBxuaWm3hicqMlfpJuiEu4yd2RfkRP69IoUCkHzXIWqDYygaTn85XQwpPGUOt+Xl
QV4JySJUSj9JuxZFX5zlC/EKCVOPWbZQyDcUPpafwJdXDp4Odxp8t6BVosGhpvdT3mIgXqM8Zgs+
L6Sh0DSVaI+reQMxidi0h94lBTQ7umruLNYLnEFEqPvfWbLl9ZMNw9/uez6USkrg7LEg2pGAQwX0
qI1E9R6h3vgicNtVHobEDzwc7WiYTWoZya+wtM9qUq18rCqeMP889u6vSZeAWQ36gAO26Z87KZta
7t4XS8+yqSwtYeBhfPa2UiVmWd9/NguHOpmFeO7k4CZ23cUk4m2xCFA8KqgACvbqhMNt4eRSvP6R
0K0JDJlgTIMCnRWp/unI/DXBRFb4tQ7ajXLhM1vlHiszJXPemXDe5o3pAIu4m14jlX6+8rAYjtnf
16tFNhtwQh3GePBCFjyCqtxT5dtIHPAPC9zihFyeqNu1tbR9MP26akl5lrH+ablpoR4clR/IOuqb
tBGhcFGUYoXNwnTY4iKjaF4E80zOSOc6s4D8GDYb5R+/ISoEtNjzjSm3upEpgrDtB0vi68ib+7Qg
VUVs71rt0vx1NTKHFtx6MwCJDdlgGEcj1CSe/FGNFMvzK23ZIs6TAygoQCnRMbuazMEJFbLXxXbm
7BH38QqsYSePN4DbkjQ4HYYJbwt6+m4dCmvc63vXAcJ9CaPnbrDfBBu5xrhjhfpWsVwh1tKJl6V1
4457JR5lAaYh+r6G0MY9UnXFLn5Y60ZfnVxx/60Lk+hu8u6Wf1ls8NkbSTdU5zgYE4ZAAl2YjWf0
xPYUNIbieuLU7K6NRMe6nQ0dEPn4R7FAmIaUpj0kY2t3F+MICUu5ey5O3SXn2CXpNJrd/MsbqCxn
ZTUpZhZN0X9NeqhQuPdgpdj4CAoe19bfhG7JkFz4mBe8EF28jobBKgEhpTd/X+wt4Td/MGnyMOuC
bJElI+Y5qqs2Qyry7lfx2eVuWLZjR33X4yVR0JPkBzG1082RM0z95HnAO4Gr4igwn/FtKg5sZ7YA
2uILh87ZJmSEhVDWJeSz2hC4CUQsF8EEZ6y3SJJgQNYFAUZ/FcbkwT7eFUtCoqUeV9jZeijXEHL5
9tr+lk1zGky9nBrmps7VX/kVRWeXWCu8HeBYwNvy3sYreRl9oGZ/1HSbCzH+wcbNrmnch9qKnoDq
1UYANkqojlSrQLRMcwJ64mTp3Qg0S6x0cmGIykPg2ukc18pAYaWt2+eDH9DcApsVxubEUxdxqWhU
UqhZ35oMpPAuTDglM9z1rtYKHT0Zu5/XvkJpeex8PCnwKDd7D9aNJ5dzUf7gsj0rBKV7Tdoop8UP
MareX0liMgwMrn3hYtO6aTRMpj6hQsvwutiEeox6cToPLfmGskq0sRratVMPxWv2qHOsEhl/KEeW
lQV9vlgnS6bkSl1+qLzCbxycdd7lHNxBXYGUBLPW2kLU77RHuLGdSPpnivvf00il1UATrL0g5wbA
chXKHA3PQ3I//1A2IdERZAKFoK/Gxlse29LwwrCR6YTZM+a5Di8eiECiyt9YNVGhuID6xFpWLwIx
BhALM/qyJmXZkKCPAxNpf8dZa1Bu3KHJcsCLF3iGSrFFCuBiZJihaj5HDokDOWAlWE9WRI4PJPto
FBWpUUS3hG0pCMZR7QTqwJrJUnfR6VkBMDzkcADH7eFJHnA/3BDXpKjngFxp9p7GyO7MHXBRmXVe
PxmX4OwZklSiej/vPKiH35s+np3oB7DUi6P9UlZrCTQffPqEKzgwpcyx38/Q3cjNxEB0IoLxTdXe
uxdDRcoSTAwO71JBiuqqsXEeCWZhj6BLr6QoQXYVpjwRpDnSdj6V9TEbpTnKSVRDQAojExMf21L0
66sPKe5DKZQs+wFBtN3dy2ULXpgtEhenrdlPluL0ZqbtUSJyPeLqIDhLX3UsCLMQn7sLIXTEMVgJ
tbbIzWKLg5TSXmRdwZaWe07wGsavmhGCvJvjx9ttdFo2tkgEEujckTUdz8B8C4kqUR029hveUISl
ErD1BOMg4MosAbqwP8h4Vtt4ltnR/AAVf/Ep2r9E0exAahwpj8k/UnA85lhJltbEcE/4Z8RcOgQA
7pcb4kFNlBi/MiAkNAxvWFYYxzXOix7bMxbe+e6YfYTn85UTTDEQlXU88R0HhUDBQ4Y3dh7+x81l
ZsFzl/okPWSEMBcdQHmAW2YYDi+crxuWbXGhR7uFzJx1Ug9tQZge1SLlfHSp7wBvpKQjsZg9Kido
SBAv5QgdWGyfSaCWXtazwCgc3v2sb4kzTW9vbkavXwK+H242Ex1JWzctM694G75s2h6wx2pkX4Ad
jMCsEbfh7Cm9vZT4zmG7zwaR5+yQtqjZW0K/Fa0UQUrcBgYAurG2lknVGJkSI1nfcUEEN3+AX+2H
XEvoEDUmIJ/BcdyvxFeQWLsKXgQHbsEWn434/ywgUJNGgv5ip/uHJvbQiZw+m/sbcswKSh9Kd+aA
wNg9CLv4wzSM8K/6v+xc88ztKawCqtW3JYgk76+WyYhcvVvktjCa/cZ1vjGh3Om/its9gL/3TwcV
qL3Go0FxpVS76Y9xkY+ylprnh26LIxO6CBNuSngi1Pfg9i9PI/VPvd2nLTGPoLBxQ2AAfx8ntlzv
D6CqmqNKUitU842JOZXHuj2KBHOH3Q7CHovS9DTxl8HOaarVugMvqD9jdacLt8ikPfCPDnH+EcL9
zuBE2MTeq0JGutPS0eLAlQE0PZA94B24OOpWbOzMGv2aDzHqhrfoZm7elM8HEjPnpEb2O3VI1/bL
tDp64Xs79YdtC5abXOkP4yVTAOX7A+7sOBH1236QD3yRyqj/EovaMsnA7i5cRO27Tf0HfFUlCQyj
d5NZkRB2dow6NKva5FoKCcHzMwECDecNUCBGbX7glhJuUp28pgGFeXqqa7FpWQqjrM02IH8bXIcr
4N366tWE9uIgHIKhM57QB2Hp23isy1CUJsv0mXajHhgDVfxMAe4qN/tV94Z2bkMlhUWx3MEWic+9
coWv2YY9neq4BX6UQxGSV4ARmCE0d89K0NrdosrW9KmiXYsLuwdUDBltDvdmryHIsoKC+Y9tsxgX
zkn82p7O8GrpwPhhLe1nZQ2h5uJ4+nVwxHnoldVTDcDdF7tzRlJgmtDfonrV4dML6TBNhrE/5SYH
9kg2dXKwM8gt2WlRFKOxFkGz7JrBM6clHaDE0NpLIIMMEc6AMyRydZck3zTON1gMguk9z54ghIZp
EURr2SvCb0iFZqyjmwpBWmhg+wT3w4/Ya+iuGIVuLzx9HENyo6KvNSGQfNkQ03bkn+HzO7GJbHKT
JH9hQ/ixl1sJAqwuoQcBsOcQXYZU6n3AKv4WhV4WHv2sTPvBhqVknUANITjuFy6AHPE5nC0+vHq+
ohphRcD0wE5rXRDlgVfLP8cPwt2FzBIPXBVTfWj8rWWl+cs2/j/P0s0VRYwkWw0Gtn62U7ztgKMq
v/p6z14Ldyx5J/6Olk+4lUTwiVKRe6xUKE0QUoRwClU5VPgdiwfkL9yYJckf4H+kKxtfhvy9YkFV
tFWcnK+ZMhIDMNCNi6Ojc3FwDN6uLO411EOg/DqnEWq/ZJzHjXUK5G+mJZALbx9CKHaBOD/QNo1s
9d/alHJlB5A0tThx60TCq9FeTKe5wE75Moa5HjUVcnoMdewUIiGuv31ZM0VzboqAs45RZUDrvEsl
1SkeWcVB+xKcE49eZOC7MEZD3v3QAJNCm7ZT/3mNXWWWd/Q05yBJRwjoVHYZ/0HP9VLyOSLG7pAu
6HmUsjn0mYNEUkjGHN91Y+PtNNFvok7oYXnwWjlZ3FtxpC1JCTSzyP+ElVrpGujfCzix8L+nzbx9
iGXjEQWj9P3zUF5qhiM5X/cwdqS6eqfWmHU1HhR2BaCcPfIWJsxzwuHmVTThbIZigSiLakA6dKu9
5NNVgbjaye7yVOFIwLzb5KrpHdSMW1QK1hMnSPz4GJxJUs058U2nSoAZZZTfg5N/eUap0QotvLjS
tHtAO9R7JLnV0BM+VgxNreiNh45fiJuRvg4ySqv57kVpHRIlRoMK7KciAZeu2nDusrzSt1KjCeeh
pWMqlnvCL5pYWqIsFEMI+KEfGjIuNFV+vbbcQv/0HNDIG9eyajzzJUrIcYfnA8Z8Wk5BRZDICA7c
w3kvQoOjWFAmk63647gXM8CxDJ4bWLj+OlQSyE/qdjROn8Y4efJIxtTHkya++UIKBdDHooiG7F/3
XBpKjL9Zlc58aM4sTSwzNeyirKFy8NacZDtJmJBIl8h3AlTVDtSH/3rwiqbrPEA7VvrXx5RRj815
MvvV1EeHScn8F+lbJWRcoLG1Hfj5HFNsFynz2g6/3h5djwxgDI5EHkr5KE62ySzfb2yxcK0QXuGm
j7HGhfOaigSFfoWzscxYjKhmqbRDQHUZG+U/vWWL32TtMcUTFF7wlExMP1+6MJbHRw7SK9bqf+sS
2LuHRoQpdk8tvO5ukZsmYmvaokxHcFRMXw8+3PUvfWo2q20lja+sm+60TsJD/tukz7cAwgz1yhRm
6BOPGYKWGfcZIzFbF0O/TPW7Lr8w6N41P4WqFur1RBECH/BxQQ5yLM0ql7I9zV2iKPpbbVMWFF2y
69E4nM/2jOQb6KAPVu9hQD4M82f23RWh28rUlINWUsPJWYpXMfhvM7BaomXMtNW6K7bIBejERNPp
mJEknxos2EMBztacJFiDIf/sgerkf+P/aqev7+rMGOGGFzYAWD/7c6JOChA7z4kbht+OkHHxuWs1
Xqzk6qfbjvP90JDCUOzI1p8GVd4Olt2UAoLLSS6xfziEm1JRJNOq/4XtyoEGl1Mkdiaeryp+9PSl
0mkv3WLFEJ95jxdtH3UHB4FNvtgTZDHq2xMsHjbj7+UWTqUVak0RVsIHtDunz/G8U1XnF2k/trkK
pTflcf3BmgtCOzznxSMM5Yhb0KJbk0pkiNXURYO19jU4kSEZSLNY9kGUQgsy0Fr+K9AYjOHsDmVy
NUuWLwEm40a6oSNV5VUBKmqxFafT4msMKnWVaUnBmhjM6Gsm5lYwVQ8a3yZHzf2mBtm7UkCNf9Vp
Ju7isb//J30TCV8ZEG6o7+p8hspm7RVeYD1MjQArpccDFIzzWCarCIAo0e95VsI/bbqigQgeLlzc
krBoXwzeiFcqrkUhG7iRIvhpR8knoOtwKFGFYXk4gimMbeR+1cpUwsGkKn3heustp4wqm7uIo2Tn
Ryg+In4a9Agvm7g7nn403/ff5zYvJN5q5FLiMXn8gq97jBbJuZHg3W4JO7zNEZmAYNLI8xbrVA1S
DNOUHeLELDIuBWXp/tX5eqybD5RU98bL011OFc4Ykzk6ZKRJVEjbvwrHi4VmK5BoM2VNLfnBEac3
z1c0gAqbVkzmf+kw0R81dPJyR3hTbjfNAGXxvtJRraG1O48LV3SfmOrhLsN0YQnIWSo/0101RMu5
XGrq7XiDxHrERybnPE6VAm2VWeasaJtU4pb2omisNIuc4+v+QuNIijqmEePhFKWJi8B8GY9rvScn
KrNjsxrnS6Bxn+fJSrrPYCym8pI4teiYRg2mul1uYlaLh2Vx9P7Z7IzpjqF1LLZ122oF7zQMOBx5
AtgXUDu5g2ZBAbq4T6al/MOfrGuKUqgkJ/cPBAMVGLj0ksd+/GFewWHEzXAQEdcA7XjY0F/gql0h
//fvP6lS245JRV+kBVjvesPvhx6IzxNdhgNU80DH1W9fNK/kWC7ddhv+r6Wa6S+8fdwTbQf0z2+C
w8sPUas+VAwoVTzg2qkjS+m/aUC+mHuKH4fhCKOy+l6pLYiixdlhC4DWtyImT0T9vOvst4LRwsXp
67NI1BpIdZo8Sq1PNi8t++tALTmqbIN2RJB2AtT/a4ePMOwiE1x99OqhGGhHBG4wKu5X5d+9TLvw
XzpHA6g4z6vX8tB9vHZilpz0Da6bPdSnfY+e2pWnsDdgy3djGSWAw3rCurTPpx8gyO1PHWh6BQ0p
bVE0+gB6mfiAhx0hPU72BkKOcFT2JD3PgTRyWH4UrSPcRS8eillTQnGykADZUSyH4yS3GpiCoURN
FJj2GQcRYcjKhHuF8PApO//i2cnj2q+nw5uiufLWq0+aN8JLGhtImbVxdG4AJIiTRdHSPBeuGN4G
14ykG3B71n3L8wLW5Azvwy22md5KCDfDL0XJSFART4zozFituYCr5y0Nlk0ncq5HAmcF1ndh9USr
o8Q4bxrkzOrR5H6Su8hw4OCQz9gMbwSTt40+ZBccQtYWAFA4bfssKKek0U0hHTL+Yh/oWwX6wHRL
eF75RFSWcjOtYOVQRGi0QFmL0O00d/94hHgp/sCzFLXOftqObU7xL4u6ZWjPwHM1AusS1Y98t1cW
EJsE0DxfilfW65C//Up6LBJKev1kgUUy7Op4koEGdFMRbEi/yGZ8ejHVcHZBM12d8DoCsELnWhnd
ue6eydw8qCnh00Wi2T8Z5Q/DV6GKMa/vXSkK3j6ChQwoomA46iQrbXyOPHh+vISI8kT+jPRKstl7
h8OlCwStHAMJaFUPxjUyL6IPEl+IwLS/CO5vcBBKQ//wqNRHls9UbIlnWCGnwRrv9bK+PhsXsiVO
mxIeMQIAJ6f5wxSg+Wdi7ON4YKMkY5Ev8SJdqQjcgUA6xUPfYL7BwnS0qVjqZQ2mwRpMCqIyN0uQ
Fiokb1kvFe0C80458V2sUm9lmsU7wZLpqdnI1NB5B8HpDGTXtmnsqJYs/mtd9vyPLFokcSSwmlo9
489ysf1Z9YCSu3fTWs8hNKj/HUev9mo7fZI3yBcVuyFRZevDTiyiLq9v3fXrcaik6yNah665xptw
U5CCy0/EA6CzhblqcyoVaeG3KW9YCAj6MLfJeBHa/MYvxGj0Yf1HAhT+DVBcVuecx+fDt/IhbtzC
nLRhZFzM0fYKa8XM/pvOcVcKO65d7e/uDqFjEMUZwfz77uKx4iDGk7hix3SosklnILf3rYQ+RcQe
EIZgms64Hw6p3vLryydOYajtZ1NsLQosr/jNbGthasXG1JTBVUB4mM0GmLOKU5e2J9Cg76L895tT
hz/VjiH4A3/NXTeZjTJrnyUjTHldYxX+9W1S/99DqU7/GvfUb5NjRuV28mwqUSaXUt1X+QRkSYIf
IbTvIvK133FASuZf1RZCE8yr8hY7BJN13bPPmfz5pqP+elq5+3dy22ycuPenVrbGGYhOUwRmhZh+
hPRUf/IIo/Cj74QjsdkCfGaSUit+O+e/Zny5K2VwgIspBWgCae92Y69SDWSbDo4FHUJ5+Q6Rrlnh
4h4u9WoCQk95Y8vPCKBZEjpxUQdhGYpl1L5bf5UJe0NQyh1ib02XaCgKJzBOh8TPMSHpS5fJSL8w
d4J6TgWORAmzBu9nMZvXIWbWVdwSU0bxsuG4i4EttdB3gSaq7aCmyc9X7cjCGJqpp92iWRNK7xrl
lubnQZjwi5Wb8KnNKuEEDb05G1HapuIzdXBjrVlqGMpsRLujk+Oivakdb11J3rngUo/CtfcQy6a0
e1dNC1eGI4+lxevrgkzJcRgMr5jP66nRMZPexqfr8ZBkaWd2X7scms+JxTR7qf7jDMr42BGGoNIi
fqf5DmbiyPQrWtP9ovQlTu89nd+djFCYvpE5AwebFoDNZArEWZBoEvvSBqKucqwfQ+x5c7y1tt92
pgZVe1bMcHFoEuPjYrynAe3T9sN6JKl2wNpOxqG5pHus2ehoECurOhPD+fJnQKOmRMR2j2tPPl2E
9fmrh49+OwgjashnhQitURHDIqTbeDUMsIVi2/IxQg1B0Q7Lral3RLnFTALiVP3GMY5m/f89gF3/
hMMl07nCrCbKlQq3UCtxZA7vzzza9Dl6o0IgIjQNSJZD4ZI30wa7SQxLfGNkzlpexzT1XeQOulBB
KbfZixe6bElbtDzT2DxIaN2HyAOlqy/fd3zSaPuCR4A0c9weVBbNynBLfNn3godN3SXejdp0unGq
wJTLcJb8VNSvmPhnEL0HHYhqqL4kc2gL+JLQnIcSmhr/1sYnwld03Om/DaYD7g8qHhZxMQJ3U/Rx
opw6V9AF4jCG+yqMmub5pDbnBEIYPLhzN2H3ziKaFDNz6tR44IWwB9Qn+Q11y3iX2P7X5HUGzn5Y
hqZKu1rXU6knCgOHLjnyKhCwvpALnpUfxcnepGt9DL+eS6fwjRgyHnddqf8JpB0nCGYMQ2Lan6fH
hZnXDScTSJw8hGDVePBJ/nVYSBIKkeQkKTmR5LYQs3vebqvLX2kQ2WcMVBX/OQQ3D1NRE50LB0Pw
AV8gNZM5akbxF/7QvE2RczfocV3pps/nI4U4DFjWBw87iUzczj1jjGuIzeidqjmB73PG4QPwUOME
BiplxdYkrwiCQ8zxvsogUcjqlVT4ytq+zfnqOGWFHyKSzykHp6o7DhjBJgkL2iu9V/+s6AU/BTp4
/ap+q4LYtAYXzxE7QCsw0Xz+9YsYIkMycH/46zC/wxGOGdKiov0jInvoHOviWvVNFIkjBVz1vSdZ
CpTB/dQKs5kgS43Ok1j5xyb4L1JBzt8jJ69BbhSBz5azUE1RGVCEcWSu6eh1CdmgwDcaHwjgTMeG
KKt98g4E3cPeBDYmGvD6EIcBDTEEuOJFUJ+JmRjh5Mx29BpNApI5poARiAGbYapTmtISzkxp9pML
4XTCCjEb1v0wZp5JcmSZfqR6m9rQnW8zZpajGgKn+krbEltTYIa+GwUkFL3bqpQgvqkbkpKl8zmc
QI4n+ayVQ5Qnx874wAFCKkiEhtKXuA7V8KAgeo/ckkcrT9rvXVC0ft6lCrqOnWcWz0x4EvqqxN5l
EuqWIDCmM5mDc+RvZuhQ+vEvG1ukXOPs8l8MKKiapVeI4AcHnHHlQ/lc8+u4OrSN63jPsn/xRndT
KzmbZjxEDnq7snJqh+bcIu9fznScttQffDjyRL0kI2AFWmDL2s/qg2EHYslhKWQeC8GyZAf32rZO
WSPKAgTa5hmtE1p+47jCsdhdKW1527UDqKpM/l1uCic6fdoj+vpCvUNKRPWS+neCtYvEWAGj0PrU
dE1R74E2Pljw5n2ADuGBoVsFKxU6XQ+rmIq2SvQ2oZvQUECOg7ihO5pgO7KmmBKDXtY8ZxSxi780
xpp3RHYIyOVNt1bBvQfMjhyvjiwz5L+cmgKjWlKlZ2Tt1DM3in2HAOglo5YPLmSPexpFkwlv8bln
wnax8DrOxYT25IiR4OeaJpziWiVbEGQ6fUb7DLsdXiCsfm5cdlNhLGSMep4fLlLK3DIT2Yt9pvUT
BwG7aJzULRlzuCWOB1/2vjDdeMx5OaT+JYkxJiGpSr0eX6qB31Vi7HEmzkMNvbuNG03uQCr1MBo1
f4sgZQT2P5ChHN15/l74aGdFq+PE2xEUf/fFN1bTKas5OSz0zcPrfdcDt2IHvFAoqrm3KVP4rd2j
qSHvHc6uyrwWwx2w3kux745COiaxBGxAexnPb4BKRxhX7n59OMAlI54laARzSPX2v0nyO4QBh9Gb
d8sQkGLZve2QxvkNUNGaVdblj3ioWypJpP8j62eCVOb3EFRT87N9oER4hEh7ZHNAC7A2Z/9y4xFD
FHGWR/ZKEgD8GwLlWwT4i+YbJRl2Tn7JtAGXX8jFWywqFUmckKxnyHT5aYpre5Tij8QRLobMR/iV
XFSWP6kYXT/ThpriryXiVKivY+ZKP5THS6fuxQwHPVHgs5LWtmO7pPYhQdCizKEt2uFLa9rWQ9v0
a12SOVH2TXpnQYv3K7zEYVjjcdsfkBq9L2akNap5Gxnmhkf38tAHNy5KQUBe9K5WKParV5+/o30u
PCOVsP9PJccysjkcJz7EQLTofoC4wkKHfpnSZyC13vRam7g6AmhbOirWTJ7mO79o1sggKRp8XkYb
aAwbJdrxUQzrTzyHq5mCY42FqTjtPJYgdqvbDCWGnt1uAsmxHbSZzik+ije/+lEor03pl7dSRgM/
FRvHrHh8iAgGQjSwJaHKIHFHeAT2cd0NRumOXx30JGMOJY0uz4EN6H043EX7QBjrVKhA8oj8UiNU
w1WZUSqsbu4EDJuKvKi0tqulXc9inPkV2tJafmKm+qDdJaygT2juEJh304w55cPxaowi3vQ9jUY/
aq0GXfQU5nruB5OhB0//G8ADL4JJkoQZL2k66tIBEofUYYD79rT/4sE4kMvE17jnKzjfUPtf5jAB
aWa7kvPm+U0S1BTPFFfNTApIr+HNuShTojGZNZCkf4oLwf30Aj3+bNCbzZngEnAf1ob/gHXPnbgx
TOde2mfbsdWFQeaHwFFW1vp4wZjd6+rh8BB7XFiiSGtvuZ4c5UygY54FzFoOeLgL/TXvLJESjs6I
B9RbkZUzppnm5EZr7KHoWeQIUYqPTO6KqjdgUJvF0udpPmbUJzxia0wunuegCbSGzYL13XGjY+h2
1LYDTw+nt12o2VNgPNq699NitjhbbW2o4O2lZg7h/gbBD5Gc0Oj8C5VZE7mWRJQulC1391juctXT
RBJV+1nvWc4dKH1QlqdXAWHSzjoK+gxt5BoxpbWb/8cwqIp/OjpCnVd0lBp+fQo5dKig/6equLTx
dX6/jZwWjgZNnPoPJcURSPCBiy6nTBDxeuwyV+Gpux4aRcui5r7M6yApSn4hcuWZblOaYnqh2nam
v18Rdtvwde4+Uw7vF1C+z2AvkTDMeTFzSMIQcT76xY3qy4aTPJHTC7mebop5fTI7nNVqll45yxZ7
GXWtK4JrfuSvQiQ3FWMBVCRD+TvB4TnAha4TO7sqEst3GTpDB8D0FK+Vccf36mOX2ovtOex27sJZ
3yZFPwK62mGWf91/VVFDTJ0a7wsZLzjMAAm8aelhJ5ub7EUT7Bq2xnM8CP4Pl/VK/Ii78A7Bqdwq
jg+mMS55WwNkQMLzz1EUfKAThs2XqyRi/7nZ6/ES0qJINOzRx8yYJTkUJeHRbFWOhpZflir9ON2z
+em/G1SIURGoOneYuX5s3SHQrKeaaqIKZmRdwRnpCamcFRhZb9bt4QWL4O5QKDiC2GWVWotHjuSP
fbe9H4rmMFgUvhdm5BtYoEGOkPZ/qrpsO/s7drAXYrEPdmOLLwSs2WhlZ+jOCEnwvaMedcv7W81S
18BYAnum8hEQgAPmdKraTfzlfMAVndViUbIghbUGcpc0+AI5tUqGcQsxL7zYUt/bxJ6GJUoESuIg
Xd9y+y7KlAYiZwEUAMGD3yJhDG5MiMiU7Rd/8FPpsficMpbFblGhN158HiyyAI7pAMwcQYn0vv1N
lpqmKKnVvjldT2yx/A4Vt463oLpemlZqiU9Trx1jiwPH10on1RThHFgO2OrjLLaGUhe333uDyVMG
LvhNnhR5ObrWkOsOBhPMLUTmS2H2Z8rI7fLFHBmUwhxL99PobCDIBMJF3RX+NQ3Eu8r4S+mqTzjA
Q0qX6EB14P3XzK1lE8WcE6lAXTZgTIddfloan8vFyA57Fgnk0EnW8hUu6mczIEJdB45WfYpRIPhK
trZKw3K9V10rK083X9n/hC7ubvrq+Paajilpbycl2RXXTmwdF/8dSfe2JmLig5RDT+5qGtfP31Bt
DR3vkAJ/6kCL7OARAroiwJ0fNKrGfY6SKNf6XFFB683x3zByB3/sxhoTs24no9oRhr5+THHFE29q
4oP1eSoM/BGRoT1JLkS7xr/5MZFt0ggWgnT8MdCdYfknZA65yHy7hHIJErIsiB454TRHsLrWkw8j
JAQVg5QUXv9MeGNQ2PRcTKa4kCjb5LAICwwq41l9+euXjtiOuMAvSxx4SRMalvuFb9Gmz88drN61
0++OKNu6Uq7awOXY/a7fRvYABANBlQgReLyolS+XFmK5MWhxB7Vcf2TN3CXUM4WyqBvaXltfsNox
cpirglkqYJ2MoFovygQu+WVJ+iPm9TehBfrDe7L+n6yp6XOdF5eyRX5WUO+5xBOpPd7iX8e6ADZJ
N9z1jkcaByECci3yovLdcp04nKtqkbx6lEdCGq4RRlSlZv5hZChUKcvln3DVwxnI4gpThEGX81Bb
qVxO4LusWwzOcPO37n2T1h4QvZ+gyfbsQ5/UhqOZoJXtOxPEwYJuhOdnhoT8HUYfvNFFAeFJNCyM
PGNfiGhGl47yzYre/AZOojcRj5WDcwuy8UYC9n4P753yQMT0jx5n5nC9R7XH+FcgzHYg0o/LYYki
I95PAIOuoiz0SckBaPCTVKL67Sd0BMibjz8jYeHRgMpOhRkYyE2CdbgBjBywPaXi7s5qR4vrZx+G
0Lx5sVzJnDtq5Nvrh3LzizmNpLRY9SGRsiNnsk6uo59mf1iKAYlek51q2FG7A82QIk8bYObnEwNH
lif8zKfEmjrDS+aMlPgrSloAI7c7n2U1+s8jovRVmRlGTgyRU4Qt7C29A2XwYG8GDz4+Np1/dIjd
2w5BdH7K7kNpL7AlT0vttiT6mtdisz5Racgh8aF+MncAGPNI/7UVfWesuobzpIg+TCKSxuNV/rpr
wT2LoTbP+ZtL4eiyzYbxdSqxmnoRdtke5VItNVb6uaIRWnu/s9RD+0JFCayUISQu+1Q9RZT0itFr
8bkCCeLqOrjz20Z1yj8MaPQ0pfdl5fe5lOKf3exjXFdzRJdd2ZUZKruLmIkZ47gH1NLNnayObD14
tp7iIARCi/4DIa3p70xkB/ZnKlGLGn37q3Mm/YXE+5E+uoVlb1Em+qY51whiW+clDX+5lYMPaV0U
RomUM+3f7nXN/CMVV4daAJouy2ecXNyNgzBYp2irtEMj9JXkvkFwONsuIsm5FqTRlBf0zl59A9Km
KtIvWa/kqfeGb6dEIdnEamTaLDGHQfHtnKt33YSvLIg6NTG5P15BgvSv8ZHwSW5kZnmmop8p/o7T
Us68ienYTYOm1YYnVR+8ZQRiNVW5G0vgloPOIajGNm0lP9Sovjz4wvof2XfqFO/s30BX3S61x5FS
U9WJTFvm2gWLy7rYUsxCr+UPsdM44es2mKpLpxv9c9zBVrB8k9x62dAlzXC8SdxemamBjoAqhglm
Tn9zwqjFQ/QWnfHjd8LrzLujwdv3L2I+XEsV3kHOwgD7dAUrETdu6izvsvnpWZOLDf2zow/FLxd6
AafUcEENPSavMGCZXBQK363DbiWzQTig4oXxWU0ro8C0C6hcDX4eNeeaJmpA91ew0YH2m4Qo14of
dcentm3q4M2EGJtrAuhgsxm5R6bDG0voPQkCkz9H6bJgs1Rb6PRzmQrXy9Sf94CRI+x+GwFlCu1a
SWhOWEf32UzC6/tfsu2MC4WX0g5sL93Wu7f8N1t99Og7D7E4YNoRaSZcwy4DGIbvHKLO6nw2SmcF
Xjh179AqCC5AScsvt95ndD184rSiVwwbQzN0cy9lGNgUgsbgIsYopBE+wXhNJvXcPKU1Ja982xq6
scMMq+1IZE7ef+YypfsDMscCeMmZXxPWSfuGaEWRe/8KmRIg3P7YSt5Jn6JEHv6BQ3kYNDtbtu4r
7Ozb9IeF0sgqi4dfF9jzjBXepru9wgCaGZN6IZvsrZWvssCLXKLSOuARxg9vcObpAgVPUYSeA8rk
yKRjrG31C/PpaswIrSctwEkwVHN7H/yJs7KWYCX2uvjBYlsZS9lz5S8yf4520TOcJX+qhMI0ySdv
TK7deOofmCZ46SZSHd5mglz23EP5asb1RHlsvrVgebXgY6zL++lxSlfqJX9GK6SBxhpKPc9LrVJr
iuXIUFEAzcy+C/IkBQQK7oc7gqAVXHUrz1fotX1/P1u4CAL3QJZHMVyFWyN+EYlWCtdZY/ZwbU2e
XCqL2p++NI9is7cYzJ3upy6eK4+IA4bWlw+XnpRMZcB8HN+oZSvdjvP3uioDeXWL5NbZmnpTmcX9
WmkbQl6tlNq+BLF+itIdAtMLjF5czPDCqj52/R75ZuiPXhLORm5uhjNYeQ1oS6+czmEvLMpfN/bi
OvDxa2HOHAYBIYo/w2dV/6F6YqLyee9lmJtyBEd+6XymOsfo+Hsns2YYIaVdRxJfRYEVmAgeqMI0
Cu87azv/+zRuPLm6+ar67DPhHwHOqfxuuB4SYdabvVWVioRj36jagBF3PDIaMXwgBW7Spw1Nploq
y6Q9zsfNTvsYkJd1eias8GzUhToKHVyYaqmHaCSlU6UJAaAaHrU/hnOw0emO07I53BBWmsXNpc/5
/dYO0z95xN5UrFOBx14V9ZBCgPJ3u6zzQRWJbqVyn43SV6R4bJChuxJORegByssX7PSXO1Hrol0n
nbD3J9TVhZLdpmTNkpB4CNcH2YM2lZVnIeLCGuYU2Lpxe0XtgM15PXA/+XYcl234pLtHUm25MUg8
9JO6X+cnTsLYn93yHfsfhrt/+1B5f2k8gKX7B0Jy/O8onxX7Tw+dLZAY82HRKk/5A5PITMZBZ76N
uPok/mXFepyPhTF1CcrnthaqrwX3VLPiznUMBo051BycxF/FmArLvEqx/bhWokit+9jBDGeD7KIf
j9WYpe+m0aZ8QYbsEF/PCs63NaL6mDoxFV3cyrKqT/l86rWTcaI4EimGyAomDL1/JMnRD297Vkrq
zsVbRUb2nY2ui+HFyefLkK91kpri2uYa2YgyCjSMRZjporWz8YHYGkjCmPFTMlh/SeAmkQkWTbmz
E4HzmOru9wdQJY2OjHiJ7qvILqDXuzAEpxZw3rnazbdJOpUiu2U6AMVGgIYWUbLObnMbZZfxVQJI
6d236EisVaagIK2aR4gAcR+QEiv1MXuFpqzL/iD6V/ig5qEY6wU7DUEbz6PjKARu/8Ssew9hPgOc
b+noi9biHHtPAbQi/VfJp6jMtOr9JA9jWW3+FvLuEdYy3/KTUGTSJj7PT/9MCnANy3nJbO+IOb72
w8W+WKZplFLsxKgkbNcC2t/8CckzQt+jmzbzkpbX74iA04tu1h2BdZpl5ZFSxllR10xH6pLgueL7
fIggXSy9RX1ROkf+yyqO84ZZ0XYrg+ExV83KpfXBr+xknXLGLVxI/N/QxVOab4PjkY+lE0MhDWkD
ybNXXInhAGQRvfNY68IR9bywJjzIImNWVtP/nY9xS6Z+EFxPAL9SRe9DxZExwUPqwsNSTsIszxxz
N4LPHf2PvkEokTZ2fOKGTHgtkuuCJ0OQEFn8dSEALvbDt7Jp4h2rzNo3yVGma0XEujIfUZJ9zcyQ
WJaKtFBWIeluGpTDXHKFdZEqg9O7brW3cdJ6TrCAXpn5qzcZVgC365tOInqoZxc5LRbNrgJvbuOJ
BYGuI0GLP7H3Em8pJ42LioyJ6jnke7aQ5HD7sizuDfFIDuowcfgdSGzDz3ynNPZHywWhGoqiU8VT
sDjBtfcTOPmILu9ICa6xKQKhuEeGMxwJiKM4ebfnUXFmr8R20zCYKeVpaJKe58jpWlCQ0gLmecws
2oL1Krszs9KvKU2Z5Ry2tWc0jLTV2zYsEUx9zF5vYzCfmOiTMJJLgdv4FjKnuEC9Z2sFlfTYkNKI
VHmUsx8PnAHFTocLjZETapMzIIlKwHK8FsRvaWEa8tCoQDsfEbxbDsr0zMSjA/Qys4U0NKikV+kx
zL+2/Cn7pYuE7VwiMV6/bz0iOgEyjUG+cRMhCLKA1uJC2lpVupk0M5dOFYlDaZo6h18mPrCshalC
oP6pZgG8lPM2E5RtqOHz57za1FXU2KU5IpqheTJxL0hYkj2EWBkN4pufp0UDYfRgln89/mOwXf31
P8qkJZvU1fSSTM9OZ/fejqD6l4pLOOFkqOPFIcZCIP0p8VG7vY7q96pdJOiHMyKUjPRWw+zvfX8E
6vkkxVOmWGioQFW61yLKs1yhJE3u9gMwuwMgqqpUO36NQZsv8/HKT6nyX4Z4LfNStfnnL8iLKj09
TqZSg+C3mgJPK/W4xIzmyg8yM1MREjx4LWYM2LINaLJ0mqEIQmoTOHEJE7VGJrmeaiS8ZFPt73Cl
SxpOMuZJlX9otek1u8vt3/OGzsqOuJ6K5N7iS1BheRrntte/iZj4Y1aBMcWI8LXUD2ZaEocNNlOk
HYhTrsOQygY1/CTgvqKFKVpSatSxQQYzSUBNacxGHQOro1/oyCxlDHk2JzxwRoPAexifCRfZkXmL
BaLC04c+Qk5q9kT3ad02w3I1unbhj4xMxCiIsDpQ9JaHFnJp9ZyJjDdxTyW51ct4jUGdRPeOF2XA
qEcyZgd7VD9r9WUak39rUqBvF8M7fCPM5ptj84uW8/QP+noXZyLbeJRGMz+Xy7xaQs/3KsyYu7eE
mzSbHwOhel2lgdzNRy2/M5Yx1RHPwIyzeFX6Sd2Jj/7bwP0nsuON25f6vWIsb7/fOzG/nmadKkxt
xfWj9CGB4psQZu2nNForerx2sdKJJZNmnGW+JMwqwU2DUX8wWQe2aaAMVODsC3ONX/S03/ex959j
mxF7xb+C3YapqzrMvy5Ftw0UHHTd9/E9WZ8Tmi++jYi9iP1VGxRbK6hXUCFTPRSwyLesHms/pGH1
keEpfieR0nxcAViPUmjZhqNPmtM/ONuYqntFvQJNWwvXgV/YNT3aCHs8q8v5wtawwSLxlBxW+nbA
Q3hyBZTAQGHcgC5qF7NvZ4Unrp+3ARczPKWjHUQhccBTKpCsYeeg2ni3X41joOSLUbQqgiFik5FR
Aswy+S9H145d+2MXY0TL/daUcu9XLbdHdIZ+yJBUrI/KruTXpmRLFlS/BNdBBX8cR2iWTbxELc9G
lqeI1gEpbCgd0MKf6cfGBAliLYucIqFeAs5lY2Ml7YIqH7bFpk+WbsvYm5cNoPld2+icKVVkJUL7
HwOSErEFgajepBiFwvFRzBh1KrGRPakXnja71/J9sBzZimWL3l9zbPuI+4F0TBmJDLGX63thW638
pSeIz161UJmci3zo2Y3UXF+8Ebkt46Uokf7XW1HiWc7LSt3fe9KybT6VVp0UsQRDJARWpZA5CqBR
2q2LXzRMCYx6BINWv3MGp/z60AsDxDLbIwasSMKKD9CrlvcuidtK0ZDLRdbYtMgOrmdE6I5bg9Yk
i5t2oOv9tP0XpYpsb1NxgWqCQ2Wc32+iaEQSwEG8GXuSlwBh+Y9Af+LVyw8uUggmPU51jab6O7eD
dDXoETTWJnvkqQ7L3oCqjNA0bUnu3kXXF6kM4n3dqyAFXujmYY9VlvQMWdOVTn0jpGJnWOD8+XSJ
CaeTYpEwXfqJwQX9qUV65Fuu+dn3ilVj4MF2+O1ykBKy7g2x0OegPRWH+ww85o6FW+qBD50jO55F
JUovv6puReD7ugGNUL4aCQRY8kJ3Vyx+4j9Ee5Um6V1cWD//X0h42CSmVhEMpbA9/InV6TDnVW9M
HqsOt+HlH+g70QRkrDJXMvNpvIYqU9GFLW3h5ub4GiK0qIj7yNo1bcNEqn2nJBJyg8dDjC4/dJ8e
8+nTI9HtRfHD8YlET9PopznojH1OayCp1HyVIHOK+kcrV5aCG+v7lFbfYLy2b2fQGuqCeBd+IIRG
/7Ez7bOcwWV18kF4BRJ7guUCn/Q2hAXd8RRCu4avOuDnbTwAOnaSqNL7m7J9dBuTi/b2ajCvuAYF
flfAZQjcv82P9bp8b8eVjWqsii0KLR+hpCHXAKlJoKwzT8fVTPBcx5zGznKhAvkA8EEm0SabnelX
eIEY3nhuOfEJ5x6jaMtl70F6giRMe3eusN6RFn+IfeT5nhmrO843L2TVeE8OIaWchAIRbfTXAQO/
3lPpsjQ+JgxkvBsxp+hB2R+cwLIdf9LOspk/JWVzecLiGDIw99VLS1AFx4TMhus00bRqiw2v5PX6
+4nbZOx1jz5IbSEW61eVJwKABCXfKcBzJqHCsknVY4P56AFGHYWO4vYVdz+2En9DubFemgDbLe0F
ZSFDkGItAvqUicCnXzl0Wa/7zZ9OUYTBEP2Q4Nyrb2VjF3fJkLalInYEUrt2jAsNRfCez3t9+4Xu
4SjwFCgF01fLYQmIivu0AB8CbJy2bc8TE12uU5xKZLii9N1rc7DTDfxui9aaFyag7PwtYccvLP5y
OaCoSGNQU8KlPTUPxngFTXbqjQNSoPw7YCTCnO8PQSge//jJ56HVNp0VykF9xT5DbKH30WqWXECC
f3Bi9yllgf+4MCgazPn5BiTHRDHsRB+RC9jN9QqBSkjkM9gvpEjM10DpsQypwJe/7TV3aFVj5I6s
7COTdmhZ9G3vOt+vqf+6tustqgSVuhXj+2u7G7OSHKWM4a46N4VqxarkREgMngeuSg5z4H+5XK61
FLXBBLxBFWv64yH+kOV8nPfVLKmqwOz7Re4Us071QU6LW65vpimpzZjxMymYHhMSqJEKLJbUDt5v
TJGJbCD7Kj/rrtKAcEqoTWDFk7L/JJkBqi0IQ0+Fwvf8l9qZnoIx/nBRmJaUBq9ErLlw8SyA5XJg
gM008u/BOkn1+N6jcsdNKOvxPIaCJdEwW3qn2kiRXrgSZSdrljLL+kj2X083GEmTfJv7GSO0iotY
68FINx08IC5qctNU68cWw1W1e6h84qyB00SOCFgXNW/E3ME7/EvjfvNpIAAtPYQBCu28atfQ7D0E
Cof8oy9NeqjEGi/NCWBsylWvvoThKumim3zxPnTGzpFi9TjzqABfiyxuFqmqEXwbRllnlJqGLefe
XAYzJJnwNwXIuIo+YhisMLzaOm0P+AlYKf8bqadHum0a2ca86ueZa3h8hM1z8SwpPfmp6P3j6RRT
gSVmcy18wSsO/SzCBgm0ls+mazyrKwRxDZWqYo6Egv5yvf3KsHj7dG+5PGK8Nuj9oyJ9K0wpWJWi
yanIVs9KKeUD8Nwy9jlc5EuY8nHbFzK6jVVGouZXgsrAY56gRRqEg5REmHqUBtlTRweQ/7Oj8pa9
Zmi3X2FJFTRQIz0j5Zu+6R2WLkd2F0r8MUCkQwPOAdglxxJMQWJGx/Zk2H1gQHo3nkluiBNaF9Li
BTd6UVgw46ehTn7mCFoPoGt5g25G2z5US/n5w6wHND11s+EYDk1o6QJjVMcLrMMhES4enZLPeRmg
s01I2q4Y4T9khjIiLhcxn13v8m2k1X5f3wzgUBcuKkzS6iZkgBiKuhHTnG9NI8/FhLBMIZbl48Av
zHcUYTtyU5yC0x5Zb4QYQYdqU1sKGaoti08ndeG+8v6r4VQAvGYB1yxzqGSxcffn3sicdZKHlYjS
1mxhDa7SZ7NLfe59nZ9bLdUe8w2ZNcb6B5D8/h97MQ7lWJHSR9XwHsN8PcMskwJSzL0YhFcTvWbF
vhivG6rTHTsIkEnOjhjFHxBqxaNH1htBHS10COx2qg+Qiizr0i8FdcFhHcCbUIOpLaUQpckW+OMr
iDX1ySfSqlLiNVIh0YLL0HklO2Ur2+xZks2Wpg0JAV9Jy88ftu5ObUjctoNznbW74aufxRMD12N3
9OV9DmgPbYef+ebuskuYetR7uTH6To0MhsFbmbgHnDfSrFu41YDKUPKp2+bGaKPcC8x7otogxhat
60yGZIg89z9TX0Hq83KWb5pntxquhOYlpDXD2iVndNE6XpReVKlcgR1E8DQ1dmhQoqR7TNR6hhcx
n9cppbm2+sPhVnuqrsCnsm2o48x5J7HesPbdBwah5hszd8yRNwq1iUnVo0xOXpQwDrkmVWnOxr+I
inaYzJxvaYpoVMn8YoYLqIMBkfQ88JyKS2qfQyZw0bptrYVj1xyMQPxD25Fxd7mHPhdZwGjgc4qB
Bu++AqpJJgYgQTMSRON6pJGXk1GXG71iuqzs0nKRNRFIqTheZK2xHVK7JnnBmdhd7xEvR6RmRKmt
Q1nubYsMUgOrJu5k1Ct/S5kys/TOeE79pWZvKPTyKo6ETxCivukoq3sn+qcMbLP358e5iQe8TsG2
UNT1WyzVrKlvQchxPE4a3Ujpstzneh+dCx6PmWYDBWjpA/kIWjkXSNx/uQMvq7WT1QOQk4UXVxum
ruJxaxwtWs7cbknqiKUYFN0QMtIM8u4CrVgrFzfdCD9Q0mcMUy5oqGzLpWx1H+ND4IH1AKIUuChD
UvQixsWPGn+hieP88v1bB1o/DkwVNjI6f2VQHGTjyyNQPRlWgwqtpyNCONbL47n003IpC3pKKaDK
jbkmIFTedmeT/MpXeWs8b3/eDJxvME/cKgkPzMURZqItET+kucqakyMYkdZdiiZQRJrjyT/yIz0l
4vFbq2zkOThz5+4ZbU5mjlDZ/LdivNyj7P/YGo4dEKFYYWwgoVfAKvNbjLQzwMCHbTT2glUMO3Rk
IRpe876vi6DiAJoZjVKngqYVl5fp9M5mDrNLPzYypRvHMtJEBdZ7qRVX670Ay1T7K2r/s5qzfrYw
ohOZ+yMjN/I1btsUmg7OFnDRescxY8DvtKVrL85pmJO+1N7ZhldHR5fOwNUP9GAHgdhtDDSe+yLA
u+LV80ng/8mNr3WY+mx87pVXWTuPdkdeyWGx3aMfrkoH3yX7GPrfdjzTBFzj+JzlDjJ/wL1WV3Yk
soeQZ8zQql931PGyGnpoQVYUuc55McoGmRPNjX2noXBaJfaUIHdnStB/jXzt1aUWn2hanqzQxj0B
B16BWFoMyBKpxM9vL3G6Db4P6PaLNqxvz+WsttXkAXZTXYfSndNeMvBpDa0/ALqNvbkPCXJ/ROp/
AypaZwzKumnXbg7cvNrbtUUHSnSUgvUT8HqCs6uzooop0E38G+Re92xpjb7nGjFOaRYxAVyrTJW6
ixRhweqvcP19ut/HlVwBPF126MJXoHQ8wkhNZQB1nc5i9CD2UyMMuPCyGpOzcN8U4BsMsalalTTk
OE9tsF+LBPdcUx6JUChQnBIzNniaH+uWPFOfRFtBmpwRpS3EYHHIp/K8nme+ygwq7VlHSHYFclBB
nrdQ3H0b7KH5XUaddP1gdlHM+9gIVpRlUH2EzvWtA4ZNz2PIYMpEqLNYw4DUWRS4wt1Y7f/jmQWu
QmuhksHi+YcDdNwjDTVlIc+HljSSzk01HTFkwu2hm7JNETyC90DYzcw2hzMGTx+rX/7/O8gZMdo7
2dLsVnpoRgPyetcfMb+GR2GDfaYSH7flYaEV9R/WX7fjnJwNDjxibH9n/dEPbn4Do6vQrfm/9UHP
CxeyJD2dLbiM0SxuHZeeHjXEaPBsJUZZuEcS7v+zIR0lNH6lSb19NzHsCAXnmr3A6RqfiBRjNyIs
Ug8+IKJNtz+d9Q+JdsWtKYut4KyHQwcYB7WLPM4tlgj0HiEVULMeObpFsND4aq2DSqkgfdJk6CtI
DdpwiJyeRCbLwiAt5UBQ8MGkNPNJoyD1wlkO10glng2drlFmCKHOaWZ9gIUJOeIRHBrTFnJDDxE9
sc6Z7/iPK3sggjktEOizUoYs5bonJcrdZPnxT8tTnDjY64k5WRp8l4CmNnyhixj4hDrC/wg1ALDP
d7h731kwZ1DhjijBmbhdU4Cd2fSDi1IbH4XAoYMB3p/0sBV2FJ7ss07cdwfWPCWIYghQJ21hilHH
9ty7elIGXGsiOgJBoNSIcgbnlazJeBRrqEdHqtuqP7jQJu+vka78itWBtQIZ3xwLKpI+C0y719sc
WRDRTN7N408p+fsNLOBLkXdWzZKtG4juqQ6tJwqAJwu1RzPvjPaGsmsmDFqdpJl2YJKh+dXKk0co
or5TA7+jD/a3jtJZLolW/H/laz4nvlBCgRF/a+lp8J6/2+WkcU4kVX8iuIaMn5Hnt88FVY71MT3H
N/MGVO41HbCYOcbgtsMr7xVCO19vBqRbVZNkwF88cbl1mwzxplqXWRJIgiEb7hFSeeoKX2vBuMUc
k4Hc8/16f1fLqwDNddL8sYSJx8cUGk1rqh9r5nxV9wDWgQ95yxcMo15zfP3elWnTZRe56uGGVPHq
bDAdFIhqzDzNU0MDVttQIIIpD4dV34xEqrcYz8FvVscGvFfsAuCbvB2ZlVIWlJ5+MwXufRr/sjcA
3tGjmz9ZzS+QTXLuXoYJvHkf3UhbtJHLEHBHi1KlDdVy0irBnVvN7946t1xUIdhy0/9xb0xPuJ65
S50ds4pz0GTWyi+3x41c5zYBNy4Z34GlFPEoVhPrVil6CtmsfhpTIP9jyhfGxS+wjrNbKSgzdE4v
tTr4PrJku5DU0CWH6J5YrJTGPkOmUKcOyN4hKIpQmrAa1/sHxT6grT4WiZI8rLAPbu1F2HZdPHtB
D1CHtF684Uw5VuP34z6aWr0J07YPsG1HYLRYejOHCTgJQ4wlEXDZM9i2gaOCKTdRDZre5vvcFBUI
aNd4gp+dfqlBQ+GWUi2S1tW70mGWb6cFLnLebZ4MVMWMo4vo8fUmMIXwTwbdtWtyVLzevYyPGxtO
B8bLhJAEqSWy0UqDhCPnqI2QMd0UQqRuoY5mlisumKfS3Baodxczya3gK+bWUk7fNGczMpp/CRWn
kMgPFo/lNdF3mm1SNZSsh5DHoK/fPR/0aVPxevICSA3fKtZDR1XqF10uoZiq8sX4JKS4lMVvdJeU
xUBYnoqJYOMOxv0QzGYYGC7JdOJ3yL76YXAzomASzD5S3mhjTn5de+aNqwQQ6/NhcqL8fvKchndJ
tFmPVRznyCyxPp8djFQtRWWraT01PIS2vF9buY30v49vgDEcX/doJjzxoGGN5ic71Mm1h1/Yn9Uf
92lhQnyNYBQf4Ze/BnUbQ9b1fNS88yBsE0I4jCYEGRyOZORODL3q3I2nnq2FP3mxc9Z5irEEp/GL
8/emJCcDM0bNFoXQOnvi0fQEKwNc9cC9nm9JRczitbHC97e6DaFSRD7lQysvtDSFQNQtu7uZTLVJ
e4c57KEQhebnBou3AQ4RPpNfnyFLJrieHqRSxRaYNfsn253xt5XSCi9Q1R0j2Voxdj4Au4CjgoKy
C/0heLXFL4F0JstxdlQFDOhJ5qCbxk4oJKivq66wEcDVTGJGuzImNIF4CDXQtj9fG0qHQOQqvnFi
HYvKsGlgm+bhwTgfcZt4BidW6KevF8gy3WFbYNOCph+bApiEfVOqEWlr4CkONTRcGCT+U3lDYoVh
N+AxYtNv8uS/+tea4rmg56EyS6njlHP2Y2YVoKllqwO5xB7oPt86+W2Z3nv3nZbmWK9/oSJMstib
Z24F62L5T4Q62UUYd+8tJQfMcokTrcIuIWdDJN5nhsEFPvaRYCoexsR7oPLYxDsM7OMAWONqwW12
NFo8XrMcVn04BtN4OnMiYBaxHYV4jPl+3eN8otgPvVdngzywBXYT7sGWU79BE5z5v2YFeHAnXHq5
ep/ugy/+bhmc1zwewNxvsg7GBZwMxwOSCT5nzrNx56EoXrYXOazV2YxYZOCUhmPJI3mS3qTOyPaD
rHuvndJFUX+cX1Ce6DkgIyLiGS0EwaffArsTM799i6Z2NY2MiiBVkW0A/3J5J3As8ytKagk1Oqwq
O96sddEiK9w7UU2/nD0RwKDC7elh3TKI4JAFahTw/liYQIIuTNJ2g+ZLgE17JYg3eb1yXscZrN+9
bO+WW6OopP9HPR5YZrOt+M/4o5NP82GxdhFXNw1XwSGbSJ0aYVo3SJHFNAiYS+KBrHQSOj58p5tI
2y1GJ0cXvW2CaJuVvfSLcmYCcQkSRfEgNTJbAcNbCQ1El/p41VFM9lhKkaV1s41+xWs1/SRj4XoW
DiqNLX0TA7O47Hvn4VHXhAkjnpLErt8Ld+3EGUYOAuuU1ocHlf7/TEPUaSKZTTcKQEpcBaACgQKt
+PTkOwFphb+dhOXorRCEwx9xt0+rbE7WUqdICdbGOId41Pj1//pJObaWbWUKzXvU+CN1cJ259ntL
kiXK5N8AR5Tbz2VCKZvQ/hfYwSC44bsVWnotitCTg52g6bEyE3QUhUYjG038qNzWqlOCtvG7llOm
HsFfF1CkyhRcdclkCFjdcxh2nU/SLEh0m7MjUe0dwqvewv05S2v5I6cXo6ndkMHLfeKo2V+dYCkj
fjigo+3p+83HYZzM/xtljXf/XfuoBJO+BUjEcGDsdojpao+cviZqOe72lrheLNwnRMy13pqUPr/a
498qqa3BFtjEgQaJ6hHC6f6HFlwvnF2r9E00M3lfoh+uXJzhxqaoq8w/g3skpnBfX8YhQVzTA1SJ
8MMRUGfwrdEnSRZYBH/milZsqGL2G1g1le+EIHtJbqbSxTD88laqrK+wlI9Fy7l3qq2RLfqMtf5O
UF4njg7FNzJlrKLU/lsBH2sc98U35N8hOqaAvVJsVmC0/UPusi46wSA282YzC1klWr/Whj7qJGFD
3RbEAWfR4/pp1Z5QCsfqCm+DxB5znwEdG+ZdEMCpxHradX6RQrH0Igt/f/xlZejVCjpOYoMv9/n3
pWLhyQ8eorZUDMwPmfcZikZNYewZR+X/A3hAKoJpADESI+RBOZZdlb3r/Q1UY01tRw1gDVbhk+Vl
teK8i0mn063OtHAxM9L+cIEMtsuybV9MAolMMACi1Xs137VLRcgl5/scgGZdRzTNS4cSW4/datiw
UbxdrJgUUVmxyAQfZyRrKCEcmKBmudapyumyy6Jioil1+LOvzZdfOv+BEvpjlyWs301lbAdcyEsJ
uIE8tyU56ihmVNJxw/0KCQWt+lYb1wmN4QFdoiX2QS3J8OEveAqOVCrtrLoB0chqNI2uLnGnnXTg
qAdPIZEScqZlws0R+YOumOjjiIrPb3a45moSWIcVnm6S8Rem8LitauTi5wmJabxgYXPMVismxIW6
ueozYyDnWSR3r+HP84YEgBmYKUXMi73OoKwsIly1ZSVoA9m3zClWodRuvzkNm8UAg1thbRri2s9a
EySY47ON9uRmlCR26/wPyKTR1W8/87GWMB/mnWjKI1OqfBo0MXZfVTK7YVbTD3lWBCMW6l5AFPLp
VRkfAz0gLrHDHGcJitZkS9zRBpT364fXbAtalxX6wknHVwi7DfCH5gR2l/amrbwMOfSZ6XigNQgt
RCkxR5ctwaeEc4AGw12B7BeOOWEGd6bs2QLd9zdilxT4mY1PKiU9biy4G7WWmrHXP+NxQpHOx2W+
z+47d3+q/wnPeetj+3gp0PIBUijShaB2lEmS9nbRFaUBnX8QTq8SkclwrMfeuFrJ0SxvwfufXQuG
mJtMgU01ylVFUadNrhLdW1QM4clrMBwKBIa7/oEF7Evn3tpcY2RPjTP3cn+CuiCuUT5/p5kSpBmy
ACfQqu48WXz/ixh2zBTciQnLgtcvaYI1f4L8+pSk3oAMxJpFdSpV1TJ8zzrH8NWmNxkd+q/Yta+U
2nKLzAy/Ve4NuS+rsr28Mck7WgMXxj/+Ju7FigxPw5+Hzs8a19in+/ATtKChre/G98buWoWpPBEP
ml5PdR6rrm71KDpA+HojlS2OuZz/yiCuB0vQS6CsGgal8OvK1a5yrfDQYbCWlKsmOUnlGWQX3mqz
fEPOwIgzhYO6m14nhyJ3JXCuI8k+uI1tHkXb8YyAlM0McYzwv91nLWd/4qixmRggLCLrNapp/RYG
W22UVqr6HwTQKhsb6f4YFHG4mjlU7M+STYbL64cGHoJ1RSTDg31eKNdGPvIXjGM/D5PlkR0k/t1E
43a7idMoEaQnu1TS3s9b+s6sTelxc0h5akJAWKG1tUFSKGr9qFu9oy41tj4u22i8jQQcFg4D8lnC
KBOPWl7WxvnQSfwx3jt4roFzHienGg5Nm6eZY3dkrg7YmwTWSwGMEZD7VglvKYSjnOjjKZwQimFF
gMbzHSCI48O3SYc4R8DmiXxnGlUn3quVbo6Y+v09BtRZuz/Dsc6f5ElY0BwVMDqNXfHHkSlNYMnU
MaUH7o+LJoykGOw+dT0MCSDCaouECieBGfbmlBGsBfBNKg3YhaDpQRE4f49MM2O9pEMf+ld2ennW
0RZjzhFqnemuMbuDKFTgWZ47dUVIk6dMpKZt7o6D/rZXz8U7hA4a9zfPieYQO4f67s23yi0leOJk
2rk7xFuIc+wJk6Tt2UikPGZuZcP+oD9SLvlOYcKzTvyr2ZIYdvzLY6jz/bGStNKaX1LyhI8sLRGQ
aoIbD7YPoH05CUcSWhhiZJe24tYe5JfWGZIX5jtInwbJStgUp1MnlZmm73Mmf8IonvQO7PvoO2jz
N4EX9cOpHe/X9totMJsw0vyLW8caPLOJxqW8TVS15J5XWk6DT5Kk8VlcyHxu2jfYfntqjoO0AdDV
PSrXIm62iQlZPjCbK3aSGPmW/86EJRlF7gAG1JYHxYevejjrjL7YXKpAPeVIzrfMu/dSX8Wcg/jL
Mkt/c1WmxA9SmpeMvOX9Mo5faMLjxzWiY+4IYyKpD2NMGi6TYKKfRVKVHknf3dJhKxaLTHlo9jFs
nVXdttVL47ZembFGWYWq/Akiy0TG5nZhfhBalYg3/hk3p4BwSiNTKJtgfutxwxk9qsOikTmROR/x
O73ykKb1jWJ/nSUsv54KWKtokRuEeWET/4AB8WzhQ4MHySRCXlhaiKpcBwL+xZJbrPtZHT/8VJDN
RuXBu8JhuxzGknvz4uh4j0XDgrWtVoxQw5bIWGPuIjBSa4thdXviihpOYBu89IkbQJwtVy7tNtmL
iPgeSVTadb3J7xuq7Z9GCHDquSVjoHmUPzxFudn1EaE609pB1BuJLgcuxHeyOcMTrtaU8ycSrB6y
7hdYwaNKVEhneFr1H3aBM9VfylYsp2hhYg3h+yJML5mYljB4Pq6KSM1qFEEFIB9SIFtBNNTp2x7R
cxIXsKvQfpbRod12+gkX0Gimye/rhkf8gtwcrWdwb/tUob7Pn8QhBqgLnqv3685DisxOKG6Ey+Eh
KZL0vv3DGkeqsEtSzqBOgX6gqVNls5WIf5SnjQle/gdK0Bitkp9TWaP4N3Q3hhGdVGHWoLW6/U6q
DSRTcCJuoUe1Omp0lStwffGnCASes0wszjz81rM3IEayhGX02Meqmbtf5tpjd58ueknky+VpAO6O
2/BKPjce9m6c0nBFpsmBr4hcE4R2uIZXRezDQxp+Cc24Ex+7oCv58Vjd1NRIje+uJI5N9xDFWXnl
Pqw3/dMdhyqpInkdhO4EA/ysQe0J6J+wWjYMj/gpFg/9Fjl06vNF6mGtmnKvjx2/fgjqse7w9fTE
IZhkhizWQCl0omPIdtgOtoMRMcnwgBW+UQ4f7lIwB6Dq9J9z3mgZsLdj+M3+9eWj+2TMv4jjCgz5
dlcCInH7kYk9d3kYO8mG5ELUGs2sLv63gdbGHz3PzyIpoVM/M1TtruNR+4tdhmzRERzmXUtmr3vZ
cKN/LIIuVhY/D08NxperSMWlB9b2ciq7vmyqN4WGYBu9lA4URx+0hzjc9ryNrhaXnT6Ar6IQwQ3a
YXOP3q7FmoNUqtyztf/XhZExERqwhjGVsLvU39B1ldOmdXLNIezOCzcJB0kZ5XeGEXkgrx1gd3WL
+d03qMf1Mip/djBw5s+EXfnygsX+K7y4HzEbhqm+wgTqSjFxMRNIyu7y7fymCY5u+BABFImhyOt6
RJ/uAjC8F3eG+kMmK8LXiRvSkDbefoarkNl2x+ugkurZdKfX472y1Uug1jgj+uoSCXW8VSIAfSwu
E5mw1ENbd8tG3y1oIhhUUzSGFGigGEHC0KT3ccWGNOHncX/lc06E86qSRKmG7g80n98AnrRu1wjA
C3Dw9HEYjKyY4EdHTl2I3HOiSPzQMwnld3VRw5UCnZMwrCtgmOxc18Gga97fBFjTyT7Fj9yRs4sP
6NizykoFsCMYmwdS8db47x2VA7E1ZfEaX8fCzPpGxojlvlezjXkhgnuUr5lfiHyofF0lpxWnz0/T
A+v2nHnV55kK1TJI+Jmv8MAXN2CpxTKR8lAg7YnKcAkYePAQsQQDkpW4YQIFGXJ5ddIu0nBq3R6R
QYlJRlQrH/AqJ3BkLag9bxH1/+AA6PMzX7Vbr9QbFsLSh0Vxgs8geP+fujrbGaCanPrAcNb8VqKc
jD6MG325tcrmXfwaZx7uf8uJW9urP6+BUx6C8Nl1PYNODTQb4FGNDoQvwFIiPblcFzPG5Arjhvdi
iY51m9789GqEa+7Vt6sPpjHDjxlTyRBn2MuiTkd7TWROa40wyNCXOxHDkaJNYvTmPTFEvpxW3c27
MviZQjjySeP/WN8rCynmVqmqHqGNkONRfwl9iwg7PXc6qjmBF5Ru2hRSUTWuHBvmEKX9lcdju+CQ
1v5x9VWNXCX+Q4AD8E0QoHKa/HrtPFm1EIo5skzmZ5pSnitRrB++FdvuRE1Kw/j7tOklTmMFT6PD
Sh45a/f+ZbNk6pasXxKdBTIJMW5ZvymposFFeOc6hg0Cw6fNMBB2OT//UM4IcCDZFgP0ebtD+NJG
EqzzopT5yYuRYXBFh2TTxD4suu6yqHIoLX8PhgtzhxGxasGN5PNwxIfOtqy5hlGSUEWfCFJ1BRvs
mC1cwdkWQtn8tZk+cj5rM+xfGKaP0Rx+SkgKC+1d2EDJwU8AKtNq2JQyxdb1fiFv3EbZ8KKbgXXB
32iQDqIxkiK2QFPKLu/061HrFQBqDMbNuUWhaYIsGsLFYbv2A7w3mwWNAURVFHp+/4DbKVjTTuXn
ZPyXOZ2+tm2Q+Gj+MPMY+7y1y+T8j5+a3WEESGHaU07I+FTIzyV4UYOMxJhEWUw87OmdM0I1WKmF
MaNemMz9zFrQydod2uAjxqnO4VGJS2PmZGp9nvUcPfeYa5exK143wv+j9jK5YycQFHpfmRTrFyQX
8wBuVg65lnaazZ6flPGAE9seyIzJeorU3qMVrty35ptPPiA2FpNYfz3eLxlkDX7W5vJ7P5WhjIde
NyaWKIWvqe42M51Gsivj59fGtKuobe+3lPjIMYJXoYlw97ubKtcG2/guR3/Qi0WcbAQ5taaIFPdt
p50K7ZQIKQxTYy4ZH66mQFdrwUSviwRt2K790wOgG3wXa29MQj547rWsHhE5xY5qPw6Ci/NGa0AD
b+Yod5QzUtCho8ydNJSqEitm3oJFRPzmhvjqzJtqGprHftR6wbuSf4qp6F18BmIQJkzt8+AWOqA2
DabeBK0/+UNsvQ5/Eh7IHd2wPdUf2lrhZ/6d3CzaO/HUN1SwzyMXLOc2zwOIbHMY0R5RtdvlNNMa
xUgN97RmqoSMBWqvxk9l4SUmwgnljuVJF+gp63ia8MfzRmhmk/mWzKI8ODfu4E1H6v4geNmHuGPw
eCymfivBwu2bxShSqQ8B3Srde0Q510eVBDS793IF07G3V3goTrfD0KIFmitlWSUKqOzUyY9rUGI2
wlxcftwXBw+dU+W6gt1Ml232HWOVWUN7L6A5OZ2o4FafMnenC42Mou0rQa7T1k2zNIPXB1PWHyIL
0Qjhuc6dp/Ey8ZSGFYLWtUrpKmQx1XSvWzMnt2OcwzFa0uGjuNwfsqIuWYdtagF8YfFoiJ9CxSHT
dAZi7bVmeyKvkd7mDF+FPCGoxAA7bRkCfIKtuPGTXrKW+l/fGNMFK/e5V38GmjnbAk47JQ35nzwl
sri3T1OrBK28XlSeqR7DjszN4PPpzNhsn7byKU5BGnTetx9l02MyKV+wOkc9C74SzGyXjfv2Fa0O
/XMzSN8X272Pp9RUK8sd+hxv/OHn+9PX4R+JcnagXGELK23pdBZYwidfhqllfr8haR6jBhr7mdTV
1u0vaHktK/HjQwcSVSEqVscwGa3thuAowkFXZ6u0/sAI/ukVw6Krzu+vnJ73WygepPaYeyvjSh78
/xPXvK8LZD44Fvui4qIoHGx2ZtRGMquuppWHnhpnR6MjUKZidCKuOcYbowQLQh2DxC7MTBYAoxVZ
HGn2003sUkaGcJZrXsgxa6I1SfXUUvMnhSe0opW+jMZLK1F+yQAOF7wkbdnEb3byCedDxI66gjnw
vlxicYHvRRRXJBi4vThZJVBD8NRn8O2KiI15QdnBBFVQLrxXzlfocoPtSbJzk2Kclh5OWcBKK00F
SAzih+Z63AWzjJO8QK+GxPHaYkV41LnKfOP3hzOEvJNuWsS57PIPxbDSStbXqwNTTipEj2cYMGfn
dtDWVPKhAQa1ShmpMxQopJGY+Syfe5Zw5Y7/pYSAfTbNk778mrjFbGQSzF3mWH5hatQZCcQL8gB0
K92NQfG6yUxSx9dDZRZ91/pvl5iRIRte7/vgccV71+FB8KtmsTviLNzTXx3xt+rUrwJohHqX71r4
jgdmr5pdyNTREsiNJ3/vcqJLnQyKXHnboTindu4J6N+zsQ6eJQznXAAdNBU+NIIxcOSMEwVE76JU
Q9V0n7wf9y5r++4uo9W1tzf63UqKamQzDMGGtr9bdPxmtJlSeng9PhnsukigwqdlZ99irh1dX3UN
uoHxfKjIlRGQBebJ0cZ3/hhhzLu8OAyFCrmknNURwK5nAVwC0AUaG8yP6bdDw9xHREE1SBd7Rcne
WsMaaOAzgIDaGlw2uKU0vAWoiME8xypZKnsyjjDT+TTQE82uD3vnTBosrNy8YaGkWnhTyhf6Qaiz
yPxdhZ7083BtCGfr6KUbLAAfgZObh4A/Usz0OzmUbUWziSg0j2vdYhOubHOiAWT1aBIjXDWldORX
nZNpOJQNIwIRcClBRVrC6uTYjwb9KF73mIl50I1aPZlVWfV2uCfYw6Hg9edRrb3/mhiJFlKAIj18
2mHvTbc/XCywwoDzvkRPpEniNCY0Yr0pZFZHnW+N7NAdBDKh37sEsST3EE4sGr4J9b7dkGEs5Q23
u6jc1KoxK9jf46zViFRCbo5aOB/d6vOujmNXd4JPfq4jZBKFB5fHlk0OL+SxvxoDcHgsArEQrqbH
R/W6N/ob49Ap3jC2miYRVF97RyMSx9mCW1YDAzRmwuB9cuMDCzb4dHLz8Io8lThKrsaAUxwbdDJZ
PLmfhOw3HBJuOjg/HbvkgP/2RemoFp1Jn2GrHjStG955pPO3Vt+2axA1JCI3K8WNxF4X4IVQYLld
lSjEtRn1gPcCrwdcLYHODqa5plg3V3xKqX3neoqsdsya8ZWy8Fk2X4PsHLBbPUgUAtg+vv+0Xcae
RqPu5xucEjTPT1atq5HcakNSl3O1pbLKR2Ga+lbsGSRbmGYicRuDbvWM1YEjTR57w4lNIW/kS8EF
FpNF+mqLGCGiTz+5WHwCncLWCBGXIOZqimca+mdEZ9fJ70FjhGpMhYOyYQviGvrkkV396UZkAD7T
RfDueD+T7Jn4GatE8MAAQ9ECmkqG2rT9swQbzsE1KS9wzUYhTuEdvTqEsqfcfFCV2ovXQ2A9MjyN
HXRTct4tcBp53M/sAG0Sd12LzO7cK9APgv50mUYXmx3PohJO3pnP9mLS9L/7fMqc/p8uqmFqQD2t
CgR/x0/ceGxmB5I/68rhBce3fJL7PpWPWpqyXAHgyB+7UrzGHRXzMgUNas0De6n+o8QDykZS4G4t
mHm3UZth++KIrs/iboSujb3WRx/qzL93V4Zd0gODgsf7VyqZrPCuP/fnXq5UboHqBtx/cDHvj0m0
xqQ7Ua7T76fQ9pe+GILTFLZkCOwLZFY03bq0Vakrj1PeUIN4OiBgbpzRG8Ru4A37v0uhlg5Q7Ggl
0hgsqSyAAyDlCamz/VBcLAJSvTsdvvZ5UioK/XNiCCR8ZBgjtaSDXVaLghyUvlIm65WOEBMW7sWR
1dE0vhJsWxakEQTt6ZWUz2x5nr7a5y2U5AShkS4NJpAwD7Szq6x20GrDs2WvUxswie8fsXi7FJl2
6bd+qwam4f1/c4FE9cCwQhlxmLA5/QUTmN45IsbyoxEtlOO2EMnCOKnVaGa+Ar0nx55pVL2a7yoE
VocEkTmVtXTUKOvYPzQrMFS1vnY9+8KwGtKTda0YwBXBLHgwqa+eM9txuvpeWqUoCGzFi88zoZ2t
sK3n7KQxN352JlyaZeLuQfixrwSwQmOBVmf/D9Qz1FaBY6KeiPi9tRHfH4ZsRjvChd63jLrPNjH2
wRLGVX8O+bhkMc9ZVkAfUU1E05QIaHcVwNxrasuhkC/b/Ie2RImjjXFlULm1hVu7UA5AM/cTeuFd
3Ko1HJpU8WXzzdqe1mByjnyMEx+XZVhNwRW/YXj61QL6beKME/6WLSMH7TXaoQ++wg5a8VmWEgyG
+Z/gCHU+V70Zq68ywPuz2ZGzsIcBund4J5ZigWvAJDsQiEMriddFvBS0YJP2eICXwvZ/aG1VQ5LG
0NxBATBMNnH/6HUvPqxP0wPQ90bzYBWPACgard8+eXv/B4wiVeCooQUDCLVFf4Y7cZAEy3+sNbbS
muJEuTwAXyUp2rlcosbfjNHraLJu3IumLWhSeCc0tG14LIPRFSoPYTI4/Lok0MnFnOjQSYFvuuqw
/m6QsEf7JZCkupNuxoihGyY1Q09x6fypKhU6L7CVxYhdapn5Kq9P1rddbv0IbhW2QM9SoKFSf/Hk
Q+zhM4kGtP/X45vCbH2drhI09Dpz4L1qGZt1H3qovkiEjuciYb3eNQKizicg6HVsfDIH+jD4o3UJ
smOfovtroWqIoVAMOcrTf/5rlZ4xFOzybuG3evtgwFgDiG3an1q/Xcp1OU51AF1A8t7CL155z4fF
huZzvrf1bmHcKo6FhmfE1jf2/xzPgXrZ9yHmtmFLchF3atzvWCFBFEl0/1tRoZ4fz4ZDyazSnZQB
KSwA1dmh2BUzFhemqF/8DoD2NqVvJOEms7+/ejXVGViclH93cOwPVG6SFEOPRKKocCLZldIeiNGb
o3TIpzYkpfFI30gkNgyhCWjh3Sm5nNypRukAeVcHQUmKmxnlAyT8/KDW8Ih2dtzKfLHWI/SqjO4j
hK+Ntwp9pg00ppeks+nwyhjMxhwjBXoj+hEP2NGno0qmUXL6bJGpO6QB26A3eVzNsDDbr9Sbdu9M
85h7Lchlh8cI+i06zabiw5DpLrUhSdF/spPWWis8TeIEtukCIFblHnLYimRaMA60ylXGWe6uyf68
SdeFUjO0eg2g2FxYKutLwVONvAMQ6J2gC620hTCoAh4yOpLYNxMMK05ivj4D22aao81XUwnHImMe
3l5CJv7UXoM+ac0wjmbWd/yy7tv/okKG7uR97CXdqE0DGanP4a3MDNS57cGBYzrEHn5Rf0DJcuE1
0aL7baJKJaTg7WbIiiSrcRMvdmi/bnYH4dWEutjn8bs4EGbpzd8DBgBwjS7uUf2O3Uw+PWXgz7bD
gbcrnSSDCsEn3TWYIhedTT8sX4pnGWb7VLNs828wMTOi9ZGwqpE64suaOdHMMHUyeTXG8Wldn2Js
zZ1k/DrXV4MtouA46OXYexX90qGWGlmKeNBs7Ekt3pffD0DOttFPS7rPiWf/caCYRchgl+F6CAPX
+GG79KyCOr6fMjIuIgkC03npJLIQZLfNHSjfBn0gdIFDpxnsiyRyc82ox4OhxTWBp/3TObFQR36D
cdJVaZA6/aShbL/+v7c3HD5EWYFokHT5q6GPT+24BgcqI3vxqBznieh3AtcAyBywk3jD9CK+RURk
mae2LT0h/RaqltqZrzt6oeA8FQjdLDaf4hbYLcgKwtyVoj76nAKN15mugV0zVgfKR5uf+xV4dJf3
pf75RuTd/Cb875RBKpAj5Hc+hDrj2pOgGkH133ZJ9KDHwn8l38q3JvTbWayVT7ViNuHlJMAVndkt
gu8OuqqIRZjleZgIt+lidB4aiD2bBDSu2UAt8ShZa+VEqkoecHDx0+wrFVgiGFaWt9ZDRBMGtdYQ
tx7B4OW8CvD3eXMjpxTIN2MZVsKiS2VHJhuqQHaEsCKHD39hBUkbCxidgKKNowe6OatIMXO5FzOi
d1lGfU0KqDlTBN0utmDVycJ/POtYRaQWpl861Ah/higRkbSsiIGiTSLDJ1nx4JIXA13bxN4lGWIi
mW0OsnwvtJiL3dfN4P9JDaYry/89KqMJ0b+MclI93bYzX9laKfVNazHlrIa50DEx/h0dsfeCp5FS
ONlekmXykFfao1P62YWhe/9rnd5rqwgj6+FVvrOQpDZfndt2EDr8SE13rGDjL7Q+JGBcNJwiWYGl
mcbyQqfQudYxfMuTs0OoesSuRlZXQh05aQmwc+qhl/mQchilh75UJP+hsgx9xE1KsvkKGe2i6eMC
NuemNm89/L76oGvuCuVMx1OTQf9rMdR8/3FQnUJLNBzty1fq6ANN4roSj9mKJihC9vY3SqAml0vf
t+krRbPiW4Dk286bXhQve03M2lsGSrIiX/5pnAclVGB5rcXYdql2k0Y1qsuy83lEgOy7YK7y99qO
UAHy2l0RELdSc0NLVvsc7PfZUxYZTiV+YMb6dZcFgKoUapGYa0YtEEZB6+KExGxd7k0Ey11lXTAp
IszANQUMm+JGxFskrWbJTct8V4FESBp7CW73JDaHqdb9uoUbuMmIXqHnPIrGptevtgjpq2gFALlD
mWeEQIYYm3dg+8S4Us/BTuoNqB6AZ3r/fgrP6SdfKrXB0/YC0LXlhUrjo6a+C18FarjXaTbzQK5F
gFjzdcn0S9IoRS+bE8Up9CT9daSp3u/kc3UWZ0kJR7dyGR+oqoL7TQDe86N9F8EwlGNHpm1wq2DZ
XvQQtA2Q4vJMRqwNiKKTIpFlbKxDelYamhCB0J232vtfdcPA/Id+R8Swd0gn/EnDwAClfSgS4Pxn
iOQJ1YYeLNwBljU/aW4e4liUzcfIUlWphdTUEmv+jaUaH0nf49QHQ00HJUTKYj6lk5Kgm5I/2D3G
i+ID/HA6I1ASqRoKoklj3j1bdeRjz2DuHWv07MbE7GiQ5UMfh7I/NtPa/Da4UJ8cIA1T5S1ra8HB
oMpVm7Gegf/RJb0ROo5PvqxKIrqtiFiFgOAaqwe+BHt88cMwXhSJ3jxJ+FFy6idNiOIISNACeNWC
/1o3UxipaS/M9T9TL0nqqXDD17OJ4wtuBrOXyFOESfWeKm94zT1H6LuE3aLF76Je56NCB5724alg
D6mYs/caChHKSITXeFLXe6NfvQJRDOaM+VLgRrp878LEZsFX6SaWWKl5Qozow90r7VAhRTCBhgVJ
AvuZosERKWZN9OY72UCQIPpk3oGMdsp6npYweISrqcUoU+GvWQp4f5T0NPKmT6j1B5TMBmD6LLrw
hpXWTZMgL+3JwHV6nTWOdNc64X/JBGjsxP+D5jaNCROvvjc5uss3teTlYH/GM3jcWxtDYT49CAyO
to9wxDjg5V1iOntyNO5ri81KEwnX/y7eSG4ZzkwnndPoF/8KbKxIaE2PSANsXsTX6zK/CxiIyorA
pK6GqO2iLkll0utR8m0ugslSfDRpwOkr/4N7j28vIUGeoR3SIKpvIYWpsLsdMmyJttwDlj/l5Z1d
jccjSBFSmG96uEo+o79sOjJ3/AGsnAsrRHDMS8zN6WRqIAGMY2YbdEYAaVMaaARG7CjvcH2qb7Ce
G2tqwlDJoF/Q8/+WIeRmmT9kknnJjl/lXoRlZMC/0O3Tl0V7c/YvNgb2sV1KYdZdVQyCPUxLc+KN
tZFdADkNlJOzZBLwYPPrj7WCKFvIsRhSB6yNXZMGe1NW4E41UXMkY8LvGTl4pYVJzRz0bfIk5VOz
nFesEM//qsm41E6N93uVnaY2rRPq77bGx3UC+138BQcZBTsRalNnhpM7cNCgvDiwaUji946sClC5
RBgCS4tAUUzxYFCBkpWVnIzBBiQS6BiXEvC6lmsR5sdlVdKUepXhkJZfDPUc5+WHApeO4rnJFK2j
tpWJVfoIlCzbGy2caEyhNfu38xExA0eu/3uQv7YYYHmXroDT+nG0EnETwar+yai+5wnPJ7qvbEXI
4T38J33Ct7YZl7p4M23JSbLCGR4yk/hJcNhk+PL8vBS0RmGDsLAHdTB8ORso8TVvc/ATWMw3faoE
b8B7TbwrS0Hrmp26T1wiH4JwFnuxS1+ztLfLisVEE1ZLC2yJGq3u+wDO4lFKSN7h0gtEjhzYPjEe
e+ob3jqFfSzL1yYHFRlFb5wrEY5gY/M7AussQVlvJzayRiSUiaJ8lAFY+dVo/oMQYXmjzkmhfYq1
EzogADQiDD5sQS8/OviPMO8JqmED1YjK0RJLb259YRg6vSHtwKBKEfoeWnqm7zBiOtS5rmb5/21W
HhaNS7VNBkqgkgDrYIgpCm6y88ffK5mgjKZM7mIIQOYPHgb749+YKinEvM9UwTLC5EdBsPLz7nE7
9e0jUtZzMyFrvaWjzLs0cZiUzY+DQIVqdEXDoF7kr3JHyvOO8IO/u5GWtldKAhjmx0TIxwGXz9No
CYKuTYvHU+4Q58Qn0wyPgRcjl4sfjMoyQiWW4lVJX1hmpteWPcvBRbB6k1en+DTfEk0TORJc+YTp
puJ2JP6TqVUfiykPMU18mf2NnC4WFRKt9j4m0DTYTei+bS1RvwkcDZv8Uz2Ah1gi/W+9txDlwENm
F5V2bDWUGZfrl+5N1gC8CnrUuATRTcmAk43bg10fgKD2O2UaWcgfv6cQeycuqnOw1UxvWALBUt71
fRobTYBwQV9Ziiqd/CPiDTGL5SYt3ev1I4BxaVkfpr7XZO2CLUt00bKtA0vCHft8B50/VSlFGKdY
mMrBHf8SzdZprBaV4xP7FUWyFTeSVNUR5IFOUgBQypFrFjseeS3ZLyfmu8wAafHDbgRDL9+/uTTR
hzQG9LtLGjSZOm0EkjGSpeax1l5FxSuHtJZm3N7vGaIfXDNqBHN0YELl6wuYvlk/0aqDtjIEN9As
tLpx7+o4Yu5ZIWmcz3IKeHNSaaPjNtobQuCkFN67NHI76aEHhcX2SgTAFg0N7eDgE1B55amIcGkr
lXyfS32eDIcn7m9lPp+ytpFlF53pq221F9fGwAXtD2DUyN9RYeoBFvMbRHi7+xDG6SDsqOVJF6JI
1yhrr/J1iiwWOqf0AHtgLRZqo5jcTKX00xIj9hUQdTbWQTDue2yf23dJwv7uciGgrOOxRY6Jxj33
u4J9rVIWGwZtEveNTwWrvEHUG0/z9t5Fv1k947W36sSkBfubdAuVVZ+IDgrBQv8b2L16lO0HY0iT
nMGC7YfHrZNwXe7sIcl6hOe/xECQJkhqguxWw7RF6cAFOdwYbAJj4DkMi7GDFzP420/sByJNqvSn
Ko0iFdpQvYEkRUpqpG6pgSIAfORLQJiXM58D6gpIRa7/iGZfeZqjP1kA+2ACjIF+B9amo3nRWtSM
kXvBtIz1Z7pVmEcsDEo/Lg00jlMrEOfhM79qqd/3lQiRoT30bo4VMWhuK5JQ1lGNhpmOe1YRIXod
oZpTQG81PTN4EGZWS9mrXN3HswOuO/4J+eu2gbH2miGjCMiEbBeNKeztni06yneF9MHetw5QsdlF
WtXT5S0SwIn8vf3gELbB2oRdscbwXqLj3cV+FLjS2PbGwP4PVSZUpo/NUBDmbORfcJT3XDN+4y+Y
Oejf99Oew2dV796vxYxE2cTPORG0wsuc/57FTrnmoebilWetDfBsV+hPjyZGOCim51qojjIL+0Ud
Ho+tOQ9WIxWA8tDVBYuBEOdGeFHgWxrwjDI9WcDiB7pGzMqpZWGYoJ7lhvYjVjpt8wo8NRpQJFpO
2ipFiHw00YW9S4VK5AzbmDyUrzL35nuyv39zZ8WFZF/6/2xHlBfzyuRLhsdT4kJmY0Ye00LPvWJi
FEv0rmhKlCp3CcU35VjAjtx8bkAJoXdn93fRtHf35HumIbMEQZkKv9mTdZrXIaICVzRLRFyv65Ih
9K1amItHXZChK6W7NngkVDKG/mEMNe8ajmnX/xYJrQQhwHdwcla9vORAdf3XDSoNkFPQpbbiga5S
kMKYkz8ZIO50i18a74mZTvkQWLYcv4Myh1IKkj0IHh48k0wiclcblgfvFwEB1NTfvV/N5JdLC2Se
Dam//m5SsrOpnzDwHTZ0UryRwyzjU0B95xaetK8wYj1rg7KDEj4XTxK9MKTs6Y3joTxsGNrsg9W6
ww0QgEeqBbUiPMD4VttXUoq8GEdijKYuh/rrCld8fiwF55HtQSdjcC5/1yhsVp5QCYk3FR5MmKvs
W4mmjyJAdf0UXqthIxO6Tc2GYlztEIuGECNxgBL17n1n1XASey+Kw3OGBuTtr+kV/NIF6bnWp2Cm
GhcCs2ffmkdb7tM+ACpqZHFi+fJCKtz3lKc5ZQ76IQuVOsLWcMXt5+gXwv+F11ot1piGsFnM2ph3
n+brcdsX8RWzSQzrHJbeVYanBBuaNUSFFnY78S9nYBQ4fnfErzGp8weUTBbRdVBn6ThGsAj7oVL9
s5mmVzQc72eOQIR1pcGWkKIFHAjULzPcQNKhC2dk5psVizhUj7tQAgH2Cn1Ix0eXvsDCfswBQY1m
CCyquQJv6ZEHdDK2Kcqz1NRUrMANSEfDyPH+o+BK5ib7L0kyKZ2rR0iHyNkF+l8TDv6sgMk77ZqU
x075MYZ53i/TFN75VJztuZwJWd/S/Wxo9IIxF0kLuz9w9HWVJxjF8f2o8WE6UqU7tuVYnxOVMxcA
ATwEsAMXclEpl+Qu1xXVmSH3KCcf9By1oMu3f/JvrU1LYB4sCY9BYo7YWw7GzhIn06ALq2rfrxSf
vnCsXr91s+34sREkzlDsv4v+/Ucu7cSTnUj6COvL+DIrYHynyV4EKEZLLaGga5JVPPQl5HDz8r7b
F4SCyzId+hWWr3e5IpBbfUNxgpeFW/IOZiyV2nDtg2l3zR4iPGzGb35UwvNOD/tSfM9IP9pYlmjh
AvtADWjl3Xp+/EuifZtLIQjwskHelt8J4yo2bTUYPlDFInXJIDe68lF+nIYUBqADNGnQ+ufnrFXr
2W7rTwEINNifo19QBpd0dtqQ5ZyUJufDWQTQ2hecnQyxR0JybhTFPgNRJGFXP6cTLSVT0g1S1bL3
1WWh60zZv2X7jDbGSYS6CSfL+Nx+q7cNi60wIHB1zi5X061z7rGB0P4DjcNw0dMyJY9CxnWReSff
qfcplErueFi/CD1q9LpOn5GGA7tc32+9pSv8Z75n080gqwDkAhz8uwxmapVplVMJG988dark18RP
gweOvFASaf4ujTKzZv6Q6hFRq704aNUcNN7NOi5+ccmuLr1rjLqJFc3ugk521m4dfRFU4jIQXcc3
TRv/X9lxCkJV3fASwUIZRAimhjXXjB8ZFzoyqaOJgcybDMR+SucZI2k7ywW5kdTFZ4WtUytG0ubU
cRxG2qbQDrwYHyPi0mfJQ9C2bFH9QKRfYxIh1GHRcLofJ4OBeAQzRQ6mvuyq/EIdU3eItl5BxSYl
Q+vgpMhouwky0G8+3OZVbOKUXbXoG57yZDv2gT2Ts+kruNO5eW5L5EOxPwvr96qKAvxa9R0PDM52
0O4aZrDjgEG8FRZ5TP0tIWk5IA7OMNQJAhHIU/uxqAf47Y0XpQGVTsg3QhBq4XEPZm0foVq3Sz1i
DfT/zS/UCnno/QY/dWVRDE2jP1QPEJ8Jk6Id240HfyzAfSBV7+7K0d4Jyq6PL3lthHvrMMjKbzi3
jO9xAVa5y+A8fEq0FN2N1niUOIv5o2UGv4GBJvokv2cIpubv1ZIVsqsYZJ9qFvMLHSVwwq+4xavq
MqW3AuKJnI3bOGycm9F/vNqqoUr0JIlaQgsT3SZzUdWbus7QCuMu9N4pgPt6RtgN1yFO06+h3CKH
qCp7pUAL8urNkZDu6jGGrTEHIeYTgP8CTPB1uMqtjitcYTzjuJ3a2cGgJHb2tLJp6zhGBO1xdp31
OnldOgdwvbxB+XeLfhKiVz0HGIB5nWEX+AYwj4FZ+3XgbZ7D67v5uaw8d9Zotlp54KOa5/ssCpg7
rkaDLXZIde0IKZI0X22y4/WYyUKOWhl5crUa2mzovpIrm5TMPwFv4pITvqgLUMk6NCE00UZvN4nx
3ew8DHgRIU2EU9agXvjuWxOgxhlOIiM/dHlXP/b0Eb2KD0NB7UJ9xhX+DJP2EQdvv7k0YHoJXQYL
fhHE9BKP0E9Su1fI845QVTiTHp8RR4wP2umfgAmr8oF2MUXXyD6QjpOUHd2PSO5hdcr5On6c9xCK
j7xD9WulIEciqezI3bfrdNromKRyOwBSKMEqWOTn6QsIcZKQymL3kP2ar5P7+ppgDaoA30nByF4D
ZhaK2MvtSaQdNADzMvJEhSzUCtE9dlyZ+EUWeznB/nJn+pXjPt5hVC42Hsb+NDNE0Uw5oOGcZZ0E
S3f3Wc7bZEkey/U9v7ErXTjt5X8e0md8pChQfp78lkOrGcr4pZg3c1AQ66CqxwSy7UTKyNyB69lp
HxoeEZyBGrprQl1qmujpb2OnKLW40P2CICR1f00plvPbkYilx67ji6EN17cozZydB3tlBtGChBpg
VsCLIEFk1+CRvnMTLUtYeISyVAhrME/VGPGf7/OMQ/NmSoArpwTJ59gShT3amHZr/EqgNHBUbl6v
I+IqSUTnG02AtO2BtSumvxMQAGL7xtjSK126TDPlk7YqBvRBSgVFwajYMWJE9CLGUVQuNEMZ3S/D
L15VH9Lewrtooi1rVDgwndhyq2lh+FGXxwmcYFCWcUUEJ/yQy+t6A7vaC89IpR8ncuu/qPKM5m+G
IiQSMrXcuxx0gXkKKx2dYHzcDkCPjZzrXbndPNtKM6Y1/t+rRi4nE700bSK1BY7p+wSFwFvCNeXn
klQDzChY4ksStxrtXw52ClFtgTlR/VgjuBwaD08Zy1nCNfjYFMh/MxezZGgfIpSFtQ2XonaHDLaZ
HhNdeWhTJBVaJ3CpV/tp0t0HDqjF86LZYimheuNt3bo0afCmdsrjM8G0DfKSsNwQef0Xx64xMukR
49Ad2HoGGtBkujtQVApS+4CeQUTbrGyraE2OTq99WW5PBrNuf902vKmLBRzPfgvOJ27x7N3IsKc6
1+/uVeyrrUMZ0DBBLFR3Os8x7amNUw3iuA1q5csjUfZsHapOpB3uy/NH0L9TD2A0xMHCyZEIGd7d
mzrPAnb/4SD8oXgAJFpyPRrOEsNMKiXKZgVJ0H4VOKVfDd81peEM6V1q7bz1sitFq7MLfFJkiYMU
NdPkbMtWo76lAKKrjIM+H1+hBcjFfCydKKaddOfB7yo7dxYbniDqHR/evNXnXj0t0Dw1FnZwXnyq
Nd81GyzZo03Q8XDde0fdN02TO3n6qYNVuiirH/5e3Ha0ticATX2s+PnIlOq0haZDCKuQ9Bsc1OUx
IDE9uFR40oWJbyvqSmGkjhA+49bRPpYw/Ct4iqodwhwR133gomsN4awKjGWQM7YKmrDn/qUo8pJe
+9fYJl4QVaDcyIM8SbxWR38LKcCBwK1ZkrT+1xqJ9+K1jB5xVdYkXqnBa8nquPbCC5N1qq/wiJaJ
IaQeg4h2x0m28d7DHF0t4w4H9sJWmG+XsZyoQAYaXyLN/Q2/iiWNkd36pStW5JeoZ1dDvqRsauYb
t3kJlsMccnODAlk+qEomDN1BmDQTIlv5fRDWs2fUEXMQdMpEfq7JUYftwAtNmtFON8uyWp8OghGk
kc9s9EIlIiCI1cFoRdc+pxGXiRaoLRU8TSY3iuJaHvfI4pxrd+jUmMUzqfY/4+Hd6nPKqw0rxOxI
i1TzaMtGa4uu88WePSZWxFF7CcSPW0tW5n2ptPDOo8KlLMtkPrtzypKloiTantF3qYPmDUqWuGOE
scwBr/MrjYCd28lbEtGgU9yYt5zHjlOSRQjWPXBKpi7zmy+q4T1utAxO0bVMqTKkcDtDmdmo5sS1
h7cj8BFIactZRZDZN3JrWdGeb38QBbJeD15oh0q3LTEhKElnQxtjuhC9Nagne1X6DKWZSQKoLmG5
0j7M8I0D5QXJXgbT84KKEQdtIBoRnfWT9PjRa4PwphofElzXdd0c0NpSR6nt2lPfUoScnf7CMhL1
51wf/w7o1tXpbHYHofbVAOpc6A1mYyKkCp6Gt9vVjj9B/jrImR+3hTPpqoXCjiLJB9CPzEwF/+Pd
7k2qZgdxWuQTc4l9yHEAZ//ha2yxpN6vwy7pirxADxTUd+1S2x8PEBzR6KwDLxpafv9PvO5j/mq0
QU/hXSgksNtEC2kVz4vLKo8ZLQa3xRpsrNSl+jqKrLxErsVyGhKYkEg9WK4dWVEaET0qlHFmMuR0
r0+sh3/RPZC+Cji+yCimKprb9UpcsNYH64fly4yAmnqxt58REzkrGKVNCMFylAEQUAmhDMlP61jK
ryYB5sRkmr3ciLJaV7uS7hgaQ5ovWdgHFhv00PNk9gwT9IbA294r3rYXgzjSpktju5ofi/6M8/G1
A0wGtjdHpYcAf01NGcywy+jo/aTjgyvMftqAaXrS+ZSuS2cCGr1tDv0UAVWaRj41ju9DfofFdArt
QzJvXi5DGWHUcM8HWQUyuDxq5GchDvGGmWtJPbJFSWT3Bt0szk5mQQ++W9bAb88vWrDtSeYbqaPb
NkX705neoqwZxVfltDYUyJsEfBsJBXY7tOkYbQtnHNznIu2EAumJ+Ftw9LIE8rWDuaSV76wiXDI0
K09gOyErIvu+ntr8T2vKLYe6puGTEyWf104kmYjCMAgH6IA5jtmylxQcov2nHpWsT1nGI8E/xSJL
Vy39RIIZpSXbU+FfPLlXiYqVjytLR9kCN21za4d3Z3uUUxTVY0qbEcVMalhZhBrYgSq1dz5J523L
0bzSk7IkUdPYZHDlUip+YVcKHZoi1MGd7yWydQDx0KlFh3h25J4nR+fFQkcNI57y/qx0T095m/tP
f62h6gxavF/uuuaskAsOS7zy8E4b0qVNOutOfcUYDKunqS1sG34Uoor5l3KN6sDPBaNyWaVZ+jN7
IweplV7UnfD8D7wF4tq7NeH7eIDFm9CiRcIUsG5v6AkqE1FM2OPYlIbxXWO/IxkfwS62Em1ijdAd
plwNWzEGn4wSzqYG4+J9D40fP5vHHiLfPuO423SjR5LFsjtUzXmekODioUjorVP65rKWNt1cnIES
6lkqNZf7fFVus7Eqauau62ThdW1HsfYY2QVvcvzDBsnCyiFTzJMSbyH4wRBcGhn36EFnkyFLs6Uc
F2a5v0H8HGtYbZIe+ifGqRQZXP/OZB1CyZ8nE40xqoCH7hZRC6B4dMzO0fQzP1QmTJC2V3eJQ7h4
H0nBDhwI1PJVLgGui9+XBoUizSeIEAU8NQc2gdjZFRKyqIbpTVbq4PVOYGDC9ZgWA29/uZacQ9/K
nN8vVpM54P0Cq+XlOZbPnXH08romgk8swsPoxDM/pzZKl+XJY6PZ7PqrpERds/qnTA4L6ZtMGgKm
75XwBBR5F33TvQdeL/c1hc0vRxnEaGK/KOqczHUpgVdXY9yCC5r3I4ZgTWjvjzqs8uf920aUrRFk
6EA5ufhRgomDXA3/larZ6De3JcLOrL7kZ/GH5gxWw2oE5oRXon2NiLFXQ/pnIWzIhGHnyo7/DXLG
VgrwVuXr4haIipY7HL84pzCHDcNUQfMzAkUOemLwQayusOI598MN4H//+WWHslS9jWcFbztrlIJy
h8tPJC+sv+JkpgxNimrTHVh5ypr2uBCh4kAsrEFLfU4kSBNTsRXj4Er3yG6/yGXh3elO4d7+p2Qf
Gbl0dVXG06tpq2XVJoJI6z/mc3Gq5DRkp8VDTm6+ynsEyBW16gErc6by5X+sHbyPVeKH8uEznkgS
s4+l3z2TpUTyXM289bxzcNE9uREw6aDhTTWkuvbSbBWUvtm93Ybuh+UIeIJMLQN5mq1QygLNdlC3
5EpfSxRJG5JGo2IQDk88CaU2TzN7a36Ltoo8f5ZmMC4eOwTGD0vSVBwvNjAqVnDdfsJWxrP+e3m+
57e1s+EM3pGq9iipi9ZoLoc5zVoFRSHcDkn+E8tPTfn/mu8w6saJ4XUGqNSS5Z/bZ54NWTwZY0kt
CfJM1B2JD/d+mR1SDl4opybLFBgTo1AF91mJatflwssfI1SBx98Ry3qFZoeSqoIRyEYSmJM4nL0h
V+1XegK+brror3CMxb5MhLWDtIWcnMfFUI294JWcd/pQf6Qcrpz7aDkHDRihmufZ0+JPRGjfzXFf
/rMcpwnvoo/fcNRmQAPGIRD9MWf2kKzKLZ9EuVJtWYXyNbIkktS8x48IKk21Kewn4Aim1JPmlpoU
s6nrMPbwbrPXAZkwKCQZ9cXV01Hhv+85NyxB4rz8QNDF3Yj5eIktTgjS9EsR1cqAMoEnKWKeK3pM
gernFI32tuSkblpL8HQ75lZEOtg8LZ5kaqJXesd730ooykdF1jsXlhWGeONzgPL53PEt5HQ+SauM
+Z43vQNstYkodormrztrjHbzXyclaDpe44QazKPvg87yAKqF7c3xo595jbgEhrMq2HZlEL7i6I1Z
hRkby91xE6YHQsBKMQK7Z2EJs7K4D4wsWWHWR7CglS5+yI6zF7niVwSaXvIdVh4RCsNKfHvy+WYZ
HtnYVNJqZde8j0ecd8S8cB4H9QQgsGSt3GBMAEZfLWL9CG8mdYLLf2WfrpyHMOXdzLK+sfQGrooH
EjL2O/QIB/ND6niadqBSgacKpg3M25KlPf7UQ5naHzOn8EfLWh4CLlu1R2MiMrotDc8GAZFdWgDT
8YKHZuCLZlGG2PiypDLT0VKMXHBqFX263dt95c9J9asohuIqu3K9JWW6XB6vFQ/vzDqQeuPKbP6e
a4EIPL8vO7+Zts6/Zp9l9R3SYEhH1bqlQvs8DfgUlZNmF0ieKpB5pp3wGCUwk5v6SOJ+x2mBr4Np
+JBXPVoyy7qFH86ckr4PZYyp9On2yZ+n2y4Jkd0/Q064ah7G5L02CII3R3V5qyklACkNzkeNgWNN
KJWLgYvIKm9ov8oe+JqBr5IyUL8F+njA+4nXmCMYYyPLQOgcXxc/Lj/1GwuksVwgCKbqhnM0lgpe
YbhLlzV/2wwfAHoDnvhv7sgQarpWp2bBduiaobPwxyJGZI2Gi8mbqYVT4Sr7pa2LgTxrzGBeFQ5b
wSzzpv1dcYSsi6GQTgws8NOtaMUbKyJrhHjhnA80Wf/c1QOMzKuTZkBAaQNpFmKeMQMxNdhHIpqY
Nm1R/398pbn2JOIBfwuSBgE4X8UCu7VTY8QPouFzGQH2fNAGUKlbuICJ9ekj4NEEhSQDN7vyYH/J
jmBmv25/FaSjw44Nukvd73uxB/iD7W6qCboj8RKACAzYn6yQzj0koIOOJ5bCvkaW4vYWa3lhDaC7
MJfP+m/EEdglyq8E7okm4e+sZHRQ78TFyhQFkoXTTvllgfCCYGFolcPgMfEByNeA19laX1Zi7I7Z
THMDd8YSDjclaeajwd7Suf08Dcv6fwvRE3NH9LPi3sjloqyVfGQ6OvG7RzbYUFSMuON4NN4AtdmF
4e/ho76cJ40juKxrM7ek+u5+Xt1Z4ERpz5PW4tk24ekCuN8kNCHlFd9j63h9bYuTPerpqfsVbLoH
nQCvdnq0ncSQMvJXC0v8rormSvkWvJn5vScmdmX7l99VmmKwGiAx6CclfV8517VU7ETiLsEYFq3e
IZKqWa9scBUA+h9aP8WmYtBRdfzd8e6snm+DtM/JMbL9es+INS/XSG7hrIS6p3XcQSjvvmvXAmx1
23OsSOMjl2hnw6dZy1rCqwA1p+zxNpBJJbGYkvYKErsKMkMF8bZ2jPvVtoHr6jupYT9wCMX0CsAM
QLTarB5v21zMIpktxtogKAgoxDmconiUT/Rbe2KXrP8k6T5HddcY7rjWJQkkC6PMkm6VU8RP4Fp5
vMfayOdfwR96IcbPBWEsRX0Xv87z+3OQn737f27L18cafxqgpozIYTk2NHcn/mAtXHmQhKTViY2e
mzNe/YdxlZi+b/060EtNWgjuyGfz8acPNKxD0p8+3o1wvi+0+05708suANRJBU7d63mnTLGf3ZbG
q3mzUVxTrRaQqUqWAxab2ORvaBeHHsmXTAU/bGF4o/kTh5og4rLakfu9uxOa9ThRlTcwSSpDdw/3
DY5/GelfGut5PdLMFPdOyJU3nQPr9vy2K3glTDiAtpEPoUDJ9Uy+T8GjYy/3VZZt2upnGqHXX755
UuLUz643wJxAOEJLRSym2viARLqD1pUJPc0IAtgd5Zt6q8+A1fkUnZSh/FCMGNK9qG3b1eNkjlDy
QwCaB4856/aSVn0Euz/dk5cfhzk2YLFK71WspCbx5aONGUiSzmpNzFhA2oS1FuebSTUkqsnmcq/a
HM2aJUFHuStnd1+IfTrH9Acjbz0lUBOVXAGgf1H40n1LPNzyDOYgxW5K4i3EHJddtn1fOocj5QvT
xmTe5wAQzG2+9sKTquSmO+cc0UfjysT8oTcXnAdep3waKT+W3VSzZgEcaz0Swc6yuywqYDxP4X+l
zGfTipitqPKjB9ivyUW9P+cGWUXOtCj1YuG2zMtrqxYr7d+52oF9FMSY+pQvKvoYfuWGAW5AThC8
mp65GhvqxSv4NIrEKxEhju7txCq56/83gIIgfcsS45Ti5XOFU+Jb7MbpaR2l6Ry7F1yth9Av4g5v
3PDLyrDsTrK76HVNbv1tJCX9VZrQxnZzr4YnWtvKv41XJYy9I8zGu7He3phgn5UhwijYiRqg35fZ
KKWl1qnIbgJlfDw3vynIH5eZr6ULKr67vrvYI9L+6WxYLEZDM4vNf0qBqgPd11hf+17VNwqt5jk4
xrTNAGWGCGD31/8dJENdELIsNv3IodhHlUDqVNXldY0Pipx2gNU9mgWmw9NN0UsC5RbYMmHRVawZ
OvzOyr7TR/oqn4ENVGOyzg+zjDVYdmI2tdc9zKGRUPzPWo0rm4ZVdyJH3h4XJ4l/NSZXwlTa3QYl
7n3bpmspwW4CdhmuHwLuxpWPTFxjqw3ELnck+PlFxSVK6pTh8PFK2k98ILQs2xHoAY9iBgvwNksu
t7YUUOdOFMzltBq3eHlES1gf0kSYIVct+liyeSTKAKbt510WYgw3x8Q3zfxn+rLNiOaYYL91tkfl
i09h/5b570Y6eYVhGZMyRbulhLS5xL6FshaicPqaIoiQcilQ7dOP5KdY9NGAdiCYIaemCWy4Vb4B
goomhDYS3w4NI2/H4tRqhg9AfHk/3wradPGFnrEn04hlxHDegb7TDmIPhsVBcGH0wBuGkQNJACJ4
VomFRBuRamqiAyudku+5OD58J57CJCV3j/9vQD73H15VOL1SXopRt1i6VVzQWYSBhrclkdDqC6oR
d1pGaj6lQbMe9A10t+sMXAYBlafnGKJhWCWeeceGA7bYTTgjnMUcdl77U1lJ3g2p3HUXUgIkqk/4
58XoiYD8RzAbrD+L7IcjH5i6hV4/Deb1YvK4xxwK8nBUuQoCcxW9cQx5DlhFXaxSTWkmbmbbPN6a
3V9IhADF2cZQqbN+H0yeR9RJ3HpfLSCRgVy/7pL4GkQ65lkVKnpNiQnlcAMEoiivTPFT0yygw2SL
CMgIs+i9RnZy6axroSa8qlPzaaFgqzL1C6AXGQJ7iGGrE8R+kvklHhQFNULKTALO4y09K8d9Ls/R
hx1+1OgfsbO9pujsAoVHEZOp6wetQOVfumy/akdlYT13dH8TGgNEaAkSA06A01fhkBSzY2lHyt9y
QOBI3Qlp2VavJ0EuZ7O95eoIK3v5Qwmnyz2oNq3j2VLzlp+WomQY2I7gYNBqEk0k0bCmBz6S/hMZ
Ar1LQNY10NzUzWeQmqHYzyvV0lck+ujFv64JYOD4lfWpOY1/HAt4+kyZFnllXUCXAbkwIEB9TJmy
KgvF7+tRs/YT0NBRft5X61oXXSC//AM5HiCoMAGTc+svVv4y94tVXIdqg1yw+B3yekrakummk+Kb
vhlBKq+upMKu/P5PxwUjiE5RaAqCMLFjxWs83AvWfnwVEnSkI/e0krv6QWOcZech0//1Laqi0GPm
du2BpEkEn6bw7gTWwT/lokjjCf+ODVgbGhRjkd6n4xEJ8Myrj/yyK4EVWJLW1RbD47viJaLVr0hw
jk4EEqqfMOElF1k1TJe8Nl66kq+W1HOdWNwbLA/9m0tY5MWLc9J6ncLKv+Nc/qpOeH/9z5Jl3vOr
CtMQq7VyH6+fcGgytylZaSVCmXYwCuZKqffBGf/AX1xq/dTWQXU7FRJ7blCj/cBE8t8DDEGyZJJl
QOZkiF9giLFypM3+Ao6k3Wb+gMjpqlobW0bLtiapg5cNAQWgjhu8NE7xvx/Hp0NMEwCM88W9UpIr
w/bB81B9Sm5nsEpH7wBwrclwXL3DBIJzJkCvP29XN+bzNZEjHg1OnWGgYHIgkgxv48BYY/ACUPbb
DE8FYgJIZRUrlkFmkQ9xLHAylFpNYePKqKIoR2Sk4ImDJUFW0UNCW6bO1emNYXzkX2PGHpsmmpQU
f4Nb76pJCzF7eM1AmYavLw5m093OIGOXNX5GfZzjSBSJPom81g5DV1Wl8PRLjaRuqVXEOi45fRSJ
Pd5xL7IbRIwd8/EZYGwosPbVHQRkCZaCc9+CqvapVp9rm/5ZjELyDqoW4qnEthsqVjsZG5SmkMQ4
8RASjUHu/cOeil4M+u9KgA/5OSy0sU9DJ7OThVNEanq5hhr5wm3CSaOsvJPIbIsKUfaBCrMPDioO
5WJSczfsu69m9ClQ9hAu0ZcXCI1C10vfV+wUzOAdxggEZZY8ZrAtIgowH8jyVIyYXhbzNEjuy404
B4RS3qUKdLxz+niotFdt+9i3ImwMGFO9qwctUiUMZwMQr3IU9mVlUz7Q7wRpuX5uXY02YMaM79Qv
MjGQ0am/N7BkHe8itpiHV89H7RFeDgA1k0c/TL3bdlsWSf0nByyNGZk2PqctGZiltQ8btAXxTHE/
Sy2nDvTY4YT1LaDmNYoOz+uUmeWQvNOpTFn5U/k4pCAD+JPWhOflhHqrIhiMc/MH+DY3lmfqwnPx
H3vfvA5+CbSVygSePey2j31umxhhAV3CIFPQqcckOSBaXkkb/GySaJEQX+o4LMI7HQVsIca2vim3
bxPVdmK/lGtslTfeYk9NTX5Lxgi+qxd9QDx6/YrKV9+NNt//X2x8pj9GH9Y3awQ+eFPL9SMvebu/
K1bV2vu2xM+eBJNJ+tOsxykf+RLH2D/u+xqEXKEgQ/Yb5TiHB1ZDyJnd6VaQX1a5vvD450Hh0wl3
yiMY/7hKFQhvdcXljZFihv25teXQVsL1hEJI5+yNnsoAB7vy9KM6R1BuCBUSAzD2mDYp+hNewqUN
zGWzb0RZyIFlN4LrSVzlgi9b52je5/y9zoGYg5d+vmjwYdxIi0r7ZWXXt0pacHBCfi4kdswUIFbf
Ay+xRtRT1CI1oVXdKTd4HS5znhtdG7TL8ajqPcGPZIgQ2pUwEVK0DrSwMC01ynBzrP1NtamtTb61
SmnM94ksVmzwGPe8Zr3uvov9g8d+rhUiw1LY2TCfH4bP3pKvYbN7XBBGvP4mM46iRHG+RAZY7rUY
ElSQ30Puqb7hHyzZEGCGarYBI5rp3dczW+uuQQ2UYUmZaDQ73O/eE2mK5BN4FhxTXJIHzcgioqRd
Qb8xm8Q7QrDVI8ohfqGHMdm4ogzF/UIwVBYXMdFTPhpH+e5u0COllNtTgpBzrMitgc08mR0hBiEz
bQTfioVsrYG76XeNSMbVYtr5+R4O0/KUWgOswLT9vwDgKehFgWffvbyCfv3Z3a5XS2HOd/fPiDsk
V61yJaxMBC8TJtx7AWyn9Y2MiLU3JKLu4XlT55M6NIgSzEdcuERGgnZ+/LXmm1fsA86axpHKAmOf
/YVAkluij9T3kPuENW384FNnjptc/wrxKuQQ5adYpeNoqjtAEF+VnRfw3pxA27KShCxTULGHth6o
jf/+yK2KmjdxedjPEELsXZl0JawyQLspnBvMs4939Ea6jHA/KUXt6hihVIcKRyauJPsvQi8Jy5Jv
fmfJ3bMekyEWSHZ5hkmy7gzVcbjsFdK71+hok2Pe6SPZsqs8i12nbNDuNNcBkNzfy/CLD2N91OHC
fRtYB2I7iZVvxva8RcfmP+EAo4u65nn5BdU/oG3b103SVJYPBwrKH9RoX2mBktdxpBGgQxW85LDb
pLOwTnpWNh4IW1M8SIHYEWfSLoDf5uHg3ELaNkGnR+rTLw0VPtdXd4FNpaqs6FIP3mG0eluOruRc
uBcvGv/HzoRYqGrs8zTBPH9DDQTF6owXiAZezXI3Mia/N1IthMh1p9cpJOduvJv5GgjXOpoOdMsS
dIpfZZHjl/1FhYJjzjvWPeL6Fk3OKRZ092674xF+j011pUTj5KCwxVAikHrfE0GzSr2clT5fq4IF
pfh56ZJNhfBvAOfH3ZIzlT26d0Nklf+lx9jhnT4p+iO0R3ODsUiX1cSvSDX568ZyOtF4d+ACMoKa
bjEo+JwwrJYpprlfYA6ixGIIfmY4kwTO2DedraiBMWJ1Fq+DS2fjUOCAGohScV6eZUVvMjWwKn9p
zhkjEfxN68IOtTfEMxZ3z8MbGSpiZ+fYrpwUMabVubdEFr1FgGGgQAHgjawFqrNYGTxxPlav+ySj
cH31MnkYtLOqspGS+VYMrChj4Q8uSzuFVpwHIImYUYOBK+dSxAOk3DayaM8rT0J9AWg8jvOYdUVM
2g0WoqJ0iMSc3fJy4KULdF1ztx8lW4HkDZEeLHGYvJ3c+QXyPO99ZTnnqqT+7FRNsTKD8wU/FVOk
v3IHc0GbbzCV7QbdonShJr3UXjYNSCuoX5i9FVtUVaAe0ycunn9vSFjbBiClN4g7u/yjW21WykpM
7gOs3+eyNfd+Z45zQ//utvaAZbKMtUdqtFg5HpceCpCKFn3L8Q6KGnTDFvfuX2XElwy54vLzp6pe
Mmtedn5dPLXhEhyiu95xWH+TWpOuJ+idwwu5wMy4Wnw3gc8ZVH1TmP6jaDYHojozF6h6kMsSrWre
67rr/sLa94mwG/m4albjKydZ/2hsBl1K3pQgO3GTE2ODuShZx82QoGQhl0U7O25pWGUlmRCmeKRH
mOOMTmRdoFbg+cGW57gQhDyMRzEWPxACZwMUQpGU6XFnxTQfZSn73QA8pIFvut2QeOt1q0VfUerX
yT5KGmKjEL4f+VD8Hs5YHGoZUH5CwuniafQhIw3yrrvDeoa5yK8d2XrpPRdc+c3eyUNHOJvxXu0I
Kmd5Ms7Xn2KaUifZO0snUuMp6f5Mgtu71lCZj9sGfQeH2Ncn558BPFyWp+446uhmjZfTjKPi3PAy
KxbnxG1mVrFUQXWHY+thg6QWv6H6JAT5mX/a6fnU+pbzKr7JZbd7g5ZJjKjGUQ97Zs7osHyMIpwQ
veAf8QASoJeZbNn4owiJCHW2p+sw9VM1AWm1eSNx/rdfhjIUniiOP+ghv2vlmG/JuN0kZgLofCet
DK8RSIw7ZS68w3a9Y/r77p4+Hjvlvve4y5juDi7uuHuk9JvruH8E+Nhs7bSeaQ4Q7/o6ElpX0XjV
PtxdZiZJt20ATJUgfghUdcCY0T47BaNOuFl2piI28vdEM+BY7pDGoXI4vzcMTU49dxb3LaS5bskQ
rtEMVy9pEXhLFEcC+L909lgU9NJdAOUmT2gZ+whDGCaHiel0Qh9WLkDOPAg5pLWaqV7mq5zEhftm
ZoRk/Tw4en5Ci76phzavE90u9rB/qXhD4XYBudOIu1/lQSAzupTvMEO3Z92r+TQsOiG/hGT2pP+S
NmxBgWZ/ETaTboyhtnmuDNH3eo9QCrhjwMNtJ2mePwXZ9xVL9odK3M6X05m0iEYorrz18vu4Cpqm
FqNSx2KrC/Hm5QeavlH2mYg6DgXg1oYOu+/CeGuop656O8I8K561G3eR7HgvqAYP/CyPWjBf0U7D
e0wjaL/gEw/jwj6TN2kak/cDkJR0EhBf9Wgziu7vK7vdsREWs9Wig8U/Na/tBEJdMnWJb5bbtHe+
KJSQxuhd8+FD3COffBLc0zbFlZDgq1ZKDvpElWnXW8M/Kw1zsS5EWYu2C3w5MsMW2IPGCALwqfC+
dva5Ghylf8sjksZFe6MOm8R2OKIjA7ZwcnByNmV0hFLpxzBJX/e7sQVomT5AWFgdarve2c25sl/y
lPvIYMjmyrOGOhSdJvtl/pkpExRztY3CCO6bqDZAmt7ykdk32eFFK/RnbCz2jM/69PNKqjY1sYOW
8UfLE6MiQie5ntGZh4UiL7Bje/SweHZ7RcGjbABtZZHvhJql7rU4BEDraDQvE9tQKU61Tn4eo7K5
s2tcN6tgHCRZipOgJ5xtvf92AmOwtpdGDObvH1wnXuy30Ji2Z9pHxQ431KKlTxyG1EWLvT8dEXoY
35jsoYRYeWinn4RVPEMJC4c93LnNRqlxCFRI+7IUwG9Cv3bJNHmR7rSpSQikQswhLNMkytQBqm3t
+knd/bDTKmFD2MWfcURO3eLKmm7IxlLqSk+LZ8NIqmVC8aQ/XTxfQBZBdHI5StGzZEXj9Y0/kuhb
dpIybrCFbATf8jnJKovuIjXtnu4pkSrqo6Dy82UWW1ZU27CGWI04m43CePLA2ZaFnR7oBFax0M2l
NFqs4uw4sMac1O+pNxs2esAgrjVgHNu7n35vAp1H6DbHKFCOadZ50rm9N0h+zD0nYi/Wq8cYK57s
AdJMUBjAg24gzOlAo4e/IpsNfrsytALV2Ykzy4iJ5BejDPjIpsNqiAxVEc4CebM6C32f3dJsxDNI
z9uAPcck4KfPbdgFYUUJAw1RYwv3cQ9zSUs6b7e5aKirTiljSK6WlFh1zdqv9M5hPUg4jGQ5915y
QdokxxnqZgFcSm2E71cdVCdhnZv/Zu5jJYcP88a4WIEVT/9VPYMSTPF+CP1o0L4wagthZASFoaQz
jKLgvJBOXm2WQyCjF5a5JKaVHzHMfh52JLEIoBa3Ocufq+zV0rPPYewWW0kaErlzAh6RWqw1EIyv
lJssPJPPYPqdc9ACvpnd/8bDvOnY1luPxlW+MM6qvOEdYEezI/QTzvXFJW/41QKC0EpUo0QvkuMm
Q2RoGfZf2n3GCivPfzmF6QDikjuiB5NZep2lRSNSC1mq/3V7W5fw9hnByhW8aFqh4CgQ0QUVYZ45
YLO4JQawI7t1pHrRzyHyIrMLC2IRNaFTTvWyHb7Aw2yMUlw7hGa4+XOx5UXGH4UGNqvbDpjXm4EZ
61TET2MkBdE960+hGVIW3vaw8EGTIQAXG4awy4hwk76lykluUbKcAwKfhujE4lgXykcvESTgrvn7
hNrenMX9uKZxEN3wI2kCEcS/hq/zMEsl5L7KgELKLKCw66tQTn3zy6Ob108+Ns9H6wOURvTAzLpL
y2T2ZrxHyeJcn4JR2dB7dA1JBdtXVM/ILDiuYp1+tybq6Qh3lAawTJKZeqpfjITPrFLAuL0yksP+
UuDsa/Q4kr0uC27ZBYGvtWDtb63L3x/tq0Hy+TBiYv1WctO9PDmpdUIaLb2q9PTDEC849bu8FJJX
uGR3rSjrggZddeRmhHhgjxUmsUwF/8/qPjKgXVsCQncKGXFfKYf8/hIFY4emN7ZCeeLlzMRdW77T
5ufa+chJsS25fJagrz5L7Qy85sF7abLL0Ka76BBcJqkNZD1MwS4XyIflmeJ9K4Z5fSXc4yWo/0fh
Ia2uqJ701UO65VGe0zqulM2aPbzrfZ83aN+t61LaJw4IN18rrY5Y4UJiKTIYai0chQmWMcTd9qcT
z9zb/puhZAVExDkpHUoeEoBBbxZ5Snu0exXByPNiRbczdL7JrXQcgXapWlDwYAoLx9BQu3lTJFKP
u6L1xt/Ex+nNaNs6YgYRAWpACesGTncThqAfUd1TZbHWmU3bFyzrKWWLgOceqLh8dox7T3Q8bc53
RYO11r8kb2oeNGQN3bztV3mktpkPENhYboNICKYhwGElb45nhuvWaylxK2etxfKRo6uaKC3bC6+X
JJSQ8xPP1P+3HlH1uHyodpW46BA0UEKaVspNyYAskv8h0Jfa5BlMr4YKE1TNGSug+IA5ugz47Jn3
5jxYYjdkYIlui4+Qaij0Hv645UW2QLvAjEhLaZrffDDBPr1cqUGXXhDMurkaOO9KLpwf6Ooi9NWH
9LuhwuF4irxH9kgXk91iFdmWkAlwI8KEKwezoi93KfGhwgwCVddpbCuJS/1jCWdkAAEAcqBWbaLM
zvoXy+UgiAGUKaYLOGe1OhjlXaHAy6HGVjx8UVYre808kpysqagfW0xwiOW/Ul5K36PkzL/VhUXj
VTUmHta4B4rmf3QMnkqTV9PF4E9tg+2n8mKgxMI6WMrZwIv15RN5mivmaTmWNLSzjcGU4jea6xSV
uDMVGd/d5FDX10JiaadoSsNdQJYYuasql8t9UpcNdvbpRtssi1/hzQiSLzr/1NuvUt0NFWCUckiw
1/zlnE6wMa9nLc23hDgTn7Rcv+siFgR+w8YirJAlW9Pa93G/+OUEVbWrk0sb8OFMYTZtlb6iHKuC
VyQ+MBexbO/qSrrRqyi5RPZ1+6yD/fB46h584J93qaFTTPHF4LXCIdhgGiSow6/o3bHkwbXd/X2U
odoXDmr0I/JtYaKZrFQZoADLjEODHNq3jVK1TEtKW05JbYCesJtowxvPnHEICm7+Q+n66RbdTXuP
mPFU5GtJdqFIv/Uclq+vUP7D5QmOni8wanzkqPyGgSUsLgt4JEl9Y8gZI2+LSasFIAzCWwrTJEhg
8tbpTa/hKjT5q/hrmKJuntuIFUV+g8um8TeZlMv15Ll6rwd48qZWSFJuaCLR5+I7/kxaL5UOwuhw
HHPwc9/HAmvBnkI8o+8ntJjxxAu8nFn+rPLiuLMUnmeZQq6voNbDpn1vMdcWc6C3QCKiEyQnEIex
ckhbRguHtTkuAiPR8WfRNfOxksrPL4r91UgheLN9Mt52AG5F2yuYyw/wvTNGm5apBvBudTlV4dW1
jntr3coh/Jt6138LAvR7SSVN/bblt6TZqycR6pjmbguDaeaZuV5vAd/p1q92gvM95Jz+6KNN9kzz
iCnhqRTVZjm2T9K3hwa/H0P+2og+B77XrmYPVjTROitgNDwezRc5azwQb99kpbbIs1ltTvKwL/so
TPOAEjeoOaaf0s8Zq8YMyArZj7oEhtSPJG1fVOazW362lwZKxhuOoFQObXveBfZ7VOwitklbHg2y
z6V6wxVgYakcFbPSKLSnzx/Wd91O/2n7o+Rz34Q40ndnfEkAqGdQYO8LGfKa1gmHLiTAcMVz2ZxA
IVLtFIJ2IeFOt9hN2jWuiP4GLUmmjndB9hAzQx/GWCpouJrW5JSPuKEYuWrj1ZQb3n1Ep8XPy1+G
JHPTHg4H9CbT4J3leMiWySYKOlCQYHGnRYkt+VN5XlpaFIHcp4N7MWgqNM/WHBbIM1FVv7VXGrsL
1fJImqDNgzJwUH6MiZv3gUQH3QngChOvLWINrMxEAOstqxCrNcHFj7+teMSOg2B1bkwT31CzeUP1
BRX1qPByMNRLvxKGTl4//zeoXtGp6rseU6jnIuAWShyViHd+d0BEbnYoHuKc0nN1WxAUXR1icHXa
Au+siceNtue0jGPSaHVubK7JHCz6OSbyghdc9oYFDJ7ruBkQ3Zd1nq7K4NUbsNBqdBHchjyqxD+H
gYKudCMr+6ytgcOkVV1YpIajl6b6uS9S2b5u29Ht0HG7TZLQv3bZP0DQAYnxTscq4pb3XoCNiROk
QudfvWzaFq5emGiuiZj0vAWGLCx5VwlAgI51vL922/1F5z3vW/uIX+dHM6TWGr1rvp8OVx9LVUco
gdtIKLBsedUQVEFCY3cUE3l/WwIEfAwSN9TGeWPB/6gpaCq4PCvgikJC5n0Z4Z80feTi6hDjJfp0
P9mTaMFz6yYP40qYFZEFMfwLP4KYN000i6kTeiKlhSxUcvP6IU0zpfGx/c/YpIazcKfLMloU1DAT
UZ1qjVpSSNCSE0JR8DCwzAS3dP+OcooLUcPt1z7NpXKTUsEETRnuWwnca69XMLo9rnjv4vx+41LC
ocjfbEpaBfpIPQamsO+sQxu28NFvvLhRr2AY3hI2B8hkwd8JNbzTFiE5X8ALttj79TvjmHIvMnGW
De0/PDq5YESZXSfVIrOSYWWjrW28tNbByp+YQaIzrMOM8dSPqMZu3GUxHiyPQmqVZLf4Mbhj5ZNT
LbSD9vRGyQ4xsZDHBQkpOfc2jFrbfxqqmMxeB3jyrBoGbRXPneMS0UBlEyPmSFskVHfaSUXzcm72
w9IdEu2prBM2HqgNcHSZX2oGyddZxfskbrCg7AqSivNfrf9fBmm98sv0HEj/V82mZJUsFy0bXyKG
mjin7JcZAAH+8F6bDNXTMekd+6rvNUF/UP+5y0O2xQ/zpV91GqnlawVs16i5KHqVZNh6aV9aOjqq
rY6C52zDoUTpGYf/pV1FH9BYu0gQ+xERSevVQFZDCsHuPt1jkQ7yYRQsS+rxYG7t42aTSPDH68TS
l0mch1IX875Th3Yko9cyR88LqOC0KOIxeQBLUQ5v3QEdZRA+84etE79XKxCMgfmqoxK6ljIZsyv+
AD52l15MbT4jqCjrYVG1dxZqqEpOzZxlRh6A5AmZlxiFOIiHVup43GX3xyRN1RLIOhXfOWtJhRvu
RMxBEaWJyMgBg3pZ4Q+DqYY6YkJCRVxu4EH0UkRw78VZoQ1m+zTnL0fEdUiqLF6HoiycytVXE8Pe
1r9yg1NGpDSkRwpuH2g7K6QeUDqSI0hoMo4/CkFHHeQfveByhhNqUSoljhX4x0V4Kd2M5ADBv/DO
sh12kjEWGT6kd+a2d1bg6rArXv4h8OYI7w3SXOjDwHo2BteSU9zSodd9mExLAmVMCtPD1lTsV5Kg
+Jd8+VkCxJ+3EAdtdr3em/VkJLPKMIGQE9g/5Rz3BWhv1VpX/5qAX1GFxmVd67jgvqAfMKMkP2dR
21YHTMKcz0kslYP7uKRv1BiGVP9FSKz4yoxqUJxugsEuVut6pLqEFhHRBLaJU0WUAtyqe2goHCAV
Id9/yhAY6sMsTAQADJN7aRwPXMSeqQcPBhfJcbTZxDlD9/fLOVJO9mNKpBO5GDByOSa8d1qqPvPZ
Fcsz2EXF14SFJ+QlbvPbasw2ajDy1bh5kSDNwoytMcb8aop1JPsc8rS6ilskY255r9SrMSrs6LnH
+MVPb+5SLAKY3UNNIFUpr768/tfMgybf/k2gdyTlX9Euv7Ot7eOq6iyscTaRlK2SdyEaBZLSNm3e
1WDCAJZY2NBScRi6PakVEx0z3z3TURMmWHbViHaGJSJZDyvuGoCZT6aHLRPPeKefH1RGGh3jq/rc
uND4/v+ZzOmh4sqdaX2vMIabCJIl4u98mHgI4xImgehVletg/eG75+N+6Jty7ZUmo80XjAnmKdbe
aHCtsg42qkVxnJzrYnGtvb02jDTuTdBHgi7ztdiHFsNFdxytX4GhHtbJj+jY8Ge74ZDv94ES+jJk
HhgugTvNpx7S1wsA7uipB8YFMrYvFZlLzaKU9Wt0C/fQQDdEEegpp2FL9vT6gAKlKgFep8+nvZV0
2uX2doxFqE1znI365Z5aaGp4iinpKa5U6LlgTgVvpSjWV9cYwuuIxqUICgtcusU4Xs/vpommSTcR
8S8SWTlqiS620UtFWzvKMbOXUsiV2k5Y7ds95Idao0L0iSjo7XYxSeaJUzfANx+RuAy9KRN9D0zZ
e/kipEIvAABS1zLvzyak4Oo7SX7oRuuAeELx7SFDSgy2RT2rsQN4HX2SZvfIRpsrcJcUHmNXkzhd
xqtHpXq7vsuAiW3jcteNrWCxOAxTgMClgxjsiMMKBOghGwyFRHiGPwPhObiyj9+Q/L3FxeehdEZT
7VPlep0iOnwvPLUXdgZ01eszuxGqqRB2AgqhQTPfOPuCBmM4aNNpFLy5UTsBWK1D4k5L4RYbNRG4
5jyWsX6gx8g5iBmGLa8ZkynlYHSMhHTPDewwAhsJFtOFTj54hSV3pZphcgxEV4XSnRPbHDJAFA74
WIh4x6NDdEgRreLz8+qhxoqgsAuO1RqMn79CFDXPdVphS7eaiepNDvJzmILf8+Y4vUwTKXXrBV7f
7T2kPN5BTHbdnQ7vTimJ9wuaZGmSns4wqjb6Auj5He2IRTG8l4WoyfC+BVXSivAl3muA66YALNWG
6dQtCG2dqj8QFF72dxQpift25i50QH2/6IW7zbmClUGCIS1LuySVbO9e4/Fm+ZKqs/9+KlhrKORM
wpJGfIqLRKhH7AUjl/M2zrGwHdKLqeJdu4YAQ8+3HT5ZN2xo22xPkyffkW45lZBBa+mJ948gVTzc
XsQllN1X6/uewukrT9buSi1uAcljYrYFzTOLT+am1N56NOQQflUyzRTR6DkakuKiFNihGa25egVa
L3dX5yIjkBQZHRfVkPnA8clrD6UALfkBPa8GM7VW0Iqh1/tgmJOq0SLpXojLW37PHuL+6+t8peSX
5hZ29SLrC1tUudxIEH6uotWTpyXHdmoUZjRPbiWLIp0nqHQB7frtF0aiwi8Pp7Oxs9RVHGhr+P+H
808cmJzecKY/tjHhrFfy9YrroJmqeDmLw09S0/WpJIirz+YjGhg+ekRN5rjdAzg7QvlcAgDlxybJ
uRZMiiaDNaTLewzJh3t+pcbX1tu2bgDD4UOGfuiNGltYfrQJ/46lpJB6lIw8P2By+zElKbWX60dd
vRSOHJpVpjRcFYG6Fs911CVjxcsT5mveb5NwRkUNztZIbmSov/EoiDTL1AuvHydc9n6fBtI+ySBC
pNji+hgHatJ0QpJQ7L4mDVuWwp+OWdLBKcsSUDeXg25u5i9Po7+BwbEfoC63kloiPM4UIZ+tdLx9
bhPHG9PPMHM6S2PFCR76EfnAWtbgPxSx1+PtuWtsMgnYGUDmSIi6yFsmLlqhTySusiF6sCguarpS
POJJuM2fB+aUF78JnQ7lY0Ikh+20lvePEaQ61wjnARFgUPPiihLcqqJ4kdCj6i1COO3SRoIVozaZ
y9DyjCQHLKoyFvued8Y4jSWdv97D0N893oZDcBf9f5Mutr6UciWOtT4XLLBMk7Dk+zkG5+Q+Dr+a
7uSJRkN0b4Ra+KWVtetHHda/vNu/ss9ia3OnbsYu/7wGQL6P1TRJRY1YNT6U3bVEMxUTtQSBBcJn
3knt4blZlmwzEHVnmgZsBmYgZ2Ud2ZCyr4nfIzF+VnABR1hm0/vgrlwYuq3Ifzds/yTdzBwhioTR
v8058QM6AoR7zspbczGNHOVx+rIee91CHPvyoJw7Of26EOVz6rKLMwttHKCklG8T/u4yH2KKZsAF
ssUm7vZ+OsitA/z5NI9eSfXOhFvOlyaXrF/P988+PNkjJ3M3wCzn9MDzTC/5LKuJce1SaxSdHtP5
crGR5KWc2WpU7Tl4EINr3thyvRHGYsNk8M6SSVIv0JtlJDDNDvdiHqs/SUcifL6Kpe7FczzTIRoU
Cv/BKvWAKFpydhzzqz6poFvYBwwQXYJXXBiBQwnrxJLnG8gjdDd+QNASTCLLJaYbDhSMIhtYggfs
7EiIW/u4iaQS4mGiHs7omCaN6doBAs2kVQomxjAP62st5yR50DQK0PGDOfGMohSZBco1aaSaBsol
pQPr1h6QnFdcFo9QQsSrfhcKEfH5GV0ks/MGYVdLSuG+ONQJR6rn8ZOyXODHigTC+wkx9WoyZPq/
f+jMnjwr3GTAxPad8mu/srU4cLSzpCeqW36PxrS/w7v5MsweyqjySrcDUVnuZrIDNkVvKPgNjorX
2BJATadOnUSzyZswbjd42QHZwLXEKgtuyAkLqeDrM0qCgXSbYmE7+KjOurrVxemREWXkV+hW950r
6zNh+Vw8CqX71VuFN6YHaJurvWA6LnEFgqdKeDarxqr++8x/GcXoxdjzCiterBQba+OkmqXqVJ1b
tbLnSo+JUss5fhANjjC3qbsFKR+yGxBB+KBqu0MkVcqabuThW78BqsAuuhzIJsQM4fmS4qFQboKR
oyw0HblOu9d2cOY9Ahkjb8QklxYx9MMcJI3CYaqColQvr23J2IF8x/hjJnc5DakhaHd4srgFXXxf
MGtGTJT33uDzGUdKL1gDY9pY/QpaoeFGqHSd+R09FmVeAlcO/1Uy0rRxwiLTMh6QltfmxAuZKOjQ
6wVQueV+x+S4X+n0bpQ6TGcaCHY+4+qHw5LmQPKdZxo3Dm9rHnDsi1OO4jXcDRMlGiNxNWYfhN90
TkLMQw2kYMroRAkZwqEYkDjpy12Ihi+8LV5SWSCqqGa88ZVpAy+FLoD/SkCq4VyVJwY6zZlZXODx
jb6/S8HzfvtaMvkI/WueZQRwx/CWw/71XYWrDf3wlo5mtBFGp4vcLw62DujRktgkpw9YMx8PAH4c
wtn6SCgrfRU1iIQP35xwMV22dFdlomh+QAUZaTO2jRXxtMdm9Q7CSsJfk0ePeLmK0XZZGyOyDg4I
tIO+cqLuztOcFFAdgh9c/tCZmwHpGdtJ1HOY50Fup+4eYlq/eVBldkBwZqUyTz6t8LhpoFqzfOqI
eP2UVkW28py1fnh51SboJlRHNYpYqIoSQYvF9Dlj8ZqwzIob90qIrRjeY2bgMHWiTHNIRBQ/j7+N
Y+eZCGcBiQ/gkXUHgsg7s8ggZq0ovRgQzYVqapX4EOqgmOer0kiaSmYvA9aQ199jhB3QhksQBmEQ
ZZbyNaemL/dfRpcE2GIZnrLCs0RCI993J3RN+DuRikzHjFX51lgUBG5F+wFJwB/iOfKGw3h3hD5S
Uc1X1saDPM430U6UQ6Goa53iidycQ2ScvWk82xM/UIWQXwuFb7tt8/UCWsh5DoSFPwOZhxrshaiL
ByQsqQmN4soKKnDeWxu0dBeelM9RQa5J6YJi/n2PPtVKtYfgnl8kM84JHN4yMLONIJsyBKqvK0LZ
FO8naroCWxkLxBbbrvy3/mz4HIQYlm0eXbDNKdTqK03h3eaQxL2y1ZWtHBl6wd08d84cyOw/2Yej
Uofzjlv9sCcE6TN94VMcmMVUA4DoPLkKOCQPPqtQj+vzGR0EpNZp4TQwUSzwwtQhud6E0cE3MR+2
j1lXNTjffCNTgm+RCkCTq1uy+jLnn2FtX9irYBsWot1/T5iDJ/Ygd8iSnvVCiRJro2Kq7PMouLlM
yEYm1DqA71//wPIo+EG3gi75xZwxzQizmESS2urb70AluDQIjJPgfmJhG+fl83U2ix/5VtLaFsWk
EwN1ZZ45wEACSJ8+7Y7IOW7yg7AN9f72Wqzj5za+Heyi2pJZpn38r3g+ViljKnygzggR+O4fyYq9
FYPTL93afIkFIS7cqwEm5dHL6klIf+LgYlK4gTmrR2VajqKKLSHvSG9V6btkw3Ctq/ETl337EReH
1E4TMrXiAcQuX1u167FVfk0SWJe+5wLWytjmSPMBOdJfNNyjPWmC5E6AWOoD7brORNrSzIACsQUT
4S4fbL9HFbRRA7bDYJEChBTUtBR7yDwlvicu/rfXEOWexYNYoDRF8W1Q1jxfej2r6ihDzgAkznmF
S12QZuWX76vl1dVObVZQJo8GUJYDvVQNSP5m9IA6Xn7iL6PplNIJ22vX8uiNPOwlI9vgXKqhumMP
WMvToCxW0du/p7BwQS6TXF3wlIvbMLcTAqIuqURCyHeT5e7GnicTse8TGFGB14qCTUP/0ItleJ9e
cfR4YRLKImyW2fWIMx6NLH/wamwS7SzZYSO7VTOnS/diYQvK4XnZ1u9HlsdxS5wE2dJ6oBskXZao
lnsCEkf5QIGSlbpHswFuRHBN+jm4f1SiElEAuDTAOoV6JLAjeQP9vr61FVMSq4cmu+0mldax++O1
Oc3+ftVv7E2VX0iAX04cAvFWD3/FTowA1WTY/ybuHB8WRSHSxMB/c2APL1kXewV1LXKxM4ccDqqI
54AkNbCSmJX59neQ94ix7RAV5h/kDk/40/2er1YzB+UWaV7ki7pHTsXztwzjYDbPMiR0Al3cB4wU
NXYPiBggE2MyMFWR+Xv4HhfEn9+dEiP+AbfSk+5Zlx+GJmXsJOSl0MS++VyMOh2aG+64Lau7GmIx
GOIjQHJaYutG0IAcfg0iodzixUkqQI4B5TlZ9xeMIrCjeUIO3faDpMH7FaUl1brUqbvYgphHB9WT
i1lnyMU3PtIbIMj5BG8EbxUYlFmWA5dEcNBUM7FNuqLU4x+Tz9le4hpCoR3fbpUIniz4nM+aHLn0
AM0h4GKPv3YSvNYk7CCR27v77hypwvCN1JiNqbwMdKmQGRqrR/QqZM6e+o9NBrS70VQkrRiN1TuN
/KFRYkq1mIxWho3ox9i+LvgUFeQachIVnhJBnxubmROqJorM/As7HGVSQyCt7UeO24CY9xrUCcPc
yxS84uNRvIhmUEhU5ZYOjk7pmlQ4pSeBmeTxsvC1881qWo5zGAfxgiY+D+pK3ptLXtAOPfC4zyUS
njCmdMRnIpyCNrgJ3euUW44OOyWzBLFO2yMSJ4C078E47+HNubC8+eDkpNSj1zD6JBqXXo3qW6d8
TzPFP0lj5YRNP9O+qIFvRryG6lZSYSgFcSE6tjQnJCrUEs4T51er/razbQJooXuzjz2ka7k3wO/H
wdd/8jIEF2iOKbDMqJbGWmcJ3/iYsN904zkE8s4QFIDI2V76EsM11FuZ3wWl2IgtiqMhG0pj7IY1
yPnlHn/RnTU8cusXqXUFuk2GPQvY4Vfwmfn/s46JJweAzpRM1/NH3mRXo6lycKdv1evLRdqNkluA
pbzid9dRBsf4myBLFjOOpAIFww9iWDll4bX/8R+ooYhDUE8cbnRwIVNBPsWwdK8qi0cwSafCqfKU
vtaWWBhh9mg/1qBbARljFIwzkXV1A2fjGd6kvFYWhvmLG/NDtStmL+sTsV4Qi39Llb0JAWV3nkk3
GYPdepu9IWePm9Oku/gz7H3fkEeHpeGKRIgaw+0jXhYQ47rlCNojNuJCXcHDy7xl4cSyprCEyhgw
81z5+/uq+IacBqnwJD9iDlih1m6Jk//HEM/XZpamzIM2VLf4PNwSl+OKdidFa6eypIxaqiajTGrF
hBqDWAmaa1azxjegEB7iftgKbmLcAFja8Fqepq7rGyi+8ymvX7uPGH+IHRUtvPTNMdCGoNPGbKgo
CONslHXnsShDN38Mm3WdVBcB66eXEBzUeI2byf17QEVCgRWWgCIm+ACoEzywb98PdFCHAdeJGFha
bQxRteegw0uMa5klJ8sHLKcllmndeZXilr0vCV/Gd8ciXFet7qlsrTeK1pHd+8z5/k/3GxZuMX+c
giBGyGuzxe9fFvRRiuy7qj/MsJ0j+30VDt5IvHYoPADAt4gVGKjyD5v5IvuiYJq4DAUZv+mk159t
ZyAxkPTgy7WVNPUsaKDslenDRepKeJZoc8bljekLqt80YekcT91Vwzrz1evJpXffZB48lHGqNQNj
Ku/iBZpIhNN3l/8D6rBh8m/kLDVsmJ6LFpdNeg8zAKrUIpY2BbAB6Gf+VP+frG5T339ckix4zyZk
RtxiUkI6B5pNkhvxVRkdmQkn0EHSQj49WMMuMU0C/q/o1UePQ80ZURg+DtihrHs2ocbiYF60zxOY
RKulwfUSONm+VVSgpCPKpYrQXL4frt2/0WDMzrjQRuQAz/h/MnujBMJwbKHIXykQj9iGUbBVglIX
Y2qpPDRWlgRPNQP+9YciQp3Mj7nRizoP/acgX7+5lRDhsLxXz+gdJWLRdyGj5Bkft93yU5hR8eFD
yhrek+XxYixh1z01Objo4CrVc9eXo1kLLoB3MUVUbz/nm//nC1R+/iB1cY9WvSLM41bFOBK/4NPR
OSmHwNmSvyiii6dh62gx98wK3/yqLZdtgQsKYiZ9ypOjeFwwuRrWaplmt/hvnsPV3uw8yQKvBTwG
0g8SW0bsoeNwABM6MZgXStW2QGzW2j/E1EKb5mQc6NZI9NINzGVB4AG9YpDoCAfT3mbeJWgaHwlK
iY2kFUtYfzMbggnl58qH9ni23akor901QPTbTEnf0YikIZV2OMW/KPQNs6i/6o76GWcscxvl4TQL
v7V+19kIKXrSbz7/uXvKOnlXvmhx2gcHx4sKD7pSwJivfktZfBbXIRZDQ7hpW2n9/YozOyPx4NcH
0K2NCEuv8IqhwpXAoPychFMB+FkqZwcK3bdhJLag/hSJcZ9cEprLd+1hYUD/otTDSaMDOViRsMIw
rQlHDb/3AEI3EtkQ6mmRyOd7WR5HBF8T2JRvVAPBOxaahMDhS4tDgEmd42t9Vj7Pw0HuztXVj2mR
Qb0xQew4X4+JMSXfnTMOrdeUgoqlCbj6vE6WJVI6HY1Ft3EZiFn0AqOrbW8lBeqn4/kJggxvyUka
FIFvlJAH3DqLAOCy27vKmaIelUEeW567+7he8XeCrgzaAI1vwBD3icoetnNri7/7Xg7zVo89s70f
IJDSfjsNq46HypEKpt1EZihmX9JKt+gxs7b4T290XKHCTrO9vY8gBtHKKIhuPGd+9YQpMnCm89K+
c29TrjvBYh96JIbeaiNEUkf5GWs1RdkpRyUgjbG7od+wTXq0h3MrorCNW3A7dxvNn+xbyQhAHRka
1+BnHdvtC1wJ/Fk2auV9jqLkI9Qn2oLSDc8pSrdLYXAxYl3YTFdT+asTBtNktNm/O1A2cruwm+K+
mpS+zAO2CvGDOrrckeiha6OhsTtglFqNJPld9ab7dIFNSvqjp+daFzemGMekCj3RI8331B3XbCwn
vTVGev1EKRF6qJXZEcpczMvwd2UTkw8vTLRe5SBBuO5zowXllhf3L5LcUw3vUkekmj4L2gdid4Ny
/H85dtIolAJQi8ag2BscUdPVDY0ibx8djnDMPMAwQ8v376AOKn3jPjAuGLFMCCwXu/y21VEsBzsy
GdKX1QN67afoiH1KQyiQBKReDK9N1F+YkiBm5Ru9btrK+Ue9yHf74BWxlxAfZ0a4lSQe4AgB9Mbz
sRh9fE922xGjsneyPuUawRcfHVrojm4BKidFsslqotAWN1uaMP5lmj+d1eKjXgZODKRtuWhoalCF
M4ph8m8hgQLXaWlhl4YPKDLF/hNzdCo8ZfIVQ2qpS/kyGsPCp8FHEzTtiYv8liV/GlrqnwM0I7Z3
nMQ8ICqPoY8GKO61VTDa06JBqcgGs7ZW6XSqcwGzhnm5ny2CjaYKJagYGINe46gFjegX6JEWMxxR
tD8I2HQ/maNEEWmEDo0eg0Qtq6i++VY6+zE4KXIBjgqBaAdj4Rb/vGbcZzRP6vpTtkgntjY0AvUl
7Q0tH6wEe9qXTBQFEk+qDVKRJWMOReqsK/52aAw6PlP5UVC5KLnb1CFr9/Scr3inlLWd4k6Wt39I
bQDFRXdmPUyVdTBWHNbqL+/neh99B0O1niR9bLhqNwPm+xGCWXG08sBAVfnqaslumUEGNcHKAzoA
hiDrPIV3Uu2Om3tQtgMyS+zGG9vEvM6VVs4MbXkx5WGs1UI2ezSRypazfCYBM541oDvjPUdD+OI1
NJVPFM0c0Izdu2WUBDfKkpx5a7MjxS1anBz5/VSH80yGS7Ln7m0b5Hxa7x5FnpTxzyYc/y/7Tl/T
UWsxySPXA8UcGb9nR1IpgV2UIyn9zbbyCWHFb1Wxy4pVrdYjeDOmytUeMIWmqLNdWVLnEZvKjSBo
U5T04zaoj42B4DRq8dsRWfYrdLrEpIxhSkXSbBg1R0nkKMfPjof7DuDKTUNWWPXYtbwwoRUqTeaS
dA0U+TIIvv1Wdgdr9p/tvcrLA9DnmK5kUa4M6ocqV8prjpJo1LqRFf2q9ah2keBdg+ylhvS1cRCX
fO9eFKSG5ejYdvpVv4ObY43Kaw+sFtnFG4wcozsEDccJuPc9IHUB5oZpiPDMKI3YDD3IhGlbjNrS
5AQ0veriy4cHut7vDFcKUU4MhqPvZwAwLyf6SQ1seFF8Oot/nFsANfRbGx9XAZN8JWxRud5aBr7n
c9qCethlauD6hm8XsO6Y2OacISOYHqX5b/zWOrUEoWC0AlK0ItP9pGLUe4n2L+ViQ60C5BNTnBgw
msxgLcmBjb5LYSMwUH53g6dvnHW32rHHBhSwmDYq9mAHtJU/o5ygGzQ7oefrh5Z0SmRnqjpniCUg
TN1Wd/g4cjDiOV+7DSK8Zr2AtS4IluHN2hj3EvDTorAhwZYQlLphxul/eBIz7AkBvFDKL/DbojWI
ULBcqxVoh/Mztez3c9wATieZO0mQFhNUz4wEktg0pugPGNlX1NinsUqdCBUR03mjPSONPlimr5BN
ZU+0WM6/6GZwFTfnaRzJfHhL/0rQ9zPDiVB4SxCjxuEgK+gofJApyp4fKV3MqINrBgkVI6UuI/r8
ZhzvBzJhuAGOhz8m8wCkrrlLXi0xP3Gb9SyboA+KpIMDP0RyCJ7xu8NipGeG/d+pkdcWiJ0vZS8e
qjLWt/ggJpHCkrrloESIvLCjuZq4hW5MIxc+WRFcd4s/p6aWGY6qbtwJbNHiiRTd0RMs+aQ84qJQ
5ZXz2aJyIYTrFuTFH3Qqvm+eUqFZMokAy7t19AhCYmoLcFi3R8IvNO+NRnMHc2uVpkvVtEA2tmac
jhBytEUFB0AYAKsMdZJpGovnQQ9FSaQk8S21HVur1xasQ8QRZkUDEAebsIrz4+iHm3F+4KQ7LHWN
yXoTUPMCDaHOcJnidpfvbZZkONNO7LmYMiILn8EWD50pbczLFzVC7Jc9m0+HWAnQDH5SSu3qSFgd
ku5wdEAnlF8bZ5pss82pa+hVYYNYpx1bNYs7iCwq1JxoAvms/nw7Lfj5LLW7vwqAi2Y9IzOZXlZu
QgfnlQKm+3Mt5BnnWrXdHFw+O6hK7EUpJM+xry6MTg2UZRcDV6lSxhVyOp2KUGtBWtXij8WDcLqw
DDlkSv020w4tQ0ir8BV0S2NFAFWj0rZiZAzhC19qGdbz3jGFIQfDPulho6/v9/9guDggBam0UdR6
zU8UkVfQwAQZ9vDFH9piJZ7Wv7k29Bbu24ebTEBibZa1vmu3Q6bcmiRWgPot5nNDQLdoCVPPshlh
+KwRND3O1fEIE2u+OReIf6bQ/4cMPEBTpcW88MBcL8MXnymJ5vdNxy1ZgLvT1RHECQ0TLQgus2CG
MUID0PjvdfNg3jo7F8ndEhaV6lx13r8QWc/bOszq7KQAAAzjnYhtBsaihWuZ9bFUghjm/0N+S+K6
ABAvpb8l7ziuy9H7/7bxOCerZ/BWJHx422cC7lA4XBllSoAzpWf8ICDYIGYHXtKXk3O9o8ksmfUQ
GdqKmaQS0T657MiZPzLbYHbh6esAt2PFSfnWmy5YNJd43Egy9VZ17hBO+NCHsVIC0PfBPIFnf0lH
hIxOIiMuSQepoG9gj51zjF82JIMClD1zXc8kWT0i2bMkTrrcY5mhOCBTsBWnPgoWeEfzCsYA+g6Y
YT+XZ4Ko4WSD/I0XRUzpanN1RW8TZmC+2EF76kDmfDxypcU36qkMPL+wVh6eZOE3LNwOKhUfMGl9
VimG5Jx4rldjYAcEhHKEinmbgQ0lBY7yFt5n2yeKcJmOktk68M7yltowq36v7y1y/NbAKp6dwMam
zrAa1PKz1vnNSUFh9mK/pnTUX63etuR7d9gnU0Y3e+dGsQ7XbAyOVlnrl/HG+9+o68WGVzYYHIlA
BCixlZT1rRTr0NOG3P3UPkU/VdRMzKOGDoUmsjo8WA2wjru1fEdq4YVBym5CdcgV8KtM2L8cHBi5
u8g8DPD0el/DE1WkMvWBD5GD7jtwg8yqxFKbOlzP725aAqe/sK7A8AG6rr0Ye6pWr8VEsx+6dLS0
9g7Qrc7BHYXUfqq5rn0y+TD6Z4Eqb61ye2nRAOrUnuUaYblzATZvjGtz2unTVIPqwOuK1P4SEXkp
5lkDkDwLd8cl6m4DVtN+GcAGhVTsYSdDmapFBwPhWLovzmcbdrd6uArgApzOvo4lDd4peDGL9Bh+
d63jMb3QB5Qlxkg6lbNy0eOlO2k7LrhImO4ij0JDY1wmV9ix8g0yeWVcYappvuq1U21J0G6n9BEd
FP7E4nhxygVrwFMbSZAzhp6zGK0Z0QJCLIDDxBdKuLJaltqd6Ekic+gVMO3UteC1t4gvF4hV0Uyp
jGXIKNC+/Ujan+5S9E5CLajHjewt541JyLILZWFajb1ozve9ZYMBQ6v2Xjo1xKaJfreuShBHh/nj
rZX1x6VXI8D3GNxMOcarlDHltCZKlYsQjSBiFvhEMVeVdf/KBTzUWriRZF/DI2lL7Yk0Vtc6cOzY
VjqaLnL1Duz/3FTS8P42rX7fOnIB6pqADxMVtewc8rJaia0mkRTZASCB1mOeF7qvfIuBnKKKeHyY
XC7hiKtGP8UEf8EhoU/uL0yOAGrohq6FS4rtr4TqlPDXo1BCxJFWHUOLGOuTT56N9Fq7HOOoiyje
xT1x8Yjq6B2LhMyyS+CohF8fFRLsDEsMpNDN89p3JTXuqa6F7lIo9G3tud/G7cRrkFjNoQrEa/fO
CsXjF8f4XlBNL1gzO5CR2OEbn3jX7X8XK+S17ea35FphYiRh02VIMx6hgVGM3QZzkNjrKC1kVAF1
qO9Q6wNNbzY6hSAUHMPKKfiJUeI2ys0uDomEOce2E6jTAnKOzK6ytIpxGnJYJmB5+pt7WL7bDJJZ
H64YFiYb9eDwmHVPGItA/AL1xNeV5R7D9Tcjz4S2bQUiy80G4MvdVs1pXtn48qRoh9UGywtbCvuG
FRBmFb1KjFNqYRjMGQDvGoZ4cuSoQWjSOyX+J67BPuHRmA36WQC5OSZVePOTBAU4S7MTVtw0bx9i
EeryhbULP6KcWOrY8YutGew6Iq/UD6x61NMwCDHsxaaQ9evinGsamF7xGMlHGCQ7JKog7gOZZ5Ie
vQPhHg8km16zX/AfPlGKhYbpuIUPmmWE/P8zWTntvZKe1vUcZbol2gpgtC3DBWntdrBfKnZICNd1
JdJwukLJQ2EHwxOmbPzxNTnS7JZGIGwKG7ErXqPpV37LMmmtCqZNWz3bcs7wa2RVmVSVDxanMbfr
LB7szJeNCrbIWIuguGe6Y/gVZAySNCgjkir9TfzFgnINyHrp43oUS6HT4k4z5bPN6vQeJ0OODxZF
4G0ZMYyLc6CM9cPFH3Tklx7EOHi454+Z4u+NdQvUiuB0/ue1eP7z91IzzwKy0eq2i40OLGmdEt1G
kcR9FfJ8IpCLnSjWUfrmZ6Obg5cX0vMqacZYLu96Fuix5XuRfv0eRT4OlI2fqc/qquuCHQCN3t7a
DpEgrK6f2rGEf2CcrswBZwG+NLB5y7iW77hGi871r5qidzR4X4TH3N9ZJ2hX0HKevCPY2ACGY84i
G5s95FB9PJjFKVuIIsdniTaGjm5rRPlJk7s8IQqeVU5+q0jLUJjHkmgE5hfM68plrM+qt/GWzZ8d
ME2j9IiZWp9E85elhHjlHgzbl4aefNDV7lGGvKi9RyLywkoFk1tjGOKi5DJKPsT3WyC5mHuarz+4
nExF8pF13zTZoZ+00AvonSYMhCq27z7fD5yPWiMskpWdni63GpGWvnLDLFo6H/Jz7irIu7OSBBGe
0JKgtTvQZZWvVXymwYHmuSCm0B0yVgzo0zDPS78/VoSWuH2vVb5MMp3z4IzMbS2N+ClqE93/ambo
Shedwj8CCol8ftUnRcAByp0uAbigHuHEIrYwD9btTtxSERKqwZowEL8btd/7brPRGGGQ24RPdkl8
fpaX4CEofyH8KDOAE9Y3Xp8XXrgkxwfjaPViAsp8N3Z8AqAAOkNoLpV60peOP1r5nNQraBdJ4zyX
l5n65n5NckmVOqh5D2ymjG8TRzifDk3lxZ3l90230rlIDsFG8MsASiEsPksY30nNP5ZNVo7V5bc7
rfpuKers3N0rtRd3tLVmILnmLCvSe3dv+yaJEUoqIeGQue/qcD9ly3YxqcZevXpBqTvLnA4Za/Kd
u4lyJgPYL8dbHaVYl9jAMh7s5xN8fYQoUgCsQ0IYF3RGGa/b8lbZBGTma6/IaF3PwbwNmyLSIIyQ
i4d5y1ckpGTEe5hnQAn966l2hcWCwTgLgWgmQmbJ7MKmJasCNRJ7bFa66KjyqmpsHwx6+Mb3Iac+
EHmSbonTsE1MG1+bbvJi86nJOGlvWVw22Q3mS4NZg9v6AH/uoSyn4BKIeRHUJ4oKYtadTaQr+9PV
DUhz2RP3V8vtkNvGY3YI5bJFP07LDrcXDbd+n9SQEanKbIUyS4S5xgzPeKeSTgWgIRq8rl7kXNqF
mSBuEa4qT53NKrJzyivqQ1axq2RUgNFeq1RvXIi85uyZlpRWRNnngpPgFmxTXkLTEx+PGMZT1uNX
3XXQUuExmqoruPSJrWjHZxDrenOlW+I/3abWj7AzTfHtLCO/lkCd4WjhS1da2G0OVdbeNWJzmHUz
9iLQSzaiDoeeKfy5cxX/x8hAoJMrg3XDPqLIsHGH/mctdt8aES6AiJ0d5KVFsP4taHQbJqidbJw/
7q1MaQlNihf5yMSKGTZ36nRSqSN9Fwoa7CqpiuHlGtKHY3388ENdVijHVQtugCZq/KSTC/EQGkrH
6NVYIs4tCaZ5dtFKBA43F8fV1VpwZHWOvJJGveTOzRl6wqk2+jrP8R3rxUq3IHZu2N9Jq3BaDKk6
hOhdGqW87Sqbn2+/BhJ1uNoD4TTe9RfsWWO3XsmTuWczp/KVF6o8hcz1RaoTsojAwH/+Bdxhw2/Y
oCKOSL2TNAaSs/O7UO+7Ri9tyF1mRZBhvkZP88SoFVAIdCB3val8qeSmFLFqtF2mCqUBuCulijUU
aGvndxYFaAu4zsZQIkbaZ0HfKniT3zXTZW6TU3wvxmsw9PriR8V/KGQcO/a5fzRLvaL243nEI36H
svxYY7j5ue3ivCnrPdC409l+gIRrbtWYqLv936szH2hy+Kt7+MLUT9gNi5lrglMaG+oINxa/PFH0
FHj96VeiEf68te7x3Pgkq2YUlUSgZYT+YQHy+DXhL5tn1Gbs1olFQPauKDFS7o1pbmGzUL7AMqQ3
Y1Tvz5Di56KtTezBz2UBp4FzuI9bcFK0Fp3w2Fle96UtRDetewZWDJbhOG1QsC9S+LYF0fTzd2/w
vuR/fJQOAQfpPzCEUz1c+5QdK3r1/TTtn5Fvzfo/R++DJoLWjsj3Yl6NS2kvLXbPNG8KUIUTPrMW
3Ze2Bj8Csfk30jura5+FOhhRfQgxnrS/oao663L0giJOLmzrId75w2sl0OarC3G9zL3KlcpH29V3
LbVhxybm0+p22ZOrRsOVyClmc04YEzKN0IjPynrljkbZy/Zhd2Mu+c7g+Z9LmxWqFnfwkBs+MXYU
fO7kDQimz/QkNrBZjY/NBMGLjWIuim6X+llRP0bmeRAvlaorRuTJaK6hoE4+ngRzSdFP61LIX5Zn
ACJDm21lu71ZPn1V+PDexvYe3aUSPYT6H0Yd4kPCCGmEbdkjuADR1140XuWT3FbiA8Bm4QFzQ1Ld
lEgPlrzpe3Lr5yEyRpsVUxg84XinvZodibGkex8skBtX+S37zuhoMhFzyizTuIH9pUO+ZtZStEWT
SGtSfymSYpOUDFTtp89H5NouOe9ANgjBmezO5katNGmPLGd/4w28wUDSN0hwsD1nGk95yFQSe09U
QOGzO/G8NZlHSOm9yDlKsn/+6n3GWHjCzqogRB+DvO54LXs4pYg5yOLu+kKjk7W8zM3AzC9NhDtA
/C9SOckwKUwqodCDa8M6WwpdVLM7x0AD2p1rSz6RVNE96C4wHM6EZCoBpej9t2RjaR2yICXqeegp
FfDI2J+AD/Xr8ADu6zC9Wr/rqxaaz1x6EsDGDF7TXxTQCL7rcwf0Jlq1VpSD2JrZePxpplqxvIZx
HZ1GF5qBRzPcG7ejvGEjrJBynXMVWbLG9Jfc2UE/yu6VcdBr/hp2KwRirXq06Lf5ALsPC2Hg2h9f
sInap4X63gaN4o5jz6X3IFuugXIjH4HU8qLyhyMPk40bTnsQcKJbsbnujCnnGkeXSz5Q8HDv4DQ5
JViCQ541symMzablho2wgDWs4zDCfOd8tNC9QX9YWaFdYakQWNTQHigMtNlLepWwZwPOklfXP/bR
W8ocXr05KmyautQ9yEu5whwb7Ro9elv2Wngm0qc5jXXY5jlMKmVrkU8R/0/V3LhQtiir3S0iFpzy
2haR5wumNmbMSwGsNw4qnW6+894hntfNl3qjuQmm1B7rmIsNfkd0rk2jYzMK8qmKclQli/rz1Gex
oN68nNAsdv2gdJl8fkCuKMpeRSw0VB9TwLlkbiTRAJrYEMV/IEvjdCD+DwvpUEq3FSBesAB+toZm
bdR6/oJOwuTyr3jTDmBpOqqijmdvqLkXKDUN4YP8G56ioPvjFtO40hbkOgEv3BZ1HWeA/jH4Sp6e
HNjtmezef6pfSXdSWsWZULO+E4pF/Bc/QES5b2eu9mfKeZmmlos8q8U5iPp5hbge0jqf+DTWWsgq
KCjeBnR38iZURxWfN7RzrS+S2IhV0+lTKgi6oK/nWqu6KrIcz+VfyKz8J588NcaiB/y4BDdLplB3
isObAlfECHx03b1WCUAdq3MigAiddlfM1fijag/qx0PO4kdEzP6vU0FioIBrbQmxeuj3UmWWYc4A
mmN0PNrqhwgMxL1SIiR9Ju0kMwi5rZib7gY7G3UYB8crpTQcaiw96W3b4pcFRZD3D2KGVb4dCd4D
6WZQ/2wS6Cx70w9YNFP/6Sh3ATQtVdbOggpWG3Q3ThhLtvl1eZFTuLM4aKM+ab6UsnNubxw7a/OD
Y3HpcM6eYozQZdpeXDfrpDNxAtpCU/sPrFySpaBpDAKh8vnNNGjLE8C6BBuwAf1Tl57IU6jFZwD5
rwcK/DW2/+n3KJBAh8ZytDVfUf6srY2PgZdr/ICdn3ePxv7RJn3g8A9kqTNItP2FeVhA7Hxw1OA/
vxYpW20D6Dx7O7VYsb9kA6sPgPl/FAJk+1LFtr+BDkbmT5tVKt3HVqWTdj+qnmWfAw7aVpPHoc9c
jTJ0UM0fEP02kQ6gJnDsDYBhRuLa++m/N72ip5UREhj81FZWyq3aR7Xr6ppEbPHyMjjhibqDLJZW
DikUdmLk+dsf4j9dUrXDSutiv0RsWbuLhc6LQNw8dveFSzsh5lAbWEhh56a2rGCBGp4vA02wufDt
FGPrcXAMGlifUHFaU7jQ0RJFNlib4+FbpbppY7N0dllT1B8oHQDFnG/lOv8iSKO98vfv8xCQKAAc
qe8lO5aFnDreab5xibiBPYJ5niC/Hkf0npvCgFpMnBEgsvNzEeOOH3Fekavys6s4TmCyA5xaWAVs
hFDCRkD4nTS278PK2jJsRxU51ZgrJgwT1eIiOgSJITcBvotcMFAOl0zYg9hIbl5/tzIUY2kkkbnb
HW9V1e0DJ2QGWz4tILj7x5Om+R6KuJnsIOykMffDt3X2e166fSMyDq2eYcO+FWEe0avK/MpWpX8m
TcGnCxJFgQGsMukiiwY1suY45zJXIvOXJJs9LuOtptCGl2e4aNq+BgKJCzjxsGjSj5liiWNhIre8
dVqMdEzVY5K5/WnJ1qJNGW+gJlUab99et8a/mynXaCnO6z643L4JTE55uxkdx8497un03xYhzAl3
kGIVGDk3Rr7br0PEnRu2KJn7PHLo/uWk2p1sDP/rhSqdJ1pA6RBud7AGkWmcZBdqKk1ICbVh7OrY
r8/dSP6/jz67HfX0Wv30j9no6XQ4HNUz7kEy17uCSXwX0hdyqDdb78LEkYwJJ/bUNxogq5N0RvN9
038FY8Jy5oovjJU9j4lwSTxuo22Zz3PlcIx8f4ETVExiCqj9TK+Mu0mIHFahrtNzzGRONpmXJ6/k
fQqbEujMdJ8AXOJW4B0QqTmjFq2scGsSUHElW3IRfqT6PNLD8hEadSRECG3x+JIGG9133IGZgMnm
iwXAMdVpzlYPDgN6UsAq+hcVYfEUkbWmIekNq9KQzH3DrNn3pqh3BYrJ6F7HCoF0e6CGP6EM8WQm
nIQtUZeivOcghXkm1AnDxFX3vIStzN9BZ17xjOHMpkq9GiWZmzS9UEgPG2w40NIIr8bdLXVq8Lnk
EGtwU6w98dBhelMQACn9GbYB+0jXiMBWVRVM2pDW7UxtHLN7rpeOSyHu/n8E4907K241ji6qXNSh
ZJseFH/SNQ96arUAME7jDy99LYfjEYa8xMyNOftZLEGclEjDrb88lBqDZBQGKvqj+7I5bg36vSH2
DX1beEOQu39WzgF4zm5X1NAyDMDJYJgbdhSc+I2JljU/XzIh/DXJ0T73u3LasoeljqUhVHx1ZpJh
klj6IDbpy9G6QNPZrEFEm9V+4l+fbcF0Td9B/6jAYj2nsOdmVjRFa6jR4+gJ9QXzeWfg0gUMz/Cm
c0QoH+BCpfSWYTWM9cZo0y1jHdGeJIWc/Rgp8ITgW4BiY53vU8yJzsH+mUcj2LVIyjmMLhQiokRo
fZb/kwYIRR4gbrQv7/usCe3fhmo9kU6Ay0HYPadJfXm/YmYCXQRjBemNEDgfFuGT2zlt843aQ+HO
J+EJDc3JxvFp4mptfkM2b7oUt4azZ267W6HS2dBheN6Ik1NbuJPCCbFly1qvlLw+OMDXQeYaYMpD
2jevQYvaBfT6Sj5XGAoQ8RlVWrOWTsZQdgu9NxDY/xBpO5RDY6ukO1eEeQ/MRcdsEgWgf+31a2ol
e+JZYXxrkjm+HF4LkH+XsckLm9jfGC0tm/Lg3kAeCDgLObsRdgEIcyFZs8lak2zg6xUk3TSMaF9m
+R5TSP5nMbh/e7AtfPkv16G0uqbhCaPmKKW4cHFa0NNHGBoSod9W/1rjvvMEi4iQ3lMxu6nYQiYx
hKyayclmu5mOKpRZYu9wdKYSvQ0mAt+Gm2ip5w1PrevvgU7/dO2xgQBg8auBwKOZwhCS/DE6SyIm
vdVxVYipFal9Z6svv6pYE/7zOWAqzqU/Te6RcjMmQp5QquXxxxRnkYi0zDn5BKqr9QKeBCgHjTjU
rPhgwsdBxVklN/DkxKOq3IElv3BtKT8H5e1X0WRfwy1DQXqMuLBftIU432XSvGjV8rnev26qQV7q
DHRNEgYWC//RkXhKx+vZ2PVGnY22WyFmAZZOl6c/z7STwAE3AD594fvRozDV+LEC98klppbY30S4
CziGXOeOyWyd+O3maoOgOOWSzS6/fgLtpta6mpgykxc3myoypvWq+N7JdpCvePM+rLi4fTkifS7v
BCg3oD/jULhIgFLJHLAuJxvpvpm2gY7Si75Vl4EsAa8pMivqHyXiYpJmackfoEl1dzpVebHdJ+T/
pzETgtW7anLYbs9sMqhK9OmMLr3BwZSXclFqUP/S8+6LW6HZ1KomGjKlHcGyf19ilTb1pi1Nfk+7
LwnsPI2C2S2tpY/pNJQoyjSOduGMGbrjaqQHCx8wutl0w2WHhhCLV5Um3oQwVmG444BTYFe8rXbi
wuqxoNzMGZmWF3ouQg4x+zvynsBLRO5YhZuAdRbzXDmQKzGcGCKjXzj8HRw589OyhJ7FF53NjWz/
GuMZTgA0HhMQvxeS6aVPhXRauTCFdAToZ+eEtnJeexXAFtkrA03NzVkP5Aq7NEYSA1C05Z15DtQZ
YGRWTJwZ0CLd8c6E8RaSRTRSzO/bCny3fG06d0+ZpL3FhygNwNkkp1391exChFf18xQSXtGsflGY
G95vXQTmz5kmBW1QCDw3R0ix0nWu3ZTDo+jqqYM/Nq/Iuc9LXT6CLj3D6AJDczQjfmNAxGtf4XYr
h5eSc/zwF0kRzlQXtapYA6E3NmP1J+WdexJ/REJnpom5fMCi4zUKocRqUe0MIZf/KgsneAIwVbKN
NRjC/Y+6PXlvRjn4dqwomYtzAp4wKHqQ/nCTW+2r48Kx6kkjFgVmhh5XfB1xgQT3QW06zdhacFol
rEZysCpelmY6+wN6HZYDHEkClaqR1QO+pvmdPjWgW1iV02H1QdMiFqDzxHIWDRqxXC3dobowSL30
UsdH4jpPQJbDYdcyEVmtLN1YPYFHxy+o6mexIOHlP2QRAHG3nQo59pC5jUIlPfllNud+3TpxW0A3
UJoE5L/J9fQRjpIhGVDxWy4nDI7JX14Ea6q7KKTIgPj93yhh/XTmfvfQ5fx9eqG6FKc0AAZZ+q35
lqeGQN6MW8sf4d6b9oZxuXtvZUcevWxnEIydhA2Zr4nxnJh49V8fzs8srbvpX37t4jOBE/hC5Yrz
V7BtZrqz4t7WuHFbBnRc38kjBO0kYEK81yToCcPt2ekkTmUEeWECmjArj7zbGQ3og4fpnzC8koM9
/BC4Y9GkaMgD2u41jvmFvxf+zad41vibJea+sXG/oh0rnGg9FeKFBTVZD160QDHiM7RZzuhSxfNM
pKLPUhpHOEwDbyOY1ii36Y03vbM5IUKv+onyOWPamakNQxl4Q4gXVZAodsNzBVfg5kAwmnvqzWyF
aPwLaeCJZ3lWQA87fqL+kyhKUChwZVOGRhMuxCF9Y+DTuoM3pu1B6rDwX6lNGLxbowkR1XDpkm70
w+lSlgCtoX6FWaO4vqj6x34IqCVGhOs+sO7HOkkjQgEb9leYzTm7/1q48gISaJ5oeQDziMTVsTCd
m+XeMIEprzRNkTHll5xjtFiSqce4rIiJMkxlOCtsEhPT8xyW4KFGK43W2G5+QcN/hX3iFeOGu1Q1
qZHEdyIuDIbQoxw1drppx4HZCLw9cwj+VU+2nM2GMyWoB31j8n6f3wJT1zyJv3W6dbnAo3vWf6zB
Kpk4NO7f8LNI4rpfpnzkyZQXS/SBlZB+Hc7EEG0haSjaYrdQyq3leURBWDXk2Ydna7YVSnqAzZx7
X1JMZ2iFaaqpBf+dxs8aaoPyZbIIbJ0x8F+IKwBR2kTpS/UQp9IoGqY0GSeX97wky6fSft1uLJ4p
EjmObpNNG5Tgl3U+2+YiBIZb9D52PhA19Jkv5an5PaRmS/Bc6VEtIMPwlrMYYBg3GAFGSOlLX8yC
/L8tFXGU4+MQCzsKSgJAQxC2Yyq/ER3/6LYZhO3ma9R9bF9dhsdmmpwvHE2jnSC8lIQ+ryRWNC2Z
KyQNhiJS2P5QNc2Aq8Hepzr6bj7OJ5xBDS8zMfskRHzjagkD7vsQVDv7OSqYl1uIK6ORyIv/uPhr
+8lcM77NhbtRL8lgRca8UvyGbXsL+ecKSpfW9liFNiSY84Ui93QfltiO8xA64HTYalfReW1oRp8g
bvcOpgMCs4Zb7XmaEjfd+6OFoSLtE+Ju26spZ2X68YJRgpuD/y1NSvgLHBOBDXfEdPT0xTWuJ5so
pK8nJ4YIJ0kgABlRub4W2odYyKde3UJ7h220UR4MXdVoszLu0GNcQENoCdQsCqRf5rISAH1Gu6Yd
mGEaMDpdf92M5PMlq0P9Ma96kPcqNp+hPov68bw9INTOSO7KG4x15qcnxAsWwC3OrNBrp8xVquhr
J6g1VXyrjylRHcRNRhf4mDP46EU4hXGmR0yLFY0CR53lMvDeFo4hNteLiA03JQ4s1r0K3D6laK7k
nUyqXH/RKOuR2nD3e0wyVweho+wfKLae0wgN0wQLm/OOKLSi0RklAhuPiIIDvxQia9aGC9moQ1CH
VquN0AhBCv6xyjEe70QV7J/WqFkgfJK6EUEFWki4IWmn0IObvebhBi84w6Vt6kKNzWBk2dc47ShB
NnvDJc7SSBYVgGZoyFNetfVrL5okj6f6DRQJP66iJ2I26jvu6M4HYpLvYWPvxRzc1DWuiI/4jiJl
VAxwBKlvN3BJK/9L0XXaSNO/59el8ezA64yYxrozUEOqcJtsBb4OPyDpXtkL7qISY5siI5BTlMXY
JUv9g6mnXVmodFdeFJvzKjG1T75nXlX21+xXhLwMYE8w4SJaiJPskPdlA3soX/+aoJtMfyunIfFi
wWWeAIb+cNKI3bCK+Um0lMdgghZGmZ2d09VL38ZDJGBz3hqKUDUIluZVVJZaC1qYfKeE8cWkZjPV
zZaysjbBzt/eBqpH0vEDY+joX5Q5+g4YEzM0gXcSwItTQhIG3K37tXFrxXxnCorLnQwmaCuD/m3E
nE3sU050iS1B3aNLYFBlC2OSGttKE32v0sEORe0FvqHQb+3bJDtfWXjxlzYPrKWGNGjriNe5e9fK
6lbLc54j+qi7iYCh8jkhxlUzyIjNBd6GZb1zhm3v8KBP9mG+fbo4ewKsZ6Ad1qPdY+BOEm5gG//W
eJ9HhyBqgRqwqepD3n3uEMfHug3eukvI8Kh0NXIh6DhxE3nmPpmSJb/8yi5xR36WJZe4tnYasf0e
yL5F/xoeNHG/IwfNaFbl9mLQXiWEcP7VOsMe3tRPed+pdFIyPZbP6yNQBdNC9/cPzapXXVVQD4sW
KmTjQYfUfLGiQlTnVkjK7bc3dc5dE4grN60vIozzYDdUm5AAbp4Wkp5QJudarPbi1Hsj2P4805o8
sS4Fe2qQFs/qgVWmtO02ekaXy7nVeowSuZFHc6pzoWXrsjCqg7KNP/52odt9NZITzoKOmtCbK9Rc
FajdKOdQZHgdHhz2JBPKrrXjRax3SwP/V1QkbTozY3x/fbP8a1mxYkApl9ZcLPD46ZTPKc3Y94MM
ym7J3O2PrmVF2nhlD8Rsy/zEbJunvmb6/ECMKzaLI/DREF7nmnJJ5vy/a0FAsNKGQGgbs2Di5wUG
pDyJsLRf1emf+1tK7L3n/J7d7ABec3zrqPDKkzJow4OAyOu/bM7dPzei19uZCxMhUfoov4dxLH7m
22UXShx94JwbMgS/eaveAyH68AamTC7wQRxvmZJD2v2EAnRrZu66hN2f9r3SXf55XVMFGpY86GIT
1lUIo9ie7r9FV9/mTQam8AUDUIDrOBFNh01g2XjLHbuE1mMBJPbtJAp6eMpJT4DJdE7CYjZeKTG5
Mth1mzE8OogVA+gujw7rseINbfhdwPftj2Ufndz0nM/p6usSBI3DUcZAq0FtrIbiViSecFAo24C3
ABaanXpNI836eLwhRw4xHkD3rpPJAW+n8bAA+ibAOLu20+0a509aE/j8ciS9R69BOKfZvk+TrAI1
HRkV7+u4rli0KmrKli2yPtQc5eo2w2vNn8T/2KRZnE/F8ndkXdDKLOynFdEUIitjdbXMVidoTZvk
Dn+/ykFs0aNC5VfwSPNoEtGfC2Gp+TXE4z2oMVOGfc7C6KK7quiIonG2IODIW4J/ZZdOZ7A6qFEU
2TrPPaeA9Vau4AKb+lwGDxt5d7uyAX54pMqrs8WcLo6G58DsxmlaS/x7/Xke8FE31+6/g672L5lI
SSNjP+/qpdTty1UN9Xu+jvjXm+axIDjIEFE+V78pssevs67gzq/NOziVTBAoKYgTpHTbB7d5nD2g
iKWTuE/Aq0G5flqWMx9IRYy3Yie1WqYxmdXt2ogJGjCJAHyW9hRdL5xG/KTKHPl9lD5sdUcvQXE7
w4Lg5GqhUum1388mVP0x8AmYvWnbpK6yKXCo4GSUmi2HA7bbc2h8EBybTbKM5x562CcLNJdjffne
YGtuUGDDa/s26OtGrRa1lmYZiDNVLNMSVhnCUXEaUUinitAyAFfSg9CYS6ozJDnIkRlorA8EBix6
0WmBn1nWy9Mv9F6ZUnw3F9ATMyLO5T0rTg26stilbPpj8hNqoTp5Hltc9FjKOVwKQwcyeVlBtalV
Fi+08JAUHkJjU43hr9+zqdYALkO9pJiExwmnYparSRi2kC2grdjeg8yeV1M5z+ysvHaPXaUhIZ4W
luakEa3R1hHdiUsSr7MVlSG6+8hQ5bpnTysXhFqjgx1OY7Xv/jK0eZ/LM13kUIBdYLK3HfqNnBbh
odQ+rqVkL4ZqFMLbSDtJsJDJmGpo5P/sjxotlMgFDkXT0eIuc8d+KOVxiPbvBs39RwDbjgZCacUz
L8EVPFZTdbQU96L4d7MB4ZSjiFbeQ+/KQe2LwhopYNeUe3H3rEl2vPr5eGR3AaLhiaX90wodfqCw
Yn9o5v3t03OZ9CILBlIwox33wpz/jEddsZCg6krToXiwf9/w13RiNV3ZUdlQq/0ImPw2f62E6tsf
nzWVARcq/kirlaIOIL38GO/fdAEi9nyNYR9PVVmEZLZV39epStUYb8s511Gu39ypaPna1EP6mP/3
f+ux2PVvCql01H9w6YdDUuEem85ORmh0rk/eyixkkb5xXEURn9qQSu78/IezeszqDD+5+XLAeIYO
SP1d/TEG8twvjg0/OQ9FreCImSeo8+7o6L/JNb+plbIrpCKIR9G1G+z2TsmE3OmU25DW4hpg07S0
wyYfldmkEPzvFkIsZ5NQ2gz6W0fCPbEkPwQvWrGYIeq/ALlErfzmGr7d+XYq+ZE0pIIOkeVJfdqL
oNjOdt0BG6uViPo5YA8VbA6V19LqtngmVov6BkXkXAMJZR/7vcvfpxNjzbDEU48aiSvRYJCkzgMU
mlEKmvd+ZNZwDKwcvXx0urghuiAcgEJaJLfukZr7iKcfxlxILxMm+hkpiSwIB3vjNsSZIOFC4J7C
sXnFJ82FSNC41mhg5OqZC1vxJwNJ6w8peTkUevopOykS0TMI5c/fFaKsN78bf9Hzftd6H5kWPHON
tcVc/R1DCrG9gR7uPUWyhBjz6JlM5Kv2H0BQnLq6Xl+eCvq+GGD7e89HmEhvbOsQZjMcYU+wn1dR
LKTiuUqzBA82pASfOhl3UTblDnaQiah5TdBzoA/qs19H/qmS96WZjHONtY3e19mAMXCeKFzXBw49
pGOusFnKm3fRhuPTFaho1Oq7IWXhfdT3x9yhrzC6KDmjwAPUO7+uQUsCRl78i0g2f7a4iou8flrL
tQob+ik9DAA71aoEIe5k+4JDRF7w1DG5UYdiMlNNBVXApf5EWqVDLNMlKDR+wMvmQVbJxuX83JkD
SwUd9aJh7udd8F3f3dVkoHPBT6Zt58ysP00zrWnq8La8BepaOgS6aeWUckRUUgHVS7u7sx3EaUK0
En50AQ39FQVnNLcwJtcY5dvRM0q/IyVm7yClaAkft/p7HmYQWVvE6vRkZT7A8ODA77e2YqRhFyni
cjcftbqo+2QXMy8i0/5zjYgzoD8DgEf2En6ND4zmzx8gCXqU4v86rx0ZE1q0gR/Y3v3fWD00/y/A
Equb5UbXCp3HR0N/UyqRTQreE4n8KbjQrAxRu2axd4KU8KvRdwgonNUmb5Q54a4HvTZi7nKzsZTg
bcBI5kibVyURAvGk9+jlxdRFw+J+ya9XE05J7wWpeNfzmOd+gFy76so9XxIpV/lLCpxv7C0B6KWh
ZZgTHqPTYZPquIoAXbXo165xSUe7Cg5nyMBw+Jcg1RTSjQIMArcC54BiiBSPnOLkBEdWBwlJRJin
qcxvBu9FA/fGUmK8qCPN83QrC3aQCxTUEHW5rWmmks6IPy6n8bAiEHtx0HOW4wGYDCtQX92ObvrP
X1Y4CHVKF4ST1gzS5xqgdIHdYmx1n0naf5Chhrm8MSa976jZl/fnuWMVWaave/KfRfz27MMERymQ
AjJl4UZK4Ud7F4Thh+9dSsskMzzDU3UnhWzSH03vrko8WbxVR20E1U4WylAD075gsh9AONsaGbTX
NdD7hPW4RJZMjiIiw4YnKZlMCSikuxerZFD6RKeU2QMOFOYzr0lUT8Wf8EIx5u07UyZaP1P38nzs
FKf4cbtBuJofBDx1YAmimsB+wIltiXm4tf8PKFxsh6MZPUX44QwAAwdQHGEYa8o7VfZxTbLND/KT
W4OTgSJlbs+SNVD6+/4gn4a/SVagDtUXw+a6n/KdFvvFr0u7rHY7n1MsxmBxSrz6mwGB3BR0fiC3
UtJ81WA1qJtgXxls4ihL2Y6mbaJvYpc2s102/JPYQ6NVzjIip4vPke1zcol6yjgSGIqUrbH2A/TP
xszVlSuzEK1Iusel0HqR3r6aMyMKr/ja8zT1eLEULN5ntjPpenpbuXN6oX5am7eeRS9BfcO8lgpU
9bpSDWRA6NcxEZGU2ClxpR8Eusdp1W1kmQcwLmXueIJjOfPqYhysFynHOlvLxWR0JuEyC1UQXa2O
6VzXou/DT0HxgwoRuGFduvlplVpQr5lQY5nrxRfUQTf0DdE9XiblSK+k2RVX05grZU1N4dV0QDU+
RR0DH0mv/g/216N/vJpisOrsQ6zMiw8BCMks5s+UnWuEWtRJvSd9xKo0UguPzY7snqox9tm6rxbv
TJT6QdIDpXMiofiSkjMaffjQlKbvn+hwdrNyQQ0MiPYoGGFYEMQteHgFnKwtlPmeOEE5wYSIrVW0
/OhSEWTVJYMqgg564owp83jrWnuLBi4B/KvlX0qMnSy4sutbzh7yqOvnybcMqXVVRiuBYVcSq2ya
m0/OkO7VBAodmvImbGg+uKY5Gz1dgaoDCWbq+/LLzIXVHo92RE3QDeZf0Nyt5Run16JNL3MO4w49
8vqdfEN77/Hq+gmhvD52oECIKmVz2sZxZbW+MxgtHfnIus3K/fKc66XYU9oDe1haO4VkPSEPUEgL
6PcD+6RPPSoeTtt5b2VlrQUJR0xuoaOlYkZNDob9olaxSDq+0c5PkSeLQU5NS8XeWKE16XAD/KpV
QyMqIDgS1jy0ax+SHg2Q0BeoQ8NedBm/7SJvB8nLmSS1PzoYBjmOiYM7ejKe5w3lzlNU81VNxL06
Kw/BACvB2oaGg8GaTQBDCY0kF4eBNVqt3nHx28tc4z7PCCwzVSyAPPYW3CfChBOrqp5f7gqdk2ug
tnQbIZwvGI5OB892OR9KfuRv22clOa63vAA8gS4l3CqU6Ph50fcWNVNhin+JS9AtiY35KGdxSUhc
tnBKFQq/7fN5CLkt/fnyWNzQQGm6mNyYbmBJ+AUuN4CBQ0Nno9rv7EXsz/+LM5gpX6SUSdOvLake
OZzxfzz4wdB8FHNc7dUAiYJ6FtpOTadIQcWSeggSvmGfuA8lpz8IgctWWlf9V6KGjDOzwW5UlxLD
vYJbexM0WBV0QIc2twgXOjWEMTO78EHGvs+A6tLRLeeb/YW6hAJOFx63qg/cVVa5qNKZpxK54qnO
by9hvsTvuj7HHiVpLoSs2QHAf530xABgRj6BO/zE6Gxxv7vUHY/iJHI8w3mkuxLXaXMbM0gRyP5n
v2VrFKlkJWqnU6LlqoJOuPzYqLhraSAoyZvw1fcIgItGDu7FPC9MAwRSwXyW0IDksUt1/q/XZp6G
u9nJjd1udVVyTsm2Ukkv7T/g8Ot3A7FuEmXZR+YTaDIZxQFkhBwed/AhrtpDYwYYV40LuZ4iyW+f
KnnqkLLIp+e6UAJFo35UybQdylYjew31gd9JGjECOt4zxHh1KDt/0FtY2wgGKmLWbe5Ei6SMSWl7
jvFoBeKnqPVlJnlTLcN+9+lsxzhS+AP61II/xc1NEBb1pMcEZU20RPbSvIlrqgDup+rqPQ8w7kTN
rM1TeVvx17OVClMrQfjfOK7bINFsCRVjb+xEowrZO63MSMyIItI+Db5VooUkle6vgNklntp3fpqX
AouhCLKVxw6k2cQ7wvfA6rf7GTDXsipZ+597FWL74gbygDKT5lX7fPwgbCUeCHd3KWpG8jFhz4Dk
efOIf33eC2QvjyuoZWr44NlVh3UgEoQWvPxB99woP3ec93nV7vydj1zN967TuvwwSqc3GGrHu1jq
k6LouYVeVA7/PnOm9u7CFIK4+Qh2ekqVj8gvBvhA/IsZhkHhZaKZ3LYso3kSSY5BJnv6ZnBUWhki
jtscQpUZxdWUHMCJlbpVTqQ3heeS4811CRziguXbtWQv4RxrMuFzI5gXdRRGmlEFsqtlj0h1Q9Cc
bncJ5Chbu80A96AX78B4oISWtYEbsC41F9QfdxidlMqdrcVFSnd3CBFjtiBo2GvVJO7eRwp7aAC9
9UTAx1+PdtMkIaU0fFDrBJg59yQslqJFomeJMvWXL+kre/ZfAJjsTLAd4/fxMeawlK9Qja0vbnAx
AvSpnsWQLGeeBucNcJIPkHUmgmaZmOBycEoqwvknViSCr71yDEkL06PsitG3O6qoJ1ONWNZ6Wm5p
894ajApyQ+x3GVGYdbr6aR6vGHFQO9UT/VOpsmC30uiyLkZzW6RvLga/lX9eCKgsaFnIFyPIkCTC
TWGqMQ3m4CSLYLbGF7Ghrlxo/9JhzmY6tkaIAVvz7IcPWtAJVMZeXz3ytSvfhX25j3V9XJ1ikYC3
jph8I9Td+BpWNG36nzggZGaWH1vMpt+fzlotk0CXwljlnbmzD6OOV1QewgghAsKlKYoGUM/w8ic6
LFEDEM5DoL2aoAR1TqlVO2oqljIKGUvpr4icKHe8/xUe07dwzjh458J44IA8coSg50BOcVymlNCX
o2Cd3qCPVzkfCL+dSFMq67Fb5a0FZc3O7vCfG9Bl2zU3B3TWrPbFmZ1grQvi6uigB5QoAOHaOHbb
9Iz/simu+9OCOqZMXRCs+aRQu0n7hynvcXK8jH+9wnDfar1gNskLSPIM5NLe/c4JGLlcrz6zzhgE
namXOrpSmnsJBIEf7cwSqUlvBcSyYS7AMER5nZ/JI8ZvOdsx0v5EJaJG/lD3P5XtmsWAiLligGCl
GT1ERrOlQ6ZCoqh+WHo1WFDYDRJeut14CLmLB2ZxRo3aEKr+g3vA2lJafsTUWkLImA+gD11pszE5
Z9m0h01co0OdoFbQqkwo73T7sV9azBFAVskX2LCucXSUsIhpIPmHzTrGe23bGp8u1WmNkEQ1wGuF
JQl0k4FmemolELF5a4mcWh5jnpQfg78qb9TMErKnnvSf4i5aqFhqTkuauspDlxCop5IshTpLFOUM
qpy9LHq0iTctKoMksS1v89fTKWuthFCNNhPQYzYekAhLzAPdAlKHwZaSCoywdB4dmwXcjb5EQx+o
5+VKmnj9ZX+osgGmnvrAe37QYIUH5WtVrmFcL33/jeFu6CYIq9LTFT0reuZp6lp2amKxoE23BRb6
i7A1wC03Lwz7MAqNc5eYdihbXeX0YaOtQL2sCpa7elWzN563XTU3URPI54hxCCljDm0pLahxIJAT
CAHfmGdI76RARUoMstnWrHWj8Fn4x5kWVAWVdrJW36r9rNYe4AhJRtG/rsD9MeIK3tjI/9TSrhDB
tJLk92Mmow0Gk9qFz3oLJBQcpq1w8cqGXeCEfjiCdaND9r70k+0kuCu1kHmoobEDNZUxI7a5RUqw
M48ZfVzc1qCO2+XybCeEUdiVJJvr12up8fWWwf7Vatv4+ACCUuX4BYdKD4UycSSFtoStpBKsVmiL
UA4qmvaB3UeSQFlfR4HqTXQsgUi7Qrc0EM4qHaEArFBllYPHorZ4iwMD8DBzdlg5nY7CsaXrAd+s
ULrduiSqKJVOx+lnBQ6Uua/d8I7ajQzhYjGe1BjJ+TqHYub6+7taCDpoCEalj8U78KEQV1w/RhrU
58CVvU8yO+9MpCijqwFQ2ZmU6Ok1zcOZ4BL2NyDpSAaJt1nzVpmubU8Le6bRnNbiWndvuagyaXzR
IiiRDyklFhvNR3YqZnn2QNJ/Nos5ge4U1yLoZW69XUv2na8RlJ8xyXaH7LmI9n7I8fqu6wF/0aDT
5e4ojYLGJApRMTHCY+e9VZcc0mreKUY9n0cjjF8+3sj8Aia7Crq2XgcOuNtvqcKlAgMVFyaU8xOy
wgkb0VJYpR7vstYh4yEtJHujlqm1BS/AwRWTtQediRJFJbNDnNQmuE/KuzUG5ZDRZaFwI1FPQ2Lp
sKeZm0gwYkfg2Iqs589+eCrY5cYaSS7qKWhb2VHselqIpyIMhTo866GdGCwN9vrNsx6bYvPpHiYS
ObzkeTDysrlcZhFg0/JCp1FV3ZWgpfvQJsT3hUiNU1S7JLe5OeVU6drNBdqlmMunnSXCXQT3pJea
tmqLrAa9Pt0SX+mGHH0l8l7Gys31NIkIbhJl1ZOgSfQP21Gu04V2+QIPwOFYdsYnCzOLh/NkgzBJ
iPe1qpxFYPJgyDS6d+lhGCac82mqRF5rBJdbEA344K0H4YHKGaZW2Onn1xVhuG68nRb73QWZOaWj
bS3zfoet7xldRbBaKOS/5VLH8pTqd+HymMQqb/Y5uh4s387qPwmJK32b7JH/8HCv8c4eilE0zvSP
iBn+iJkJ1YJox3mkJ5dDKFxxCqVs+pRqMEWyCDYX4POv6OvC4tbkwUrkGPYGNaiOT/MBLj2C4+GL
siglD7z75YVeUT5OQKYfscu/MPoG4CeDRhKDEiByhtcZ5YUQleEtHFOrsQdA35sAR00JQWYMOITA
pUZDt2YhiKCksYFtnbH6OsH11fCoZJzpo+oH+ioEN3u9/YQZ0UnXldHBGQc0imH33JuZ9EyRofNy
Rc46MPgoH7gA7NNs49KWW7pa7aIwOh5ZnFrIDM+mmCdW5S30qOCMbUjhw4UeFZxaBZb9zySkh47k
kWtAKcNE2PKTi0U28nIer+ym2wpxaMI0J/JNyV9xxstd3D4rrCk/tLXUARCVmNbegECcZ6lMtsmQ
k8ng2QP7Ni5u/gpCGxto6pjHCHLbDW68OH4zOtNe2vLULOlhxFNH06PydHf5MZvNVgnNai8GhVIo
EDKNuDjCGujZW9oZXFSgn8Wkw+cFW95ReV0QvT1PMR/aO2DxwC+D5mlfpV2nEPBuZLecznpPQ9qo
VWINNzv5NpoCEZG4vGahye3psJvsujWlrNhDcHY2DS+rpyMpR9u+/sJ9eXiTNUfc1qV/6oLRK9d+
HwAAi6kA6bVv1IdM15C6MdDLaX4c2uAhdb2lTJmqAXnhLKqoIjv4I263VJfhMkXXCwEXQJKtEVuV
pi5J0g0ufMyZTw++5TurB2n7E4SoJTALYdaySIVGFCYLQYg9OexGEOXM8XhYNd+tT425ael6ohr8
kgrGW8lhrtzwsMyhGZFX6G8a4+B/QyMxAri/JpOstDwaBYKmdfKI2rvF5fylPfCPpQNtp5gYlHQ5
8jSXEQQqpUzjN67j8N2ZlU74UJwYFJAgiAgbR9Wy97rvGlF2glqquT8/VSJoJmd7L1LUT0DoFr89
OKbNyVrHIfm6xPs4TdJgGwzt2l6RGiSRBzNJJzM6GFop1oM/+odaXHCQbVAAfu86uf/qTurc6NXs
A+jCbNq17bhozF7G23VXsiNx2R7GZ8Spn9uBlti9p+3U5s66ViVrCSv6uRALJjrJKA3/W7EkDHoS
NiTMgmijO92Wpf9gX9+fuj13k3+Ois9zIehZZ5JwwNIz8UlEzQeSfOrIk+Ng5wmLzJzHwrvpdHBH
tl+1n9yOLL2WgWC6lmgYeu9SZ1e/d5iC+Y104BSDZlT2mZexHSfjb476puic43Zi4rty9/abCEPH
vXjIJ62sRlqfwyFZXXA+GDHoLXd++tpdHJMndUDUNWAqvzp0YDz9R6ixZ4AMlWpYFORqCmAacTfM
KfuFNzlDVoJeseKfFR/1v8kTvi26DygpXbVlsOwEKgEvtBKYFEtSahVuxESCqavgFlxuLoBHUxBQ
MfRSi48sPg82e3Ozm8mbqwWIJQDEC3F+gefYKvpF9zMCA95A4Ax0qwaS3fZ6SFL1ejwOJev3OKpw
K7PQ7qwcu71pcH3PbUFjTRVbV7pBINdSAPptr0ZHRss5hJvPbrSpeUVvzc4ozqW/zV7dB24AmLtB
98M12SF1nOTlRHkIn9HHz/nnFgR0ahpZIVZLaVOudNsGfHk9DxaRlDEaJzb2u+fYBJLpxvNg1a/b
GZE/TOh70p2zh3xu6ZU+gfmcTOqOIFhRMBL15fN0h33ehFwh1+UEI77GRfnD0XYCiu4fzaaNEMGu
hVGWqjG/6nBBvkLW5eRv8fh7A7uvop7jXb1YG0twtgonIS4o6a5WK6qZim+B3ioJ59Gz84NbNXDG
UUCOPqntWu28kzhSa6xNHcuJrjtpeG4/NpM4g68gHMLP/W/VXOKKRaXZweDIUWT3QQd52dF9gdPu
pWmIsTSSm3W8CALAjHBbYLiYiA0nl7l5a1vjzttNp52MvI23yqfZT1ny8ncK4fcTVOtfUST58D9C
cFHQyy9RpP9V7lBiXa13ddZ/5IZGaxRMr2J0DR5mAe3HnzOJqgsb8/C3DkjU5gLmLipPJT/pQgk2
BUm5NryQ2e6NDzjNhOPTi7wmKrB3WKv5pYkz4asdygRBhPBknr/JoZqv+4ZEuwsnsJb4vwILIwKa
sFc75C4rBIMOrUPWKtjTOC4uFGiHnOCXJ9Y1C7PApEDy/j9Ss/ZLILxmw5BoAVvcYIvRqNqKJs5S
zqcGsnSXVgfO2nt+M/guIFewDO8OZQO+0FZCKEE5TcqRENkAZFBwip6IwFLsLS1lNN7WIVX1uErw
w33ssX7qWhnIYFDrZApl0DaPSALHHI8his0UufF7qnXj1sAQaByfUoFO4QrOoAJimJ6zjoTy5m6a
zulQpQMPQH+AprNZ/6Sw/mBbHvNJD2TZfq2LkjYPJ3TD9zPGuIYdzhcZaGstnD+fYRTnyG4mgAUg
aoeyuRr8lImL0oe8EuKulnws0xP+lDX9NtRI72rQMCmkbDd5yVNnuhTfk/Zkc2LHx/RjZZoCzvgd
PTBHBnnskkEFpqWzcoC4HHhTuD00GSEVkYBmSdjEFzxVKdlZhmGGnTAseuWY4//tKdJ2u54jiZPo
pBkv9LWbxPW37a5cb26usrW0AcwgE7BJ2XcDPZQjGp6HrRC6Xu8tIdw/qYWf7Xq5+hrbIFuU18YT
crIAEzBcvEnfq8QGv0j6v+NtJMfQc93p5MjLG+YmsODUJtVr4XGe9hVtHNEexSZSEmsKjG8hVP/V
57NBTdeBvx3C48JJfr4N4np9fS8uAf2xN0uhbxjLLkAycTBmoaV0Yb+Jy5cXoBUVd2e440Fwx3rD
LikpN9XwGNGNAXpku4bKTUqk7zM+RehdUS/IgBMjgIMQ3/xrtsZjXcJ5q9UepEJmOV6NjArSYrNv
t9Pba0IRVJlG9xGWQ7z7KX9ANJkZeLSyueVwGosKZRYFPBUnIaL7k9P0B4wpCp2mzFBFfcNkOVbk
HmmcG40ZUwx+nOfphf0364ovt/plAxeDFYEyGWGrigyYrraSqtNW0CuVjMhroQynOuXkUFn+Q4fy
Fw8PzMQHpOCFqJZt2oYfWF9wOF4uNpzRXwKBtQpg5q658H0MVI+6u6lctT6Y/aF72DhQYECpJKsm
CH0o6SolLwl2Yj8qWpawoIF7FMP033rFi9ItCw1OV6Z7mLyZ1qZPCfgbpR688c6PJwC6/DpuJ6Yn
omigd+dYSyDWkw2joTOghtZad4Mg9ekQiwLIAwnC3yqjiCJARwQ0OWykzS3pfrgNSB/93Q18yiUo
A47PB7NmLDBW9ntexHu3AVdJIF5UiBI7VPzRFjIlsHqqkkUZ2tcMuRFicE4boEraTf1vlrBB53pt
74hp1b3iVY7+rncLP8MyMDrBXoFMxUio9V5yk+sw8WPu548O3G7GUX0vZM41YcE+tWUCeQrKGdsE
rD/fVio6E3A8BAgetBLRXqf86D4aF0ze7iVGxo70Qep0OoA053NWlc42oM4TdiJbQrXWss4haj1x
hKclEvhSX010TLczq8qtZIJb3urvE5mCWKk2GtbubzgEu6C5ULWsR37GVb6MAOrsHdoMy559DU+j
q3IY9lptQB7TNHVypr0h9o0wlp5yasn9d8nrVg4plQjW0NQbLreXHpirE6mbA8as7B7fryqvtUS7
eaxW5m56sUjzmLcCqODost93tTl8KkFGAR93GZkuWOpQ9BWH7Zbe2Ovl208JTBEdYvGY+9PC6NJG
itI7mLt4lozt+D24mTCvDBca2Z0qbeQBj0cMcJ8KOPDp1xrzPWqwTR0je10bjAiaeVoiPBBpiZhp
/zjhunCv3K1lFbKTmF+zQWqhUFdApdonLFyPiUHxG+cfHUnbvIYhC/niDQIkzYgUQaMlV+fe95UX
/NtwWktNbTu6LFcSqJ5iEjgDm+tRW+QZ9viqi1Qd+lHhPnH1PzasjcTR/qLqrKsAAMpZRtBmWv9i
OL10IsMq1B5Jg54NjaLIq/WQvxXBFT2hqqys3Bd3bKj8EHyQmGHl4rfwM5v4Vs8VyC+3D3sJLngP
Oadqu2yhVYDRb0LMKvGVg6R6Gbt3V7RVuuHiD9Afpap1hwvnlWpuaZNV6lUfT4beuEmNfucqRn+m
3qjBo2rvrpngRl06jr6fUzeqY/kcFm/Vu7NRyWgizgXXNCiP9IZKPSuZm5wPyOySK+TL2h8kaQhn
4a44JpwvXZ9H9Y2X9ruPKtY48POQn4+lKqFEgd+kz291vGLon2Qifa3D4voduRm5LKSQ6qecashG
t8gUBb2wb/9WSxalWrNN3F6SxYQq+sKAPa8AAn82Cks0Rm5clLXo1IixxNvlF5SqjLvhM8xy7zZI
j36aVBNjziwZJQToN/jV0dqE7pMze3Z8JXzNZh7S3O16mTWVSNNfe1Ar5x0/9GVG0eh7ws4E3N6f
cb9/fuuCAtv4HFoWDw4sxiV57/JZeWqrNk+Rr/PYTzyJBwXQGGgOtLDaI2Eel1rjzIM3Zh4G3DEv
1Di6Byt/fPq2q4kiwGnYSCgKGW8r+diwoQWy67xHKA/PjOT9QnXlGsZM8u4tN6x1qPrU2aOI30K+
kI0HaBwh3a6SHJO+X53ch8QUuJTJCbudHWqxCPKIOIevIcWMJiexal83DWt90aegR7iP8rota8bo
feM0jlRHAKdDuMSwSNroZYjRSUNprey7eeoylo70EkpM43LNFNEjds+lvMa/rFd2LbM3oa5xx0v+
x3EG/48yGxZulqjBU/5cMiOcY9l6E4EKjR+lYDY0F7r5jg02+i4kkpWV7heK32jouCfWUtGZzvyB
bOamd+vuSTN6MVJ6JwWW1CX4DSWWyugUtpDHmF6Cf0LHxdI9I1tImTttFQPdvJzAoEcUYq8N5swy
G5hwiBV6ehs639yjS67JM4g3OyZ28dUfS2nk5qtgzOrFcO103R57wzJha8myhNTpy2MlMjx5R51L
SIpP+QwGTQWnkE0aIwp2Dlq+nPbhmr7p5Q+GQajb1s+jkBlb2nBQo8qWstgq24IjKNxudmAYRq17
TSes70b8tn4yN6NNkDd+wwoh1xROExZJgsvfis+EmatWqWmGjzHWILqkykFVgXAVPZsXvG9gSBJN
DPc3BFIT3PwbkiH3b8IRhIEO/KJbrGeDe2lQecaUvIPK4NRmveylQYx7yapK1E5B0RBW7aYFqQAP
KQ6Tvm+kXX2U3cqi6SBG7JMSllkxwi6/ehwl1uHy/vFRTJBw2Hw81QQLUcC5RaSHloc1ER7tyDCN
V35QXvnN+bC0xJy4bBdTKMZlu4AGkBEJ6JW3OAndAmrjPG9FYiQWLCc/jt9zpCH36iVGP8t1EUO4
ARMeQI0Q/PfPXWtHuHoJ2XElGgJY8r9t1W/V4i6zIXkbOJKrXCrCDDUQVaflzhMWMCFOYO0jl05E
5rinjPQZW9XfSD2TiFzZbsyR8wgS9QMOXSzxcVzJuklboIPzOh5RXcYsuVHV3KTcBCrSU+l4WbYs
x+o+q+S5AMvQGPOdc3f3IOe2/xv1EiZkxJhA0/gFi0AZFn3bCh9hzAXWjNxbIfTIRDkkszFFdJTN
AlIc8HeeGxx3CjzS2YPrps8BXBmgk+b6URajDtPUI+b+qLCur/xWSebQkm5bdH0ESX5s6hgPGZ1M
0ZRTr58N/RJaKBjlAx8GiWBxT0MlwEnSeLKGC+R+LOVZMwSm3CHh8N5spPlQY/Rpiur7y2W8h4/6
KnRUUf/05UwFgKeg0slD2sxHSbJsMtrTYObFE0A6uWMAlVDLS6j7QnVAoamLnmdGtH3r4NplsrTV
gkaW27oenUwT77QhUiAeBptrcPFlghsXuQ4SiZjgfZ/V+zoplehCBICAPDlrWbrnaBJmZlC8ZNfv
9tL3Ug30wYHWADZGZRojP5Wa3HSBFloG8H75lmsSfaXZPLF29wagM2lB/mZmTUO/AOVud5Ytfrqe
e8H5HzWX6qcdaVpqKNWvyfwAct+2miITROIouvXBbZ/CRuRCmj+VE1fYAaeLYlD9eyWcfRI0zgf2
QIriK3foGMse76h8H018CoJK8LFT/t9m7acXsTvLo6rXGPxO9Q4IbCRhUXbxd3b0ndHJpbjwlsTw
EtmQoDpAuF4yrSSKZuJMRHA1de+ppxXGOe6JPU4SV9J5TXtKkxXd/0XfbzGxGY3bntR7Zv2iwgUS
kaNt79g+CJWWYarDfE+Yj1EgtIZJRTR7NT6yG6Fc1tEQqeCxZDjY3PMbMMXGMOtniEzFt4bAm7GA
h56p2quuNxc7EVhll3EGCyuvQSOpIvXmS5nFRYsP0nZcTwcaCcMp1l8f9c4j9bAhxaUwjoGQKJMH
oSiaL1SKDX9QimcxDCMwl1kUaUGha7GfyfAcLEFhpVr00UdjmrS4UAePlNJob5IDN1w7VjRAcMMe
iEJ4XR07kl3R1p48qXHg/tvNJ4Qz2s5kCI2Cqd3qmLVIY/CVUY24Azeb2ErFwcxIR/PIq+CQYCKd
psGlMx5ErYlneQBYT9XjNJU4YsI2DWvdsBuafV/vuWryaf4/rL/MVmf+XWXenAgal9IUw2kzKWxy
vbI5izjE8IuOF0jSCvIRpCkIMrzjbRwYi+iE39X16DT2uxYF2xMqsavmwnVKa2wv41A90d/g2k0S
t9zsJSJ30a2hZHlkdK27Gtn5VTPdSDCKm3v6p3VXq6+9YAmvNcMmEs3iMelzNXUf/G28sVdYZrQu
5UP6H5JgEZ5ShIKBVSD4WNzqXIEYHPJ4t6cJtAu3YQc6ZYm83uwWjNL75fDxRpt85/uGgso2cq5n
NjpZThAh2wII5xvjPp+REKSFV/RpBlI2l1vsl6zaLMe3SQ2NboYG6fKds9cAwVlL97oaYovK8TcY
TSVKOOjynwZSG0/PD5dPCbcEu/5/7AsUgEQ/skCsfltyY0nPJQlBg5ltEoACD9Gp4NIJPkqKSLI1
8vPLiQ4J8V03/X3zN2ldzuwZxdhoRmbY0Fk3t22kuXn4CDyLAp+u3f9KyboYuI9hbqP+t4hr8hRX
XkXqkx/Ui5mx/b57u5PPqyMHio2irB0CY3/g0UFVcPyGQoVAklrBVo4wkyR3NaahqnSztzOexBVr
8xPEtZTOU0Rw9OV4fRrIa3vb27/UH1Kk+LJC39toEDMJf3ItV35jC38syxBL/7O2yFZa74OFK4Sg
r/nodYLJyc98BJVVQSNVfUUaFoQBNfChNWfMSXCiLcKvsWzz7kENgug8IkHXd+RSatA8AwyiTOsq
fyd5ZfzZTBJ23sPyEG1AZyNmYB5+1oSRmaZVCpKkDxL/KufGRIqjyw5WwRnUqO4xP9S6soRJlHAI
939PzBO4K1ltnEj4+4y5ey9NLivqRDbu0aioTDObD42qU6EBOtXo6cC0jozHLy2KpbdqZEEQtmSK
/YifEvqW5ZXE6kOAjA2DaJPQGGyDRS2Z03j6b/GuQ4nbEgrYxBB4qyL0NaA8FABxTYya1naEqXx7
weSB8N3swAdmqwlL7weFMN6XdNfL6CB6HoOPqYEM/ISCgeeYRXUWbGsHZzMTKF3vANjc1gYkFbqm
iM0RqxOaWRP5mxb2UByofKMZ9vzcNqJJ064xDXScio5QUD5Jgq5k7ActOXASqox3WSBinuNHmL+J
1YFqjLh0G3y9ewlJjPjkjelyk4QTxBns5/yuzC9AqJiGNt2fL/r8L0rM5iGOElL5MoMMbrIqPF2O
RQYGbfrxVhVUq1xUbXBv3AKAgKxsNDJJKPwijDAQwxvWHsNPToYodG9mHHLXsVt+SkbzGpXBtbMp
701gmVsF05c+CFiOhLzMPyimc60A5+RoC3HgvwbI+P6wIrt/lSyISQC55puGH+AsizAH7T98/DdV
VIl771KpudgTzQFVaqvxReQNV9G98Twnm/9Dml8EYrgS9cVbWnsZXuFkhHHUh3koDqqAHvZIkSrB
eflulLAz4xYieQx/1KYvzh8bMwgfnIfdmDgdVowHFpsHx5+tSDvxHfjnOtnH+mggQnvkHtb6VZXM
MA7M+Mfv5Bcolo2kCWKwnQ+GGmHfZSJ5DcSe9EPbLx/n1Jc8fe67N/SgKZUp4qULh7tdCLCD16p9
BWKxB9Yr4msEG6kfO9irwp2iwm1HHmyqzUBtogU/yjASum2E+rMO6AI7cnbJnLq7rGPiiAol0izD
mTd6cVC9HYVSgb2VzOWjwL/JD8q7aoF7qf13FHgv5zzJmb0aO/BAHbCPoDqm1BRJAFXssT/C5k9v
3dCO2u8RqkwEbM3m+pTXQyr+t9ihpGXDpUEuTDhPb3/ue4xoWUz90JlVjHK89HEYiuI0ue/yI5dh
9rhz72+62RPo8agjj+UhvOJ0t0J3LH8wBUM1DITb7Bx2aF9GZQzApjD6C6c5qos3lKcC81EdHNwf
u0uAVRy+enoXp0fConQf3Hk80aFQdroZhOirB4g0RwGKqZDATN1qLYOrN0BtqYiMPhMwSztXOw7i
uaUXUCk8BYkF3Av051J2SLCX4cvQY6pkDDustUtbbheDycwY/iPIurg7+bkNQHT9TpnRWwxIRtlF
ks1CBvxEcZJCYgIoiSlQgIZ28fo4JYfg0fWL41K5OSaho9RFjxhAupYiODQ3q/OL85bJz0VijNdm
VyTGpZig4bdmNLJ7H84E41BZx2dVKFUWyDqycJ7AfyVAsSM75hvtGgdELkoDoKoZbdLrGkD0NfYo
t3YKqsVxjYDc3Uz9gw8VuZyoIAvknSCGzrY4Q/rm/wmgiUHvh8DZbl1BgjWsWJ6bBpIFXKVY4i1s
TxVw+EldT+uxRmFnEh4l9sssct0AatT2PcvSSbFOIPEtkewwOj3TBaNLL4YJwwQxuVIFYV8LLDJz
VKHwsqx7vcuo9QoRAeRa6XMlUKbPmPOZVABUZMaFqtCcWQ02shOjOAC3Ey2GGcuFZUroDNoZ/bJa
AgRECYvNyEXrDoIsYyOcHHK8cfA7ETiEu9IKMAlxtQimCbau2Cx4VwKU7be13rGLr0/ToOFe4qbX
x/k6dUVVO07+xYfrI8G2LM2xFMC/Cl+Y5QzfbFSuIhJqJzyyayIZeu+IppCWjwued6xvQnX2twpY
Jeevzte7K2O8BN6rjfcCgp7HD7AFx/Od6ME9l2Q1z7z00h7ssCrJ9qTNODJNxkRUAbk2CdE5tr86
0NgphSJplQ3AX4Ntw0m7LdHn19mQwqbHWIJsiaXeCXYoeCo+RVtwkszduAwxbivGtC+cpB6x8WIF
oh7FJ8f3IJWKq5woQk1N3q2T2fh96hpMc0KOVWrF/zXQ2ZN9f+X3VpVM3y+2KOmqJyvmijSwIf5P
OIHIy9jcoqndE7FWyvOpB+gmSn7w23reh6p1LCO0f24llz43MZYfMjSbMD/ZcghwT3dz1LstoDt7
v2kHYxLNsyo0WlKsZVnvvIo54tXhfmJVFD1z8OL2wnd4JZFxzP+3RESjxD6PM8FF3G0sGBljj1qf
iXmfr8B2U1hRB0htRTUd66kqoDuYEPoQE4vAUC6G/ogAkIuPzWtL3QfljWA2dBXAlnAaOZvoURjZ
ES0xCzQH/nCA5qHJ0vHFNaIeoc45MTkFOWUdr/wp4EHqRFecdIPgFXowJcsAq9WUOJAXlKoGFRCP
8wqMb5m0wUibs7dUJC5Ql1ZQNSWGrH+JnalDuvxH8dP8Pitn6qC5GA5J7yAMeO1iHuRWvYapE+W8
OJmuTrtey1xW0JV8SFYB0lcovXnIv7cHt2ZkAW4BnOgegtmXqKqcv1tajUpj86wzBT1sr9trTsqG
xVT0A9rkD+GkBt4vZKHtlnwye8UtTnTqJV2Tf+4VyquwK+IPwBmc9iBF48deDbe1i5imnPdUP8aB
vQJamTVn8Bnz4VonnONnDFoHj4orHKa+EF9vuQ2uQUXN1HOsqgJvDAv/xaBc/7ULoggRnQoLAaXS
kV5w9D7LfbQF+lGY3if09F6BglCkpPUBZFMlxWZ2Wl9Yya9kH4oy6ctFGxhEknocml2yqSXNLbtG
avZwwBQiYiiYPZROXzydOhW0CXZXlFWj9wVSYX9pGSDi/Jig28HEZjwjCVNOKp1pk+G9lVYuqZbV
1D9sN5fs66rmInBsK6CKV0gVBMKh8QPUHz51XLugFYPOL778a9ec/NWaJjwb/o44By3BPvZcmSiI
CVhxW42ytlx2ZZzWCidcOwoFRi4GuETVJYsUDlRkRKjaTT+3OSgIXBxYShP7kNmIDonN1nbG7UB2
ihy63/JKlie1XjUPPw+BH8p1zZOkEaZHUn/prlwC//azaEb1BDZoEhlmq7EWHrN6z6xkBxcU12Ju
FHqo+wQ04/oCdiAyf8XXzrAnkKspJ4vNPGkSgpivJO5bInye7fWEEdo+AjM7Yjvw5xfT8P558IzS
hSZ7O9/q5QxdWsfRLDkoTj5Z/uyw0Gi2MIy3Ck062eBIRLbL8v6F4jNWDANS8CxP7zOaL3qqVJvZ
ZKfXlOTC3hHMY/t9SMNaIN1LifzvPJGCGYwUB1Y+cVqI/dyBwWyIgvsi9NEHYXkcIkwbzMfbHbDL
nOT86B0rICsc2c8eIPvDtizQscg6N2KQUcIoI4+fw0EOGInKdDYICehxbzXNGGa5Rc//LIpqxZ5l
ka/aoQTIzVQzlwFS1ibPrWWaecajmViY6tCxOBNzyG9UeLjUiLRNbovg1lhQe5QtEzeyOX4oWFfM
wvBXuYeAQWA1aPslzK70rUO2sAF/tRXoYQYulE87Z/Cv4T0W7oalQyzMmj4tPt3LLsrO16IIVVje
BhkevTvuIPl0WWK3dtnSKihjS9BaVtPD0b1kEjIZZ5kpB37FnbkuEiFz2qHARPkXspqtvK58/qyz
wZI+reNZIJGkZ1sE0Ee9RI65lY1n9lZcTA0S9PwiW5tBLSo+cBcNBorB/XpwwtvGt3/U9+hToa9f
ShQgVek6cc/X98ue3LGGoTeUzs4ZL019vlWv+TFgu39EC1PevVAcxe+wd0FxdTEt1VSsOXMeq/1g
2rBFiEJLgqHuSJI8oqlsokMigj6MoTbIuAY7LUco1b2re+K6SZ9aSOz9lE9zsfW8t6Zh3PhjTkiQ
pDBW9CdbmfdNvlzDdaV9nBsRXlQpFsTVKsGXm711wWXRo5+nlpRI4pOr6ZDESiNylnnNzdhoHJew
NRijSkKLJ1oK/5Z0oZtjrGWdLTZtscrT6+ApB9DqTdxXBwc2V0rB2J+L9ANNznBOmPNqYfDaFR4u
zC66OisNdHUq5MEde3fiKHdv6Lm75EZnRcw4kKMiCwAn89r8zkh1hvkDnaib2YxjQ/ZuUGmJUQPa
QF4FrPGZ5phHpOr19IqmmaPQuHkcpul5XbGicUi9HBM8N0wBgwlvEZ0OjLDwjvBm0n9u8mh6ZKC8
eyv+xd/OcE2YV/NYDmzp2nXurLqy2mKHfJ42KUhzxB43S0UHfH7fFDsf8KqKxksQyZtKYqZbiM1g
N4FNu6fnzGUFFpXpQqFNp+S0/bviw+0AuY+PiKVEmGLhmZRstC8524h+Ny5E9AMImzPgFyNvl0uE
Ebdx73/WtTvYifRna+qFtB1xfqiNtCxVoUhkB2loTAKYMiaTzvUvzfoIWXyYOuzohVlvRCcpY/Jh
4u4M+1vcc7b9O21tKKagzSnkjihEpxQdtzXgbWcuq9GTeJ3n4nsOPTr5hvae0pEvj/BzHdPALPEu
buVj1SGfAyNOwmgxQyRY4NWoq6dUctrnYOYJdcn0LE4piKI7zOudB/r7T2YoBrA0LgAzfiWHgnSl
LqxX/3eKdCTUX/h3ByBGImgR8QbIV25F2ITR6TzgP3JLTFdFzpe2SN2joU3kr9qHG2aZO1Qs2YAN
80RfMUMTvboFkgP5SEzMpIagAkgG0QLCBsTSfrd0I9PtUYmArfHNcygCIx+X7CWMitVsnWRMAKjP
oCfM/nG6mQtibVuWLOPXg8x+0PVPkclI4yN2Vw5FBAz2WCCTLMjaADwsVW6IrO+0V0kiPJv4e8Qb
TK6nnBjcSRvdEhBmP9cjTddtv+kG9wVEIWF0ZyizEGSOYhvTVERmnO1u7EwnhOBnTz0serqYlEuD
EYSrtC5YhWgR3es/HP+Fn3zj5a9sgqFgerdFc8OHEx+QNiZUPdvQBNWeMp86qPAqFEpq/3Znl1V0
2yA4amccCrv832acClUevapPJdWCJdze/Lbjx4uKUkwydBISNkJprqv9lZU+W8RiZXo8VS4xw5IQ
LbwtfId8ZXlUrwRjGuavaIBS5Zn2pV0YiEkejnLRvVvuYG0dxwuzSdIX8MXviT7LacGX5hMAsS2R
pxaJ3romvRtbna+/hgr9tuk3s8JTEheerWzmi+MQPRpdRk8gkdzSwj4LSsX3k+Ki16t2F+K5RXUW
Uk8syxTKeCbOrIrxxFCp3Ev0Oj++SUft2lSW2/AfV+a/SmDob1PMSF4lmORwjnQeGKz3SyO/wlsG
1SCRgQx/0Gx5VL0rQ6pQ33EUU/ca8WTwsWWcgWFFFWI80k40JNwDJmbTYs+O05Duu/+dqubqN27S
8+mWe4nO6X43qtXgARihDypTqvvOXm6f5FEHFBa5B7P+hBaDU2Fekb3Tw4K4Cueq2PBBXSI8R7+F
KhusaM171KHXHEID8KpB3AKXL7NtyK/bI2tZBW5TYN1GR/ynZ5i79tTnN9oQxJqnzMXOuj73foeD
xJcar0Dg3IbEiNltoVKvpUdN4NzoKg4w34m323Y4UOXUaUGfrL4djmFdTncf9YvgP3hNDhXj9YE5
xAqfzPIiqMB4kDNBapp39eun6lX/sbLhbUOXsyUWZgCUKuFFAFeLFXGcsK0ddjCBRfh139aenH4r
LAudbjos5y1LcgxgJdWBYRoGMRgabvpKbY3iS+gUJ8uh+0x7j7ajP4hYT8EJIYLi0XQFq+fmCujb
hg8rnL5Jy8Ny3jxfuCIRl98m2a/oocm1smprjnyoLiVh+HS85Rj8puh22S/fYRbAXc4vty5cKsUD
ba2mw4ZvyybOVJPVBTaqZvEhIxvy9pa21HadFjCMozOC6i45OV7cYBm5EnCnRjjE8zY1r4wvmlEA
NOWqBnWxsVPvxXaRUJeYNL1T13wfUEAUdyaUDQgxf8CK1F55dJu6Lo127LktTzvVnesENi+3xdpL
MGvCHpZgcTkmHv+Pa5pqfh7DX4f8oNPAPylQ/sqT55uFo1YO1PMZVtf4stjpcmpIZTh4x4yZ9+OD
pK5VE5BD1Aw73D1DWx66GfAkCfY/LsbmykfZw9mnlh6gpBfpsMI5B2lic6unI4qQpPbShk6+3GtW
ROQpJZC8d9GJf7Y76j0ejpjQC80R3aM6G+CPhocGuXryEgRq52Wvb3OulKqcISnn0XPXevXg/auv
VnDbuQ5H75GAhMJtjzKb/juO1mlROl/MgN3Wz2ZFVGKwOVCNi8vbCKlZxw+TKBfJAf6dkQcYEI9V
fgP+TeIMF4IRhRsdhlkJw48j8Mf6c9gaYKu9ky84nCBaiznjyvsTS+P9/w2QvxRN3IDyBiQAt5+Z
XTMer2qKSH9zIoRcFCnC+uVtIGko9vmWA3+F8aMQgfHkFlGKn0QK7yafRkKxRiLRZxhiucebvX6Q
BBvPDj7p/nep2hND46Qg0ADZjpD5uQL9u5I4tITRJfJe9QIVH9rj27ab8fHW6xS0I1r5L76upBK5
0bSIXcLIby9Vz2kRDP9L6bwjKDXFJe9/3hTUxyEgVLfnVjkbzTRgoOpJxLqvN6bRlORFfD3FMraG
I8YGGtFHJ8Wg33CmvssZ3MZNlo5c3mdzwySfRw6bKwZmrbqbvu8vXWnaWu2YAD2HQoka+HYL2g10
QywyXR6hSut2D+tbpdpkwa8aGSzxywhglhxTysEed80A7JhGQpMv87CDQKUahrCEoxXMkcOflguq
WKmEEupso9zvV7rw7sjMhyU6da5LGuiuENOH3jiMd3Ukc2HepTohCFO7QZ4P69GHrknruxRMXvzR
TSJoxaWQ1n6Mk+tUudU3NaQpt9anCbgnpPOEUiad1IE5t+NDYyjnTzNOHG8lg1Rldncs6PnYVEUo
SqMc88/NyHkJY2IeO6GusPK+5Q7cZxDWOUe0eBpo31qJavvfc0EESVCFCcapMkG7caZBQ4DhRZgH
CzzkIN01t5q4QXH+DkOFFdo2NtRLgMSd9AtTrXtZx2+0LTXQVKSL/rnPOEeptm9XxlVcPvNvqRMI
eKuPeIU94V94/76zoBM6543b8UXogvJifoyiAw+2TL+KiATrrO5vlJmGPVQxpROC+xh6QR/omGT9
j0UqrYbnFP+TXvy9lZkRRgoRSrY/xuUfPKCkOE78BUYML0piAOlPfavC0UgxmT7Nn1Gecgy591Et
gSxVKW6oZSjrE7x/D/+5dbfcBXQjTf6LlO0dWHmwc9xxI4IijFNbrvtGZo6gLIKECXAJTI4KktAL
IZcadGYFMC6QbCMvbTip9yCgJMrjMES/n0hDVr4aFzBNtfXFGftnJtBzcvz3CkPNyFemme6Tany5
6e9gsFcVQiXGwtocZfYgl4/d6/RZP+gTuDMeOPyQziZlV4JZPaAtEmOOQJsNdx+Eq1l2LodFuW0K
6M3qKZD294YulE3zhehwWUO6QikyLWvwREBC0Q4oEwEzM6o7o5NHltkR/2YJMTPVYFtZMJfrD0NW
M0rGaIfq83hAer6KCXwBGtSQ0OKLvWsfO89lU1jVMCw9znOKHI7nU2DzAnyZetNDoY6owHE3HEma
Yr7k1OA8VQLYb2UcKLxrtsSrpJXXFrvuGyCypDuhdT2ReAyn5jM8nuBJLBx7lOqaPzNCyJ/IFGgg
1FMV0eMvz3QiY7efoxqixWO3ZqfjlNmxzICIjzBN3W44lNdYljyebD8NcjEJC4xq4LJv5Iy9csXv
cEPKxEFLQ3TCzlOQBhurqIJdCRcBHzIHK5OQbf45XzNyB8R7CazNcfzWwoNgTwjlC7nx6B39DuL8
WvDxxsrcpSe+6Vk6YUh9NqCDVh3LdMB/iRSi5cFmDpk8FRtZS4QZ+ryxLNg3nw2jVcsz2XB4rZa3
Ie+PQS9yp8gAXDK4b0jwJBvfekoupLSx8HqStBVybHknrXD99uPH4xL0NVYqy2/vcOcGEOODvxoZ
rdGwKxkadyAK+HdN7CMAQPg9+7rkFZ4dhND7DdBWywqvo0xQkkynLQ6ciXfRveJFoGs1LACESIAe
q3Cq9l4li79bF2d6HBOeMBlQWZh/7AELXs6zozqK8kBamOINbOVrrRwgHhLuF26ayZ5cwjmU7fKy
8GdtFGITbYx1gZVcBuAnGFbbGZVtoOqA9Iu8wfZSCY07NrMY69qPpZEtC8RzlqXzjHz2vZhMbOBk
Qj6O7GdmoLld9QffM8VZF0VxJ4wFEEq1aRGzy+/yIOiYhXr2r4beR8QL5wFTpr97Lb5+NsiJRHAn
wLoD7FpVnzulzHrqt+5CMwlbSiCYYfi8r7K6AywHXtl0DNovzvZOsZt64nXT46aTNvF5m7DXZ+lw
O6I/xSi9PXuiUSdb90ghuUi/K3jxHA5MeRJL4a3Hn5PbUVtGakei0THvFuxkBLiEQqQ+Oj8Ei1s/
/7YKL18t4AK5QHlex9XSvEwHblG1+70SnHr8Ll+p3plz8TbrPmVplBCdK6LlTo5To+7eTqaePmWx
xcOOSIKjMWn6VhYWGed8J5u8DPRLdkQvZerc06mK6XsHKlojIVZzbO5n1fJ9vnOX5Xo5tSeiPQ3M
nm1shP8qWqVXfkx+421XjIVVMgXSRje744WO/Uk8bMSjPZbdLkNBMC/Bo75NCAELPDEAHPwaOHKO
qmDC+hV0KLfpQ5G7PV11E/E0t7GBLQJeRTTfjFyO/MWvw/1nlNVywUCZuYtvn/Fa0WMsfACQDXRT
pmmL8XY53dWsIcjP5MYAku2OLKkBcutAUbiN09q77XexcC2k7gpYm20QO1KSytCpcovZJ77ayL1F
rxxEyvkeyWQ0eC+PWbhqF2lThKQhb7MXgm2KAv8AHja38R+Xm/UFKFmRPtqoaQ5EiVcW5TF/OnB2
fLJ74M3wOPJK5tWlTevAWHQ2V/uL+fcCGM4Lw4iTY5zLL6Isx/3rnZoU4tpczEkreiD6pCNr0li+
QUSyErsTymlpbr6we1ljdvd/QYjZW54QTOHEYceskMkYCTWgIDgL2AV7qP9kck5+UszQW3n5MVoD
oaFMkKhf5aPx3zArx15zwKr2qklsfhD+RqrntlofGcrrNCxZxCIg2vTvAGAdSI+l5cWyEtWSExeX
GOuFQZ1XFcOYCFKixx5muFJz+E4CpfdrOZRuE/b0Dy4la8u7Dkim+xK1RSj8vMwupa965pjvx0Pl
sS9ZcKPS83ISG0CqSP/7w28m2g/M0fSOtdUrkgOyuo9U/rdAV7ztdCAgU3JIhrtP7u/+2XyeXjWZ
RHb7PS26LrvhQmJOx44o3II02iMMEr9wTwVAy9FlPvjguOz5Rszzz/jzaJ8XXaAIYEMqoETb2s0L
YAGKYi+qul3xxi72LjRluzYUCWUR9eRjBlv7DRHOA7A+UeOfGK9oq7ploM+tVHGZK3oF3JLKcgqm
BNWPOcVPdVu2hiMirtQJeH3NzJ9gWhz0snF4HT2DreA6zVSi+3ykH3w/UorOF9U+8Y7J3fClkJ3K
A/ORH5+gQhPd9ZPgzQxpqP6F6Zt93UkEGqLjcUtos4xa0Pjl1RRbvjDKD5laTbzcBqDCAiXHRTtZ
8FIauuN7Taqhxeye+KcAGRfkmRYPl1XUA+fpovgUkprM7akoT4dOrs1rkErlaigZv5oV41NXbAYt
QQNwBjFLxOgx0NX8qKQYTTvMtpNvUCyEuyg/I8CqXL1S+ixry+oNfLlze8Or9fjCS2FjUZvv/hEd
R3Pe8/SJcwlg66jEugHhTR99gH1GL4p8PA/YnTCxdI1iYCbN0j52DBbewbnqLga/yKXtXBmDCBqn
bhYT0wuUiQnzAWkxCTb86+7E0rdjigVEttsNhqbCb1of/5iGFqqbMqHvEJ/qUbL8De3DQSaqyRuX
gzEXc1wVK6a4KxPlQVADWHi3avWf+lyJ2fkMP0sDPkkAeyAAlwFlrOTaPmMW+Ch0aav/k2Q+MtkO
UgZhE8xAA2pZOEJ49rXpVpJhDIlgA2u3I1lCGuhsLAyUD7xYvV6wXellviMPr/saAiklkmq+fpvn
HWMmenntp1HZZqmbOEaeSRGsl5TWQ9b/ECXKfoMAY5t9z2LAqkotEKn4X5pMiDbR8Z+xo1gWANis
Ap1IHw4oFM0jIgYXM+cZyPz5PR558Kf2NydpVT+ThY1bcQbWa5kysdQRYe/CiDZlAdD6Jl7tH5P0
Uh1AZb9lA9Msn+QNo7T2eMZHQlvstkHDFAHLbDzfajS6NwYCjSX+u1M7m4fN7YvJBLMpAUMO1fnz
rmc4o/ADULL55DdT9IDtZ6xBQh44Mu8sbxAfsj6+Ry3qxZttJNbbMJSphp1wNxj9c4NLfWcQVwEN
xdyC1uoa5OpwuNPLnOSJzGAQRcAePB7OhUxrZ0Dne+toYKnPQAunqto1uVm57cFQmrvHWO44+ve3
hjht9zm85iu3yDOl0vFvoIf/uXNgkf1pcCHqGBrWzj0rZKqAL6y34sHo228F4j+t5fU82/XJygiB
iEgBOm+Ph3FYAlqaBzKM8qXO5nPflTICdj960lILZvGiggNGPEA4aESNwUmNWde7cmDZonKBtUMH
pMXJgeMYhQ2aP34hipyDDsdcxLsHE1ciLVuXHzrlUGGsiVtlZHStlG2yXXaW356MGf8F2g0Yq0EY
8US470MdKKJKoBoJLFUAP7vTP/i63nNKJzcOUGv0Kl2UbaeS5s3eXGETEvIFG3q4U1GwKl1QjvvW
yWlkcTe5p8dXtGt8n5iAWq8LSjEbxRUULJSnc7nKW5Zj4+mqp+MVl1KDbW6MSKuKHluBcSVm+10S
AZrjMQ/vi3zSS1FGk/PpAt8PV1B5A5qku7RDnif5PCs+n2/J2EJaedLFAJ8mCPyN+Nc9iKo59NAk
2fSdj4yWtvgpB3dqy2oJNi9rqysH1ysIbjSDU0VluUGXaZ6XfBJgJV6PDWzeVEJ3e/dEMDAf0PeQ
iZP/T2aLE51UBuYs1DyN8U3jj+HfcoRjUZLyPCWWOZnyBSEooatIq6h2OEIJq/KPBDHQaYWFMuzL
k80GYO7paBn9fdZeP7zg6PHyTmWvR3bz6VfxsJAFzuy7o5jh5sXpwUjoYn/RcBgrdWlrzsv2VhyK
RQYJCojbW/3pBBlj0P1265wUyUDH+a7GeZXQ82/b+rhPILVFGcubQ9h2VAZjaSkQ8xPzvDkBRRkZ
Z2/2bMk/NHXrhTcRFMqTvoaYJXl4aSfsWzou4/nX6tkBjvvQwFO97P5t0N3cxeo/NiNqMAXgIN6R
Yog2fiybAZWczT9ehVe4t+UEjqTWvXs+VzlsIy4Hz1A4ozm1WQ7Ci1IejR5bATJjrFypeaSDV5C3
E2BfNkjInrVouQqD8/CxrggjFWssMHkeD9zqRGSzdHpf29yJH4haXdpKjg3MsGklxRojiXMwsjKj
RnM+bAnBUtlvmXVGXYGyezL1TBij3eq6J+Osnj4H8jD8Vy8T7cbqSEy3t71+huCNpqrbQlQsaVky
Ptmj/LnWdu3tcb/qa131L9nNZnahhOq6LJcbjr0sWX/rpvakza/VZS3YdRJ+I2Fzn4PcK1eepN7h
i/7L3mylIX7rNmpS3C27Jek3V3av040E47uflEqyS5wEMh49ZLC7ZD6N/Z+emfRdOCgXCzOaH9b5
v9ouQ2xdNCBzSosi+zqEDMfBNJOSW6KNVwFgHao3K5EhnWx50UDerT7pRuZTURqbCtwb3IlP93Ji
92ETkcihk43OIC7OT9lPbG+sco+o0QtOkGDrxQI1+7WP0q0qAYCGyfxKuZjp0UAbUiKh6LxU9dq/
ryJZZq11r6KelhRtMgW8j2iIP8tdwEGFKZIzuiy92axxxBwXJR0XBk48evY/mT0t6kBjdH1+t0BA
F9wV7r9Xdghox6xtU1Bzjh1qS8TrZJ0rT9b5nwin5l4/YL7BUyRzxtlY46RkkEeJv1kTQAKbiD3O
YlhU+sIBu3O4orcO+1Ws0zmrXr0l0oMCduPyOrdDz2MVFWu53e3bWlrVgzXZgDQWk5JQ0Gr2qy7V
6gkQ/x7FKCq1xaIAipbLdJbXNjCS3CfbK0C7BkAjzJQgNPaxlm74QR9oWxiPjq/ZMmcMEPAiwPgc
u/8sgIr/Z1LPGblVdNYUWb+RcSgU14CLQdA8YrCYMSiKeC56HNa21WClLBsdoufLzijhVCYXQ5hO
SEUo1vGK3XDrnC7Y6HHKbXvlPQzg1cY9RhSXg/OR9OXd0HwPHBMYzi/ipOzzpifWqSYaNqvgtPr1
hx28VLZBrmt5caUcLlO6o+oXgmYKruOxG0lfb7fUnicmQ/7j62YGbiNi7HmTSo1OEr0WFLn6N3Y6
Om06mR6NIODtF9eM9TnENGXea79+3XNIgYT4nVIwNIa33JqNfyRZc0CWpMhrjkrEI+qg6IDlyZIz
jIMb5fItJiwLdE9cPwUCCxR12zrXTRPuJAw6v4GZiPi19QBhhFcLI/xUxgtBpXNHHzDZIhPIY2Jt
4/WqVc6hJwfayditVD2Y9sxIRgiOOjEL3/2JBPlNGVSEXwGHnNHrTZSc3pjSh8ZwVx9GnqxOcP7d
q5WT17yPcPCIu1yF9Hej9IuAjjlqNUpcW4cqAWH/JRTTBZpLLZj3kk3b0ITM2Cr93nZ0TdpWK/Ej
QR6fWEbCiQFAwcWxKp+CTQsYQSypo9/6n9StE6IuSLZYFnsaKkbXK/bXibqVBO3dtixt1izRgQFn
vtk2gvutTMJhKcS5tPmACHLTQegou3s/U9TQtWodHqBn1/mWpUSvFj7Yx2bWm4/QQyKVB3obmfR6
MqwEkASTFgJyfEUSkBx+aJUezq8RQFEO0vrFYE2wkAc7pgFwPtMr1G/l6sfx1QW7PNKANH6FvkeQ
ttdifzaNXr5UG00rKbIBcninIrAPJRRQUAS1uBYUgfrdalbVpGjvgxfsFtPMpsxc98UAnTwIYc9e
iaEpy/Qs2IbVzcT0gxxns2js5PFvcn5oPjSuUyBOGwdjU3m++3B3apnhUqTuE1b+Kracn3ZY7zmx
hlDm8KQDSxDeNdVTWP33aFwWht5lsYysXzJnjMhiZ302LypGa3UM9HCDTu5N3KO4bHMfnnmZyzfU
bUNxAeZ4kdbaXUnZXgFxPmuuDD0SKPZ4Y7iHH1Nm1xFRlJ8BzeiLhX9EM9LUjih80M008oJbj5xY
NfFnT+aoHQrUofxPk5XXnbVjsI/+x8N8ADeNTqiYUeextOgwUvNCqXF3u3OXCdmNvK+QuHJLmAgp
/pp8hJLx9hIMr1Fur+o+zxrl4gqp3NQovUzDxezWB3Z4gfsxXO1cSVeT9PaiywyS28OtCckaajQm
j+OB6FYA09OdMxbHsI4YWAsycHFQ4xsd08kxrSkyOWtsUI2bDOp501dgZP3DUCjy1oQhnL0dfAQl
5l8vVVQopkG0JnoDRpQhfzq9KBqrXltNpqwEVqAxKJgR/cJOkqW/7z4Ni3/r6lZSQEPIXmCFk4hg
ZROaZZt25vqaaFeGvq4r7tPqv+7csC5Hly5x6bp4UBIDRExxlXzGAnmXVZchMdmxU1ntHc+jUIht
SXC5LrMSfAavqjM0AOmT8O8IaTY6VBwpqqb7ztilQw0t1JEu7CVVjbSiZrk44zsd5TQhztDKvv5X
Dltmo8A5FQ6Sh01RuIepEACVEU4EZEif0eXBlXXpisfgVyG/eaV4vdX85+744rYxqYwkFyFKM9Ki
7jj1/8ju8XGgehY7N3o6XBF50gM8grB1v/jtSoco60466Kg3ETV6pcauzsqzsxFebG5OJZ3SAFX7
k5TuKNIFWZjdIteNVV799mx7ZhNYEP6CFXJj8P+IH+nM/AaB7Pxt0YhMiGsunztWzgAZhCR/bfLO
5qxU6gdFqF9gNMF3e5A+jEF6EzVv3sFBK0xAlhsJoracnP++XkoKSTTXs1+U43oCODZH/en0Kztu
IRZjTt3jc7+zeoenxwAtyxuKP9k9aw96o6EWHAtkk2cJLJ9VimVjr+9D2pk7EAcNJ1H8RXstlvm+
LAxHrca1QhPN0QoLROcKQX5iiMzcEbCdPNoJnB3+uvRfru7MZcF8GEBPi+nsktQE5SEhHyvqwQ0U
68JhzGR8jg9vATZ5k6dRzx+6VIQA046ZRut/WLVvHwo4TrIQuOMAlS9h251/zEZ2JzSAMt78AfAM
+IKdD+sT6QHUweJuExnfz7c6jLS5skekJkQPNFvc8IPk3NX2g04ksp1OZl0eiPKmHr7MpNrimci1
CpdAywyVwE6HPrFdLNNfWOVrJESdWj+5wVX1CZsaTmSbjKLj5Ivlkq1XmAol9QkVbVeY4fnqtXWh
5kpDzNr7dWVGdmI704nCoX5jzpwkpTZEhjC6rCApMWSa8q8sFJdKCOlXCgYfg/L7pZs5ilnKLtrs
EzIbBTjK6i8BT4X6AOGwzyGw/m3xsjHlOEchFixxfTxAuQd6PYgeBRkrPGyHnwwWqjKRborzq8Pq
9Ajcxjmp6ctoRdLLx7FO1NkbqlXqWdLgLpjpvK7JO0QIHe8cIx6rqT6nvmfT4ZpPFdTS8TfFdzZp
r3kYoEVMS206QEBTVoe86j3oj8kWx0tL6vY/mpA1TFSj0yvSz/oEezdKfgdLXHAIfhe6o9QPOcAf
4C0ldcdV7HD4suhIiUXjV6Eu0JmLeOeugp3mu4P2s58wiCLOYBJxuUcnFB1EGpdVxWY/pNNaO+Rg
vLaaDFgi5Yg2ctmNgkeCENffmRLgQ7xP2I0Hps88oOdQ0F/RCCSR2Lhhw5UNM1AdIJJpymFNP05K
ALq0LnRyKAKu/rVfwfSoOZQc7ug2orfdOX6DMxGOoGCp2/umhZfLj2MonFxgchMahF2rlRH2YGTx
Nxx2b9luE7DESX/pxRz6idouH7FSeC7U6ztVJgWtMA5U0Co7x3/D7v6FsYhaGZGdYZVhoH9ybUXg
zi4YIT//sTR0/Z/qO3l5g21zKxGFsgAPydBk7dvGhgRu+jEJ3yyX0tlCyT+m1+oq3JTqNlgf+EXS
ApRQLCTKRCbiHk7E+At7b656rEbRS3OCGxKyoDnPTLUCeiEzn9Tn6eIOYU4uYQoGwqMpBRULkhek
txZAoA32gB+lYeq7b57NL/szHZAVHLmWInAiWpfnhKKZC7ExL6xAH0hm1yFOz8fZEJyxLnIow+bF
kztvwgF/UdbhcsFAHb5E/kEWMbMwCM8B2t+rGvW+PZBT2kk99d/PRMnlPGqC4Sh4l3wMFO5FGLSL
4GtE2Ob9g0n3vTO5PTNIFYKP6Gb9frwviEiwlQ18cct5QMcWjIG8y6xgPa+vtc8PilhXe0ueLwOQ
JU08Jm7iTcD0S6/vYocdJR+oxkH1EnxLQtRbMV3cl2vqHn1z77hLbkkM3nwtzHDU0nPDkADtjYWW
JTzSJ34kDANkZM2N/WBZ1btOSoB4b/gvIODFQeExxTZZnrXKAW6Ljwf/fdOoY/wG15BlDhwq5nFW
EHH4FIUhQvI5grs8+7C9gPF26NlxWqwNkiyc8HxcNJYRT0yy8SOO9grSOSXp2LVuNnSmAs6L8oix
CNIKmV/CZkW7L2MEbCKAG7q3u/UwAR11fnmp7a0SE+JohEHcTxwh9d9US27LNa00mSuZOVkVz2bL
BFpUbv/zJiaONTSQMIqfFBdqWsPi801MJGWzZw+8d20hF8H7HVuv4DFoygI5+aEJj/ZdH7tYuqWG
cwGuobs56pBedfyo5b4k9SHjFYOzYLMfLI2E7uyVXra2IUNCF/j2XDZju/idNG5Nnc0lLGzvW6P+
L+MJp2iGXPVbOzPHCRisamYZDWpf5XeUxg0gscbboXyK7sN90/zbSnUJ5LCAQzgNoQ5aVVKz6L+j
oiO1mzQCKv00HfYgXmFLfD7eZmTFUIg7mu9qO3sejDJ49H1s/XDV2KLlN0uF8HBb+3KTA141bhcA
uoSBeTkE+CuVwPwjbnWwCLywcowjQmiKOHPCbtEbNrP8YzFhZBVtCmniCqtVm68IgFYLpTBtb2dK
qwRNiXxtCpKe1Pxjm+3YPFLcmIA28DVhRSs0omyd31JMwUbKu0GVt6CjOt18bcIyP9auOwxI7ujN
Sj5Nwf4uWYfECyOSnGg5YKVqApI3S7dxsRTf4Qc2+t93drMOEdyvsnCur3c3i8X7w7igBdYT6X6H
XvfCD/K/JvE7rg4Wv5Oo4GeQ93lKKIOjGWCqaMzaL3eJpXpArGa3vEZiMcysEVs0tXJjfQxTuvca
liMKtq61oHGG/49jx4zlP5Hnswq/vtdkeN6fgaREtAzKelZ1lhSXmUznCLap4dy8y3H/BB+0duZd
Pkz6krQtaUpxe6faZkAFzV3dFyv1sXU67CFwXRFD4I7mAWBF14uuOrZUjS9aCwNHw9GRM5IIO9XB
paiSPzpYgbxQvFifuogqSiEpb5AphvCBqMsDuCzQMNGssQNt88bNfBL3UKbJYfQ+S8G+tWpr6pxB
KW9SERqX3/dsTxp5YatpU78MsgCinEU6/JEdjjL0j3zDyFRlGIqsa322IGwsCA6tBAE3NsUeFGPf
rE/RFqFA2RDoRbO+4Fo4881K0qLy2dw32AMjmPadN4yPflGa3y+J37Db7/fXPXCvK2Ho55HVp8h+
4xW/WyxUVYSSdcRc5O5VUBxtNi/iIti1xeR6FWs5rmB4kPx5U13Y6FL15HqHyOvOxESs4CBHidA6
QJbc8+q1roGPJMXFaoQPUicwtqIpp9Hp9JhpLCYdgb2y+QJfWSxuj/L/PIHBPz/6Nghw5o/x5mLg
YJLc1tvMkuWr8lCIPDoHdZP+mkl4O7MHvhF1ckPeTwa3U+ZOLABKSgSLslSisaAnxGLPnMkX7rsW
rBRY7lQMEb0UmLc/SjGp7ed4MazPiNPsO/r9FzgwGUDJPKY8rsiz2oBAysQHXvR9pnhY2olCgK2S
T/88/n4oRqJPmm8Puv10PK9UDn/x3AzWsvwWJtbZETihpcnRfbltjqNaO4x7u2AYMzhQTFlP8wV6
T/wO8iLwg0aYtU2214/o/4a60K2kcu8w1rWh0CKjUUBIG/nXELW1PdqqmhuEoXtE6stPM3uCJf/7
aXHumQW0TJt3YKsPMKNxylD9fdTBM+7ih3ohEJ8MMrGvN1myohVkob7hoQCYR5iSf5D7VTx+Tyex
s9bJzr3JJ9D/q6knV374XQsmrwcJQbroOdeBsDN6Ouv1stl4Yz1CcsjBaXOR/W8EId+U51tVz5OP
2xqPPrWkHk+ecYyLkS5pR9bkSD6v0RqOlX4Xq14jrd7zvr1BJdm4cvI2EdCWkU5XX77gpqP3MIO+
4OIblMCpm4ovu/zKn4XEn46ben9jDraQCXjgznFgG5/oVtEqXg3PtbOsEzMk0pY6k+MiPMP1grvz
KuzGd+VpSahxzQ6g9+h6n/unF0MaEf3CWxJysIxGsB+n7kpa7rZXS0KU7w/o+vcjDdnbnPlkLvyG
zClj2r6LIOqWDqojYAG8sNgm/tMnYno2CwQZzSKliMNQN+2LHskFXXN+fyQ/navOwSjUNwumBSgw
YavK0AwJ2eEKTQ73XjMvfdiO5IEf0YUHDtIrRLUub3xfNHLd5fyBTKOZ+Ee68ueHMJTWZ5fGtcRs
jIHMyVN6qdWwS/FiTWWLbZnbeqxJWexLXyH9AxfHNK4T5jeHp0Sn+hci3wn2RUpGJVAPF+9za3Jx
vXhWSa8Xa9T2jQEztjVtV2txkzkc6499Qgg+kogbezAWPee/Z5dj/+j1yAfBBqojRINQJy/7u0qA
KRgZCrxw7UEC82N3GcAQdmQMnaQ+I7icEnhdeVGwtj33EncRZWKvzaqWuLO4XYvDJmsYei6IwlrY
lAiMGumFCJMioTyP5cNHXD9JaPefIZRRvYRG2mccUkGqgpOAb9TFzspLH1MQKMgPJ6H5mPPF7kyJ
ANjGjAXbnt962ZilsMbZAQcfKqVbTncW3hPOEp/r/ZwNxKZHe22A96UTEbglltsXqke7b9Ukg7DL
276JrNewDHd5vzEfLk8njcfv1ttF726fla0KR0pxN9k0Vm1DtFUOAPndnLT1miTqWjFjQIVrb3pv
+1U5zMVS9uiHbK1PgXP/dTY4JcplyJX/MrVLBxnTR6JCHZ2E6psTqChs4RJHhN2d3SQa+16q9wzf
NQd0Zt2ImZSW+bR8WGhxQ3Pj9P5cihTIOxkwYrMD9YWbuJ0JdZ/tTkyJvu6obC8m+hG1WlU4CRvE
iSX9hKKFu2XZyZ0M0QeSV8uhpKN+Ay/1WcZbIvJRHvzX/OjtuyD5mXGuCqRFDZAgtUzrHiSWB9Mw
YUoFcZB2+yPRUGt1O+Qyd2hEJLJhJUvaAijmfeu+yxaULz5Z50W07rg/WIgvemnA0sAOYv44X3/b
ZQYoQ70lnTee24JC7bFAsdlhE29C1AK4KJvbuBtz8ZdclL+rSqdLwbpjhOlq5jI8cLmYRtZ+u5vV
3gWoP4HPexRj9vByjKWCxGAXuTlvJ3Hmf0jqDYJjCEGnFixKqZtHdSiMVAYknTajILaxUGYnofox
ERQPpBIChjMn8dRg9DlMUSs5cWJvq0ONjOjtNHwhk4K6u++qi4/ctgT1g9k+jUFAm+FuWfF1+j2S
PBRlaGN45d2T0TjFzvE4belJiHvaOTuQ17U5MlLh5JVev7JIkUsyfhSYcT3F6M/14oFefE6V2HLw
q4JVbYpJrDpu6yEQ9eItsyxLwpvOKYNk105MU8iM/OtOqmEWgXmZJFfDpYbQqSJQga22zPuSqdXB
hsl9adYmS5h2DLZ9pqFLpJscyzJIS2ncXToBrwj7JYazjflhHULkzkEd1IIdE6i51kh4PN2VxmkE
Pwj/WTcycsn8O3kfUJqU0Ft1wCUmFFTFTaPAEqmnRkdCkdlaA252T0jIMUDk2XDVWT2JKp7DTHIS
rYaUn435mkh+FUZnZPs+8AvKYsAfHW+ddeeJfEWpwIY8X8VUplcUTN1cNauZmA3lai4tjiG+/Rd4
pw71NhiDPW9NBalXhkLizK9yOBn0WFGYbQt7jI84a0jGEN72VoHQdy/w3x3OL8ZITJf+h0aEapwl
qp4teWnMVxjYm7qG2bcL+DqeFv4/KFKAhIxKV/xZMdvT5fQYXDq2Xc3gfps06get6USNq0mXtXpW
HTEWm1dtWs4CReDoB24bw7pUhGdd6EHCYoeYhiAP1Hlf1wdz/MPAbHf131Kirqi6kVDpNL8hAHOb
FG/tLqpaxXu1yetYyO7BcM88DUq36o6Z7qAzkw33GSKdpnC7g/t3ZEUOLvb8geneJt6AhHA+KTO5
PVvL9JPAOdSSY0EUGDMe5rdPde+llvf/skyAluW52QGmJpayRwdjl5tJQFWci7UMvG8C3IwA7y4a
awUjbUuC4YktrgdFR5ggX5qO7dmJqNQI24sRRIIRH+HWAuy27x9E7zOVa7leJNwDkdfMdf3udUS7
JseVPPuTMOra3x96mRlErSc1Vs0jT10bG10rtBY68pXo7a76G4irhRkBHUn9rqVZnmHnLBTm2Mh+
OoJSaCirZRhhHt5RD6MGN985rdhOfqXR887R9IQfDMMF8id9S+MeUf1pMKq6Hw/nv8+w5E7j7CQX
0+TeOmsf/tcW8JENcIEwi6xVffRV/5ehYbdNYOOFoWdiJ4UueQ4AC88qZXAI8eA7yLOKEsH43Uye
tAlmLn3b/ypv5f8BqKKijxiLVpVy1Cz49g2BaaCJx2NVFN4kisCQWu2klIP8j0gb0WrnSuGhinv4
gsp3X9eIq/ZTgvGuXG7Vgux31tUZGF598MWSXt+drNY8BrOMp67O6Bq5i6EHnLetWWXTAnNWR2W3
1I6xvh6AHBgyrLHZFhZyAVYiAB5BpIqH2dWihsLPYSvK6x00eur7EK9E/Ytpw2DHgjLM60E9qDNJ
SE/LK2TICpbO2qqyeO1tTXOVdO1kf9jAcmy4i4gLytZ/us7NGdOPXocs1xwQQ/yNnWqcDOFq3p+S
iMjmKfoQQCDF/92mM8frknCDNNhdbN0w3A7ICAh2Do9lzMdQ840wnow1J5ToWZsqpnDuqLi9Xhs5
zs/yQMlbTEh9KlBUOyWDQNZw52tCjXRRCq8bbYZcLwgSfQW21FQNzwtml4iZS+j9DlEPOCkKeepo
AVNmT+CuQRJ8BAM3GbqLbJ8cmbHEE47nXIueMF+5MzT7/4JxwzqELI1K1h5843x86KsqbajcP3qo
VHOXWqgVrE/TWUHUW/IRaImHCcd7ckI+XiOPHqj5BTdZL5a29dd97xfM4TogTLbbFMVPObAg0HAa
U9MM1mXVkB3WOpSfpQ9Eyrnuwwy98hKCVfr9x9sJiZWItyi5XCRqcOkryTLHaqHjED2+AzNpLWRT
u4tPcMCe0sANhNgwrEGZVLIfhXMZgaGr683WBma0CEOPrkCTo/Ia5aeLdbzxlYvxraWbkj3XR4Pj
/TNaiFZxfM3neHSfdVWPf5HxGFjePPKd2ycboR4HLCa1nM0qZX5h2UQVgk7+Q5bBlvmAfDc6pMX8
WMDk7JzRcME2hSM7DamZsmMGMH29Hxiuos3jwMMCCJFG0ZfSd3H/PqyYoGZEoF83jyYDr0pTL1Pz
jSLmTq3ROUyopLg61XmbcgFUlU4zpHVBwWy82Q/yZPCCJF9Sb3Jw49mrK6/6kobiP0lkwg3D/p2n
mc4Tvx+wwQ7vE+ofs2MHoLmVcXhrK8DUFP6vnNgsP/ULfOvCMAqOYj3G41JCdaZjygbRa6xRmMGS
IsxP1oVzqxaJvNQiaGRXHxwfMmdfZ4dStBiKLAt8J66XZFnyST4hXWMyR4gmVj/G2EEk21XbIZ+K
NbSqVV8GcnCHl2eZDm4sB4ZL3mfTT9pWzZv0Orq0+EUTuLKOd4EnMpKP796CA5n7cxfdBrYkEBC/
luFhGN9JzmFRX+9x1ZcdtWGYMlhK4ifE2QCl3EplOirf2q3B8Xosz9UcI+gmVVCgQjm+e1zQ1lxB
sIoAQ0HnbcSn5iR4mwu8/AjgXOM/Z9K3PiserFdBmnuPuQ45aei6HqhFnT5P6fEIfJnsJ67cP+lM
X4Els16VDVuisGKZLx9fibKnKXQIT4HGQ6cPbV5Q0JS/yb7aQOC8Jx+79dtoWdnwne2FZOjdOES+
4JwrYVqi911FPIo6izxLq6xxPvLIkoZLFQAQjgT/ESzii7VtJBYJ62q6rCrGdhLOtLJ91qV2K1vK
ZM4ScjaU+2//sa6wu8QTOG2CaGv1QGk2sjBjdXQywks7QzjiMECYT558q8P5sctLx+xMWxytgUvS
slsO7s0Rnfwyuc4MfTvReGzApr4MHJE5KAS8tj0nfM7mperepO/hQxXpDB/llBt1zmSZhxVLtFA/
sgfwledGumLXnbUo9VH3WXpynCCnjWYbsHbeX8dXeLR3GQG28iTNm2Ca1uKGT5ZlpiTFOh6vFnRt
+blQ7YS3BR3KceuWeYgipQtmGc7upLBcwvlQgXBhwmTAnO4uHPIGCxuLMPOV8G6qUu1wo64K6gpU
Fib164ls3udwHAUQo2dm/c+qcy/2ocVk1+UmKLWhVApImLR8VWAsV5TO9j7leIDdCTEWod9SqQ45
wTd+5eDiazqgLzUSaSIR7O0NNzy3BN0s6+rmqzmTys9V/+MreiZeEgrNh5jEWOqQyUwFQv9Tf088
zmzSud25OjT+mCBWyYAQJo/wOOHHGaSFoXI2ZK8ULcwJ75TXmpdHsVGNjuzmdyElySY0je7W5F9r
Pr+1hMeOqIVjGUlJjxAsatWZEgiNidpxlnVmRVr3xl3IeQ81WtI0TAjaOGfJYkHt7JFIAhMMWtq/
+9OiZYoeAR5cBZUXSBtnijk82kcTp+bo4v4hSW5rGWGiI7dmkbC8Vmpih7f79XPIM3sW/oX0Cayt
rsRxOMDp4zophoH/sogo5Yp7V34K0lCUHYgWc18ad1L9aT8k1Ej7/wM7TBno0AUT8Am8t9cN5NTs
2D3MaF79kntlNJnSPXEbg8yy7oYJdZPg6bH9YSlxyZ/2Naa73emkEgwpd1uySIu4sg62MJhi4+wT
DGCpRL6Ez/IAI73Ff9h/jK4Dxr85jNzOTUsfew4jQ/aUGetofHU4xsNhYaym1IsXzv302Vwsg6kw
gydH2z6ehONyoFTtgBzkS8oO+nM5GWvTkhKacwu4CeKPbg1c8W/W8D0Y5TSHUoVv3mFYYEG3rFc9
jxT2A3dF5wZ1uSvMoZnX+r6sQLrgYyyfNL5K29LuYQs/BeS+P/YOglAlwSICMI9PBUtNCTdJPMJR
DGJ7b1JgeRxCHFO8wrRLjBhopQXo2fCYu5Nts2nL0uoXnT0ILhd+WH0Xh78CmDf2axfKBgoyk+ND
m38R4icyZgeRvLdCpqSGjIJORGcCPsCIDOpOhaKW8byHoWsx41Uc+jN8ZZofgTptYI5kc+3vmTeI
xZGHLnWgPyB7s4+qss4pTTtmLOOnuV08nfbLmsbadlwljozHayTWtHo7x6gyI0H8avLDbWrJMYfv
7TOGtpbTbDDmC/kayV7tS5qgT4Jjvj8DQevBJdxeMIuc1PVMbKtheblJa2IAutMjV80ryiYGX5z+
mm0sjHGldRNqnbVL1ZgejPpDboqiZNSSf1hXbkz62aHskghKVhfBVGIMxTE7L42dXL+m+U/wjvLe
MmXegrGNuxv4r1D3FkLN2EkESoRa50qg3v33T5zMw/rw4Jd0EBi0sZ6cuemsIgOuD7SGuYRmUCYv
Po/jr1k+CMr3wOafRqA9azFWTVYOaarnIHFHE2e0Wnn+3MaYVU9isbbyydO5NVgc8d6mMxp1Wrj/
AOWulOOxOlZMb2qQxPlbIPKf76Pj96XfdjMqo4ejBdrI7dPoKzgjFyQMYhQ5m1stkH6JXMk0o7b/
7+n7rkwIsk7bpnh6jaS8T7peI7PF60oqrPrBdCleuzz9wq8aw0ZaUNGwNdkfZkJj40gdqzfjEDMT
URO+b2XS17aU9COWnDeXTTORUEsosdRUz22WI/Z3ISFqwh5BToouPdynChh1M2+N/Jmq4rHrDy3I
RzvR/lY3sV9sbqnZ3Ee3W60nI+sw1i57jQCm/0q2p0UlPJI7E35DxTisoEA0OUMkLp7WyDqSd1dE
b1o0hOgSooHAZAdHJeHsBlOB0FDyfg5Wr7yNceAZ9ApYPLwt9fzXLnrO441Ydk299wXn7MRiBP9H
EuQMHYZpCP/YNY229dVucfoN1gA5XxlgcJ+1s38sXKNvoGckof3ryYpUbigJ0vod/bbrFxkoBQpF
c1tddK1AQWfEC1gp/ftKfhfU2HlRUB+Dkl3e8Hkfb7m+RVd375xe0oxQFJUH/VyGY5P0sLyYUBPD
fCyBjJVk1f6ZScNzgGcmKx+82cKaa+38kWQTTUTIy+bgTSlJi5KV9jWeKWUzTY4vFMI4ok37w0Wz
zf3psD2PkoHtBX7cUT3BYMjWyI5t7A5/BHd/x82WgozWKdLiYa9V/iWsNA7O9Z90RtRyUvY5WM4t
zxAMxmhmAIi55/ZCOYP7NEaMYpoUGz0Uv5By8bKtHvhI1dYWX2+oavLcF2WCmyOx1lQb/T8dpU0l
48RX14RP4t6aXQRApfvRoAIFLWFS1H8zjsvhLh1fMBQ7NlCdl1PaP066WnKxIfI7mGzM6hGBsFMU
yhh5opU2HFAaEXTwHd/z4DbXWrY6Xi9C1MbX4nbz03snVHwKLzi8nR9Sqt+BbW+RRQ4179qY4yU6
rNJTcIa9bKTejJRqZvJud00VlxBDLuENcLVN52i1tCMRHCldy+mQsicxygyV3DjuCUN8ZeopY1pu
AdSqWH/SiW3gAeDHxUy1mri95uFXJN7otCV9klvkJB8MKZujY37+lp6qAJ1/2+Ab9uPWhWhWgWRd
AtNNvVo77G98cQGFTK7hOtoJv2MAayPSBQuAX3UVwdbjhI7KjLzNVGUdQ5CM2q4dysyoTILc+zmm
EXFH0dKM0rrLVphREVBuWII6CZDyBEy4FZn8ef1mgLKNRaPa82xa7qoatEAdWkme7TNMNxTQsgaD
+Suovy9RxRLtUSK9N60llqB9+j3z+4aJ1w79N/cL+apQu1/fbLqiq6hOBBF4zytG58nD6FF/qorK
YWjPuXBjjk8N4XOlQ4utxypkomcBjiOiCA4wVjVevi0pHd4oTOD6SpNWPL7aQp07Y+mm3l/uGPcP
8igSQPme7/lR7vCWaEj9f4b5uzWGWkJils0dR+c4Ed5PiA4ZJiv6gGjIee3dKPeXRrSYpzBECEdX
uHNYdPEiUnHQ48qB2/x0Plf2F+ivMb0apnq17om//HgJO4r5QgzZrJLL8D5hEy88LcSKFRsrnLui
Uwv0wlxow+pBYDsUJYME7yH7pdKVwLSvRpSEI5s4wicQvFdg3XTGcqOVd2ITDMkPHJostuAbOxc2
25+TRyCtDtUEab3cK7rUIR18DkHJQCUxSsbJKl1hP27P3tL6Jg+Thkn6gY+q7bbZXc1Ujbaov4pQ
fnnOyokkpXHM2twmMSSyMnJ+hb2xVGJu01jJ2XyCCJuqvdIOJbhdOm111ItR+BNv5y0ezeaMROFR
Vx7McbOeLheJEw5VzZFjAFDGHLYBvdCWMl5YaDI7MxUlGReBHXSg+dRSwvZ+k/Z5rhbFd70Remi/
HzfMl4ehjRucenc0l5nJwmqMfN8UejVPK3KFhMlP7B2y2Cxf3ZFzeEBV09wQH/lqQ5cpKqcjfmMj
Yqz0b69pX69MC7kE6Sm0lLSCZgdrI4G3OBEhTItN10kuBOFdun0+z85qttTp9jh0lU7rNyMUaAJL
jWPacOinY+kMmkXnJMsFYiptbrKCxFpNjGdSKUXBaFwAg8IdR/Cjd3lBHnjJlGAhmrPBFOOGt38y
LBJuOb4Bnsy2rwBibjDS40YiXFnN8OHTjYuhtxhYZOsoYSCS/dttZvHLSNNvRMBer+GC1FEROhUW
ef0CmolVcv2MxPfsJe0t+J63DQIHL+SE1OSr3M7V3QDo8Bu7WytYPF5Qvw+sONWZbgbN/juIV5kb
mSfOw0QiUiXoMArHbgFIOw9e7qGdUf0FxWFKEYWNGnJKfSSooJS6ktFyDRJohZnZwtzuy15NRJdH
pXAZ2z9M499GNEGkA/3YUyv8BrMVuxHePAvgwxtG+fbhV4LUiYY6h1xcwx9Qm4rjGG5dvZBWw+WM
SbPo7PIadTlconF3AmILkeNYW/lIfSxOZTOZA/FKN4Ueg2hYiAsyQpC3biGmZePKfXGm1Djdnfie
vcPqlfYC0dIYsmTuIbO+PXcS+rV+pFuSDifMOt8pl7hKKCZrHcObYJ/5imfEAR0RTYKkzOQmUtWF
K5hQnhrhh44VIInc7lBFQVXpgmOb85i979xowSvH74Xu/0RcHsDBnhuKhgbmFiTBE81Ut7gB8TMz
4tyoDFsGkfYchZ8CP1yO9WJwSoXQvALwULuGXUfrzugQdKwONlAtU+HvnT8TeG/vO5gFskBd6ODQ
dnerYTs/d3DePCsICz3HBZDNzUZZyJOgc7cCyITThkoWlWX8EyPfwNOdTNhD2JkcfHls2bU8AGXc
gukwL6TwDBJPmcA1uuQXbdfttzVyOaRu/rGV+seqBQPh0W4ov9aSEpUyrHVpcf0hBl0Iglm6Krk8
yGSkh0G5OUDneizoywfKRkeWViTrN6GThFDftiN2xtcS7Eaa8GqECWhdcihojBMBmA/UoLefTD+C
7cYtjVJMi7SlygXt9urCipKWZuoIFn8GrEI6jMONSKH1ldgvfWUWhoCPgCAWRr2FED04YRowhDnW
JLegcC3hP83e/CNnFVm2+szTdNz/ioMtKF6KpBPNfH8IIb/IXdS0aFsRAYCLWqodcMz3OKgkWVvx
pYyBkhaTR6tT8p6s1DkbdjrgSLH8l1voE6V1H5ufwQ+1G5kteIloBapbOdsL6sFLb45UPNSaFROy
H8yv/mOmeVIX1RPlqG3xZLCG38IMPAKMcY3JWXVKi6mdBwgHsHksdN1G4N372CnttucdeQk3FQEH
WsWtgi/uBOqXoapGy/sdUA+v6P1FYB7mGmz5G/uV4wtPXimj+KDjzcI0KH5LUZOzASeZJhL0qjv+
F7GPwP12/vpD8dq7IsFjmvwh3x5D2R2Q7sWE1r09c2rHT7utJTa72EAD0Lf0JNUwjD0wcEuYWNn8
vNJ3QZzY2LkXE/ajlHaZFRiNgyeHBOHsz12kvFMWTBUSOZYykAa6ujRxF5VqpC1cPKJGcg9400pH
rHdcdsyZOfAdUGkiiGQsL1CjNOW3tAKqapk2YJ7IZzvI9rI0HuDotMclVChltX3cJxi7/B1Ar4sR
mkL8PeQoZr+L6Jy2fjzNiX2ZPk3uAB55hiTB6k682R5/tTSkWDrbkf8aoX+1v+IssE+F8HNb4z+H
1818rrK2+zCOUgps1krtn80fF60SJWHC4Kno8iFDCa3xzhtbOhx/RnIJD0fwccowXhFbR7/K0azi
qTK6thoZyvwrHCPx/QNobebrP0IIh7m+1iSjFqZafCKGzPbIhZZ4qPTc1m+SXBn0LAicjt7wrUaK
xkFqIbuYrfRAyU6jDC7aDPFdCZw8+sOoVMse87C5rwr2cGy8sU+yRaS/YLN3SfVKbc3S7pG9u/PH
1nq+kfAQrmprcS2sQhieKGI4k7VH4xtQjkG852zhRjlyNJfkYOC630FSMleHK4mW/F8H3OQWuc9c
MJGx8dLqjNOSJfuaai/IEz/A6UM+40baFOPE8V6FbOpMft/7yALpSJmWyZu6OtydGvKnnzvuPM5u
ioUU9u+mHJuUEyg7aYLlR+BllsKpT26cvOApc5DeQZRFPcy92V0elB9Kx1wnVlZ8GzihGaW8/JEu
IEsdgRtwCXjHwEy0XnUk+SPszBr4M655eNY49z43Xe+4J3HSOo29yWf+3+vVDddVRI3A6uOOR0C9
D8UQquu8Xst9VtNB78OPsXskoF6oCZzKHat21If6sdoo2MEl9gEm3HvAUvqd7YZUK/yjs/X2oyng
eudU0jzap9JSz6zc8dzpomh2G3kW7bejsdzNnkQ1Ug293iNlQLNElHCwZfkgXzfAQAILfoQMsYRN
S1n+o1O1mYD/OsO/Z77ZbdHBNahHfeNJMM1iKUhB8fC6rQpf6E6irk+vzYBw+B0m73sEwkCXfIzN
Xmy03BnoBDGYkbnCnLA5dFEYPLk7xawJoKt34kRE7iQcB7LqQ/sxdpl8wSUzmduZ9v7utOlsqrPq
XG4nAsFgzEDomhzvxTPty3Iy1Lp7GhJrCjues0lc0J1igeRaOQtRVTkNqoU70mwoSVJr2I4y928Q
lnB6EPEgmq0pAfiVFmeKEago+RrvKqrFvcg6MEUxXEOA+CYQDF6VbRNftZ/Fn+r5qunRnKCzXW5L
VNwChSvvpE3sdJ+sAC40jRenXwfcsAqSRtpI5Zu8MddrWb+q1vDRdWcRa+PADVR28FRjQ12v6ilm
u9JUU51cW5/Xz9U/xoNh4ljVDEufl2sWmRp1lfTZOrpHmnUeAEIHJxzVGF48Xf9ihwTgqNS+cLor
Z02j7dIHx2imp1wlmR+/AE6yRPCfYeIE8qZIPVg/cSo6P+xRnJuxS/tdiRDo0xFliheiYcqSe5Mj
TX6T40zPaS+bUBnLhM1iYQ2nAsbm+QawsJLw71U5JKtpxHNa988P9vZXXnRyQPjjukHsA6jVd1b8
OVrYgjC2ZQ/DIZlNdR7JCWfqZr1Z/evJnvAbaB6R0Cd9AGzc3ZCloEzzDDkWP/lBDGJpIjrO/way
hDrZz3wq888eoX7ouIcx9gGLwnQE3NR1/ztjCqTsNLeJK/s39YKHYn8dRJeaD2e1OUsxOU7X71tO
jioUdpc4DCQwymM3t3pGrpy8kbZxWygjsT3YnJ6S7FSoeJYWO7C4zhnxHqYIH6SPXcGXpsvCsKol
rJoDLXqWrDPhc7S2UmtqhfH326tbF+mNx2nClGrIeHwXcCiEDewE1QpjQw4lv/65va9+xUVHC7LX
Zff0ZaoegAnreEAQcWg7y8dilflGutz9CkxD/aW5S7JkJl5Sv4ZKaDlt2eEARmhr0nd0f6xMomPW
xJer2vHIciDE+FgnnpSYgRP9jDvNiJbFSMc/mW0xaPX3kBjaRJeFNvk5FNGQPdOCl7otTzgM60fD
DQaYa4jsXYDoFGHMx8TD5caFabaOiZHoW3ux7x3MalUpwnyc74VtoVOYIBj5IL8h9hJ6qqy2ZX6n
O3yPc/31NTOqDPn8ZaHoZ6IxRbv1ZpzjoJwd7HwQApB5jjA3LpKQhIVOXRAfQzz1WYkTuZfpxaMk
gTlf5I9wm0o6WNhQR3wexSBsdCjN5Q5MePLz6f2eX5ELAXIUw7IXkeEOU7HxU92icslKRcDjDipN
2qGKJtWGo3jx/wj+n8Wutd4+wRMZNspejaGqZ/L+sAKo/Nv2NDRDwBXNGgimsl3eI9VB/+3yTEgK
wtlObHguagaBex0N2HsrRovCEcDXzAmKS9ZHhDi8X36StHYeObWKgPguqywq+cNjzd/16zVk0eyJ
iPSQc+7EDycWc+zMCC4NPmAxkehyLt4txO/abc8FW80HebeNrw/xCopLXmuaEYTH3on+WlSEsXS7
jKUn5erAeL8KDhG89Vxegei5pnf/ejxGULJG/rjMIlSzB88ju3kLW99KrhgDs7HQqc7JXiHmjA/E
WiQSNEUf87q4d2UnCLS0pc+eRauFHhpexYUX5gCImwE8G7AHTRQyxMQiQr+yXqex21n4EipGDrRm
LCxbEZlNMqEuw8Nu0fN5NTV8HPbP5pWxYoMEqSZZVnKbNabV+lBQ5jZVvszK/GUjJlejm7V1kWLu
HcwY9Aj0p/znGqHozYcpzOeohSO8AMEWI2llyR95+Ry4hyg64S1B4ZgZZJ2D32zdxiSvlKodPvho
xipePPbxyx9n7EGLbjN7LfZM/h0a1zLoyH/O4TsUYSBOt+xqYtmNc90+tPTb2nCwofUh8wnfuTFJ
Dh5O0Yhr1rgSWILLrr4Mq1fGcLyY9HKIYBeFgUXb0dPQWjuzowO9rCQJRQKJwGHOlCt4962jWK/w
ajFLiDH7ihpcqmuQ5PvDYoaitSZiJfAvYgvN72Z+vixadKvFe2NyJKkbPIYruLSiNxhsgLq0HW6t
s24rXgOc88R3r+VafnyW20TMR0oRnxDWlKw6GtsJi5DmoaO1jzMIL+I4x0nr9I06WSeGMP+szRj/
AZXP57rYhPZNPrH8U+3bGhRbZ9LlCzST1423o9kRWjSLUa6AL/TFG8pwjxHBGYBUOrx1wowCG5vH
karXoEwBYTZ/EqI3lhvomADHE74ox83BPy51W0/dwPtCyvRXP5ojIUvO+UnVjbf2ZyDxcDmktXXR
0u98Z8vSz6Cqk39QQTntz2GBp+nywc5yoln88U+cOt8Pl0mF8DxnMQNYPhRO2wtDbaCwS8m625mN
XbArYLEuzuhrOJ1yBJkiSgfVPJWorOG3HQ95tzn6Gl2ILcpaPXdXLdmuXlLvc76erUelUEAt2guw
zrBbycNM2woceWKle8i7DolBrlW7l3YQE6YOMbQM6RJHO5f8R7HgDsBvXWDpD+CuzchBhoqWe23h
8FyQrHzux6DGtKFc6D7xQQCXibhf0hRapL5x2y5ftmCS27X/BUfGEn64y928BGp9eajGFuCRQq0S
AQbDLX+6U8stdYojcY/h4amnEatsR1yTeR9K6MjceR4IqLbRA1bykHL+R0RwgPKf/hNxcqrZjmPk
WuwQTLAi6fhg8D0MTGsgrDpEdypCcmVmmUyDPcgqN135IdhUO1I5Sq4lcfmlihoAKPMrA3HC67KX
hwsAHQeDE/Ol8mJwK+GN+IjZE9KpSg4i9rbO453oPZtz8jg2hBZ6I1uqhwjz2yH0RuRp6HjMmHMT
7TZ9tQ5cBWWPHK7sw4pwWGojAwK5EmuwCvmpDPZvE9v1FkYgdGbiJ0E4oQCli3GZm+kOfcE1yaTU
MOHteT/zwxHtgQWSz1EuhCgi+KigVtqMzfoh78XoLUuK/8D1qfAUGV20ynniipXv66F4B68hjjKr
Sw0wOMQ1OJ3ByfYjxwe9yiaANhBj/28z340jEYiXxV5gaYPeVoQbSke2ggb5KTNBRaPG38m+LDwd
1yWdbkF13at0IeQeWfwBHCRRkzMQAb1zHwzKCLQrah68LNEne6ZAKfUphk+XeU5WM6lIybEcfStI
Y3Bi3zVv3++aBNL5JXfnQ0ExffbtKEQ+zeperso7bpfPWWyEiVJe66q67/ovE5izfvHtA0RoRGo3
Mts+312E05JTu87BiZ3ZWQyoqpFfj2ED/7MrUAy4UE+HLEzvMwkJnyVjDE+EU4BkA8AOxooCqbDu
w9lSGJ1EKa4764yJShrAwYaioBmUwDI0OZUp9ie8ZQXjdD0h+5GafXZrO7fLOTFqo0Pv/P8XplS+
soY61g5etfOs2ImTK78UaY60+qx2iXOLxIcmSt7022TQqpb45t6PglfjeiOoYMlLjg5j9arRRTWr
YG8GakJxZzz0bhbawwFae84TtugdY+xtpWUhKZfjMt6rTyom0iULJ5KP4vOyeiNLOhmryNlmvU/I
6yIsFftgKJom/1imclu0ifcxcbwdR1yrLpiQlcrcHZBgLFx0MsrnqBJKPgJNEPvRwjJ2zRSPsILH
s2UV5KN1/miMde/YqNS63bnu8EuTPch+ZZfYaj2+kGajQ9xuedMaFo/7ePmAwSZwyxHbzC8UHce2
4w/ZzrtGq1u0ArZRPDaWhlTLDYnojpqIW6DxNLVw/3w04zdz8izS2orDGyvLEz7xD8FWTeNl+rKB
l0oAvQOQfRdc1+tdsZlmhZVgDsqevjWnDnhNsM2KyPmHNmAx6FTtRmn76LThAN/BRkkuQNjaKys8
ufpb8s6KLol2XfEyGByc38RpRSGH2hpMTtLgiNEqTNsZAgApfzUY2YJj1e9DK0LGL8lZwQvhzT3W
NdD+bPOMF2M1hXj4HkfExqHsryZpYEG2zTCxQwVCQsp9JReeFEqPM4/MPI4djVqeU3/7dVHhKhzP
3UVxo+o+PVy9/vtgyVBcl693NXadQdnDI//DUv075DTNpvhD9SFT875pwkBYzTwxs+WlAe5SjxZG
PJmc25FCVf7dE3Q1qsyd7Y0VUjGxTUmh5kYPaE7c3/0vQvy0jvsxOl7l/xy8G+bV3RFJyyNASOEr
1LzWlUXk4JeB87VPZ8vyAEKprho1RZNLSlwI1hFujGrszmCc24Wwwmx05yaNgEJ0A5I0GX3XIp4Y
1QDCc6OEXuwQu9cnDGxUgPqhIW3mx6FQaB6YELZfGo2R6FikVyfYL/ai9Dal9s7J+XgbTgWel3Lg
fVo97c0emAvR+PvL1wbbfgN3LVTNmARZsipnZDj11ReXmIR4jr3raoEZakV2z4fryCPclXJVmwWk
YkNj+DoJBGOl8RMsTaFDBnjlaAzJNpRO7oi6lDJQGe4TMt+sULp0oKEncIWpZWyM/guuluZLnY3j
mJGcUvFFY1S2houEtz3rWEYZRwsLT9kTF9T7+hGRG6LTi+rm2uC/35NemvT0xcITE5A2ZuD1P1v8
qsdd9f0588+6TLRWWe64Al7xXraIjWRY/rrH4OdorOt6aGbwNuwR8aVhxjb/iAYgNdzv5wfoNtF6
m1hw6LwRf+0BRMtwFMlCI1qMlfhCJsJzwsLtR7t8ik60omRZQuh7VXKT85zQaFczgyQ2OwDO/wgx
gbEtwBbI+MD9zfi585tmjtysGQLr7OA0CCPEdk8fpd4i3owtwe2WMW2SYm9OsWcqJ9MdQ01o9s9v
2ur+OBYKrIkAj+N9Fyd15vjcFD3Ll1vN5rsZluPkdSpY/jlwGYWBGP3qXOmumDCH2WWnZZK3v9HH
um867wcNJn0PzErObJsUqwsZVcfOM5XDUB6nzA054hjSXHyt8RO20+0wRtwucALSGU46tNTUUdUa
815IEl3xxfVbAea3JwfnqgxBcPUuFiaYBir/U/k6e5r5xnWrF3SgaT8nIoftw85BM95xAdXn6F6l
DT2wTIPc6wNONJerXT8oudRDKkDyuJvuWk1tdecDamPi+MFx5TvPZI+3Y0kfSjBcjvcMMMU8X0NO
mdAOR/spFnlTndEnJq6JoeWrmhbyQJi+7qUbn89MqQyIgqtdiUl4FIbyyLhWAIxEjsaZnmXzwwVR
8vWkGED8rarcX1P8AdKiDYC6ZxMEu7KApysZFQPy3JSDmvXWPKH6eNp0oTM4tBETZRxuPGIvLdzU
mRBb8NWbWbdvr+CgDFkVlWMdqhYhIGEg5XCzbw0ywbctj8As5oaVcJf3pqfaAVXQKQz8eP7yScFg
66kgUY27jqJPEjTIR9cYih4jpBTmtRPUkvtD2WDw5VBMhDkAgIlc4CJuDihPILUVh7TM6ci6OpiP
OVpLB6dggFq77YwDVb5PRJCITHhgGiTrH0WOfdMDVRenuB1Lkn/oW7ZM+qIQZJcfy40CGhLk3KrG
jjZ/b5C9O74KRKqb6IVkBKJfapOyqcN6mbhSeOZrS+iPCUa1skgZASaFme1pOJARlfoDJqPwbhFe
XZ7OD/87N/WuS3r9ajwzSBWnxSUgKyF9Gsr55wPI6Vm4WZ5w8zQFR1xE+YqzKQzt7/V0MAkVfUDC
YVkFlbKZ+8KOupAPL5kq0L+iVYnv0ne0Hklr9e9q/DnHDnM+TwsbAPUmwFvNeE5G9G8C6T984Feb
4LSr0oHccvQ9dlOwPavOv8DCdgZaXOVjX7dYzH8dG5GVAHNLZR871r5q4MR8HT4jdxC1PT6oGfyL
8TZPQumVonh6RYkXzhmD4UjSVL7yCRHQ2qcgEt/593fUqgRcHj9h3Yg5tw9BvxH8tj40gG7Pbceg
A8AqQYlYN9m4zNpQvQ3c6msjXXK/+p8uNqGEWa1+Rzn2DeC1gyHNOPkN8tLPLHB1lEo+9OULq2qx
rHEag1Ga8dYbT+WwTQWKa7QyRMXzs04CIckXvtlEgODv95hVRVU1uwt0KU91faZyJrCWYO/wIoue
9pv7mvhMwPA6LfFZTYbpsVByOdFNKw2gPT1ddH6pOc4uOcOC8S7GtHVTM+vzKTMqSGVPr94frPke
+UOophfG5whH7vuhcG+GHM4mkDfDuAriHtOSiO6BHX8p+MkpcFKg4hPFNoJiHVID0NPS+4AuZQcn
9p4vD6Ab8Ufq+QJLJr3dLKBEKVsqRIN8BsQO06DghuFeLYJaLj8qhtmqymFY/Xph7Fn+59tsIB/i
IbYHvQ4UrSiVKtFH5/aXV6U0XUkIpxYnnn88I1m522iFunII4RKlAu2/XV0XPvr3141mMqatyH7u
UUybJasSx+ftKbt/ZsY7qKiXPd+089BFUQhR30XPEYKEa+edszRbMRJTpgu4ypnFPBW2t9JF4MPv
OvZrksyUqSm0XphJVtCI2yhGSBS/e7svbc+L1xsr68NNFcBwsheIlwmAXs7IpgHDbpJTq2c/kBDQ
AccNE9hR6ahkW6w7PW9vjqGxNoiUMEcaqAPK8ELlNmMPBm//jBQJqljoCeMTahmOqSQGcx0fnmRX
c9dF4pnEaQKQqJUzmi9ofUm9HDTokOMWoMmX85RxE79N475mEAxEa5tBBoc7UhOr7Vu0y3Ncfxos
paBiayuRAb3k4PsIHkyadCBhSet4L5iJ2P3llouvWjGuWNxOCpDiU5GAOjEUEbFg7Dj1iLxMkd/2
KYaeVRDyVRq+QZVE6uAP5VVFaHxG4uUN48x2qfMYEVZ777vHiTHAzm05SUxDtOVdm7TJBkzKavbK
p4f7K3BDzmgJcsVOQEjY+kZ6YUfIMZbAeE31ejEbhiOyJ0NghXJmviu9ytRkWxZms51P3VPH91EG
t1lFsAyymsfwp0IPvt4vXP7vm3c8u98VavfrOlaZlEaK5RLxEigvmCyISj/6b/Qvb1qLzT5tueW7
U+HpJBZoABOTNfd4/4AXgGCSOF4iy8KG0PqEm8FTCYX1CRG5gge7hU9QE7QlQq3t5OoB4xQqd26k
IK7Qw5Ruh229fOpsAkO0wjyOwzGbZVVdSxVD54+DTYgaFQtE7z2AINzapFkEG8IjGHUFpAeFPTxQ
YUa8t2R3sNSwKUdMS0xG9wYb7DDimldTbkYeY1lfAi06KVuthTcpPj7iLQPv+L+ksFdC5pPF26tk
qxrVEU+Mt/2vGMykGbWvUCay2MCRC4b0BQ7G2zNYNoLlHzvGX3NKHwJzJ8W0/Rw2Uqd5wWsiuYdI
PzThYHCrRGkPgBITRuA09XNrSLhn3ibgMPj7MlP1kg8adw+lsdLt6OzB6FwyZVEO4hhWfBxW2h4f
b8HhmpD02OUi/BSgEIFWzO/dZzZ3vyX2LiZR96dxN3vDzhcXCeEh0SerZR2wZjDwHbC1w8ubZ0oB
UuZNXnHMWW/1UyqFZNNsPsW9uzzYHd6QwwdZgsg5qRz2xMC2ZtEPWgEA2chlew7zPSSGGvcOFZkk
kt7LZG5P4PqeamumrgmGw/Ge6XhAzCpnBgmzG7XvJsHWJBPmCCCqnHsmd7586hQlxFc+s+oQT+Iy
kcot8Gp2ENw7W5Kv8ubuRBQ30+/wxPMaVlRSFo94T23x0y9f+2i8RZ0bCgmh9BQjwl5p3YFvdty4
OK3mHLvyIdJzWfz6fojLCE4GRtVm7gxJMdoUbbI1p1hV4vDMQe4efeLaMCeQfqjfwzToO1RLndIE
rMmqanRP/t34xaR5EVK6TQklM9sJYAVqdsMNEXsRUdv6irvPg2ROZf80J3BWGGbCJFJeewzf/ppr
w42tXKy/b3A0NZrTqoXZ7pWFSgjHgo33k0RskcJ2oG3FGjxCw8B19qIp2+R+sBR9hsEj9ubgeDE9
F2OPOaXzZ8QyCcZC8jY2jJU/OHfTHYjc8nZwdwku2m7NmFk4jKFiFATECtgKNYhUML5elpNwG5DO
NiTR3k81wc7Ys2he7jLvCIZfV5IUTq4HvnYaN1Im5lDsbQV/Y9N+8JRslurXGIhE2UE1YyIyWej5
PIMtgnoDW7C5taecf9zeHf2mlmTrSxbmcpCTOWD6TnHzKqBfoaFTKvzJYIaFXFJDmwHJj27uVlHm
KrGMQ/KoJqzDH4GyBOvE/+upAL8wk9nF5n7njbVXfwXpC6qOEmsS0sOJqSCCII+Sz3XT6SmtgrKk
H1LauxZjlH13bne0sIxC8aaTNIhHis0JYvGrIhJezzmseeLBqY28kywSMctPSSJ1IDvPFsHmQHIO
EWa1NjBFql+ZgIBMvoIwCf8BjVLbhZfnhUQOePIloA4Xe2u0VRSueWrhs06N6x39DMaJWjyWE/5p
uI6AECTgtNCoAgYNSXYryak5y7iBd0Bzrix4bf/GzrYqcFrPT3Og3L49bmR+0Ml96nd4H1ITW02J
A0ca0Q9Q0URV6b4nJ/tI6z8FplMhi42SuWsdsDttAYxCw/FLAa7X17L1PCJfLMAUFEDYbm14Qgvx
TeQi0GEUnNU7HqV62e2fNtLTzHeM9tA7+DJOLd1BwWhpORrwlaFePvUAD3P6KREHMOLdOC6xw27h
Cg0Go7yOVVPodg1eRVwGO1zsd5i/y5T5OgNJwQic4OAmVo8WvVKf2pcAfITlWxsT/ktF0uvyKM6P
a4WJ0BRkJPaozRJoPWRecXvArev/FwD9Z+j1wEuH0+RUHUO5oOdlrl1Bk7cUSlpwBwYsPm4q5gCz
IaWx56/cTgu3oE4+8h1f5D/aRhaOScBP+fCHj9w/Apy+2RHKF+z7MmpUvf2vA1rmN3V01/D8rpTO
E3AzEud7HO4QGDH2cmf8Ap1tJlcBtr9ON/1Wg0j8HxoTQQlrwg+VmiCR35+ySvE7sbwb9ziBfSMX
oCJTc96dwkTxXYhTZLDJiOlXkGcGWA18WEin3rXQWAjwHdjfE2V6LQsr6QHZtUz5WUm5KRRuLkbI
lNDA5TSLEk1CeqjcmaMdAZZIVs2fWvU64fTDuSf8vlZvyHQVDmT3hlf7eeZrcLKF/mxLzZCpVQYr
bHa1BfQCB11u/PD13S3gu3RHlWhUAqwMlkt0HYLk24JY0HU+rsC9VkAKNWBuOTCQs8JX8Rc26GzJ
2XZlTukIGa3v0ynwCHgmXfNA1oD8jemnvqpDcF/3tgmHJG3tQaUnIdFEyjynigllVdFNxWpiEhk0
/UlWVpqxkKsSpyC6ud5RhSMK3hiqXbVmWhibrZ9iKqQMkM/mXp3ASLUck+WJ3Zi2QpeUSKyKUz5Z
8uRTydmaMd7QekHmzksHBp+oZblavS8aDk8J5TfX/6OjKkPYe7S9VhzifrxZGHwfolvbZmAarylc
EN8qPA+8J3NFcYxuR+WDOXw2ZwMFfFx7aUGELOYfT0VsTTlrTZGldaK+hwwy5zRw9EgMTfPi1WBX
Gpx9ZxBolhGZakM7Ha8R9J3ThD0lVDeqPboOZK0URIoUL0awAL16YzN//x6N3Dc0wJaoIPxkuePB
AZjddY46Zec8TB4Xp2N9RI667EODiPCW8K8FFSgUiGrwgEQdW8vpLrW7lJYD+oL8bleRw96I8EP3
BVZnu8Zx96Hoj2fteEpOU1fYy3dSlhRQrdAYhUHAo+T8hRCFODF4klhAw38stziQH2ghAYIISzAV
urSNuMluTcbLpSAivAbw7qaANBDW/pmWoEd/zY00jrfOu4/x/Y6gOmLMGD0DHWX9zUnu9gW9/iTX
hVK3WGUw7srjanrdHVmFQ0VTo0mlFUYT7iUKVeKvzeepcGtTCF5fFO+Rrf//r9aHUf6pZioJgUtp
O6HJfLZIeGZ21ghrqDD0rvvOsMmrSVWkcSLpgcBpRXye2FA1XGJKBe++3bvDZZLOw5td25QNyRMK
elWucjwzbBcD9f3xBbggZjOQ0iM/i8+78Vqe2NnfzFjXs4/nmLmalEfIN5psDy/Pk60t9ziIxWwp
mfMQqQWYbePSlyACe4b5Emkxx0tj+1gZMX+nDGJJ59zG/uAqfxsfMtmrmY7/i9uPcpC9x5Xg1z+f
DLGmw1z1OFd2RuaFgDnPS6W3uSl6NarWS5LXFWYAEB2NVRgCOY3HkRVxI9xLCrMOSmcUuyXd2/jO
0X3j4BDIcU0GbpG9x9MTUkFQr3FElTDme/WuIkTq3gJgMBNWaUt6/21OaVzb5DyiBFEPsnbJ/7vd
cdO3PjGzHaa9zkZYTEE3pyd6ijNDpywoQ6wG1X+qI0irjwP2hx+PGVJ+1GWBqebJhWmmN/f4aH51
udYJkecE+h+uBuMj91JVz0hdAGzLkEREd8jkYraQtzKTugWVPdDvMBQv894oChB3Byu3/T6eyQXR
vYhfniL5kCVY4yeH2m341LX9mKsoigzFjMA6IuQCuVO/ujcqo5Af6FsmiQy3spoQxMYDP3yjvXQr
rnPoI6OkRDfSZhPMIY4Jbee3R3/Yp6x/Al3/+QdmkUqOTQbHHsFN9TXDIZLE0rPOMMTklLj+Uw0Y
naI37uKZEvUbQRGNXnV1WheLuoFkzmhoLyLXHMboQPeM9PTN/VOXHsmzI+C7kbo1xuz83xH4Z4ej
SDLlmpDbisU/b+1SG4P5KWbc4PV8xAfiZPyKNkIAQP8qbYCftmjJ/rhtGqR9sfjDVCDMO5YXp4X4
vUh9FWz7L+GFZPnrdKsMS2ZhqnzTaXwuQ//W4p3PCqC3zJWrWvwbz6R7qo2J5z+lGZiBwrDv0SqE
ymj2A02XoDYLVkM6u/Q04EVBLa2khIPYNQ36orm8fK8gPjF0NXFykbevM2jvinyVmtsMqdEHbO+8
NbGHE5KqjVqwxTKYZqr+WCVj0J43Oz/tYv63ovVxKHQLGWBRzP+0BoA4Z3rCO5HITg+OzxPRr3kY
wvDMeq58tEhfnIgUpEao2WXD8PlE5detdMCVELqnTuPbBDKVA2Na+CBdq6qwxcYw2zgCbCW0MRDL
rZfEFsu4QDnHZwt450J5cPD76VN7qRDowOe19diKzfNurUu4tQNZ4SEsvpHUB4i3rZpxu8KQhX99
LsBwvv39aTSvVWzg70sYPBliFOysBlpOfPeFUR7b/K+CGeVS18TToRwE2b3lkCNRP6UGQjCJe1zi
7lBXXoFg1AJQPk1kATjmfMsC9ZqKZHJitooP8KPHNahzc/uKltoUwM3qNVJPCWNnzvsymREQ94En
pJWabQj05CHCW5946PfICmtv4Eo52rmXcg0zLVmYty79v2U1t4x1/21UR8l6s1L3ZjNcCGpbCBFs
eB7FKlKJTLOLxwd6JlbmNnMkA4WhSrxIZkp0fMQDKuUqHgqv8Pqiri/SNfLh5uIugJa01uJWioZe
yC130WUYebOdS/E79pKKQ3o8EEMurKQrF5QiCL07+Q99ZKP5y7bx0O89ugS+4cgdhEjDlQfQYI2q
+tu73QA/6qvNdcIC7vJzvcSjno12ZeTkzUzxa4dJGOgvryUhOtBPmv6XR5mY7LMYz5WS6Us1m4ug
2aDoG3LRxMZI+NuW3tPGMjbxCUi2g8ArwQTFSZcde7Yult1Zg2BYSCDj6H7exoAcVhxX3nbCXfXf
19QLxBwF/416e4cs0cZreFIhnJ1IG9L+UVlVEXe/DgDEp5A9YoHgMqwIuo7QPr2KlMjROOUQfAv9
4QYOVJ8h7Eaop9gltBiA9RzoMPhNUWlsXsR9I06l3WYPypouvGhFg7giiGL4O52Cr9mN/U4yLTMA
oVN6CBiMLYJEuwaqUVT5bLVcqbLkTgk5YRx3/lhv8MpiuASP7dnT2H8tYrq7jIk+EihIV7cspEKU
Fq6UiDmCQkuZ5QqDULaDPRnsaVQmIg8pNnhx2jP7kP2ctoDg/tDwQvmwqBMDDpvCfnbWkPi990S+
/gNPoi/SqlXtEF/ywWi/yXROYbXmxxM/iK0qqQJTYeF/R6mLkBCD3C1vtp4UoP6/uB2VJSeXpjrm
V/g+PFF9B7+hRnEFY6qYWF0zi4e/CVwzDSpLx1sXUaoe+jZeuprGHwZh11Tbt4sYemAfEEn1mpCf
5LakQ7gCKMWte+rDXH9PCsOkXLDdlijc6jiHwhesc+0Rl2tWqy3i2t3Fhm5NsmcFXGx9emwo88T3
xZwSQkiDTqOWpg0u7wyd8vjYbDeQNp2WMPYW9Tf335lIIEzEODtRklzUomAoV3vulIP8jZBOqAXx
vnp0LkCunhZXLTDkeEwiKA1QRkoKc53Bxrsz64U/LUPZ8SLWj85HUXJNUd2sf7KD0ceuhBNwqQQz
2zgwpzq1UJk3UknCwkoBNAIdjPI+34gKftF0UbExCr+YZ9CtmjWHMaKobQY0F8LL4ZEwCjHkHnaU
JmgGQ+UEgNRgCAB1BVtK7NtuyVsHpGeoI7qkSNb7CZUytKefmwbV14JrHBgUBKWS3wTEtRrLTRU/
HZz4jI3IHVOZmxZ3CT5jmNV888iwty5VUjKhb6IS5AOalNCwJfdm4WZhpXJSSH9qJNVdi5YOqubz
/Iswl32uDvw7vKWFTLq/Ub/COlMxEh6lrF1QIcWAiH4/ZiS4Tbv6vZbw6pM58jFD5cK6A5epUCaA
dexTKF3BEgz3YtwYj/qhAmx71zizdVl9cl1rzw0YRY/WyXhxdbSoH/XL6PnaeVnkNeeLVYFjREUt
s4xoTr6oRgFJ6u3pbDZa8qEIeMSxvS9O3g5HTaKbkOB00jSBG/h1uZFVqMmHsUTsCaYXIXujiABU
R+4HVngfAabviwSYJLp2IsOwKpO53T+oGHBRRVWwoPBIkiR6AUl2uJ3kKj4YNwug3AP9L3RquxGF
37WileWLp1s1KzHwhHuiV1BeQEDrbgEnVtFQLEKQtWYuoBgC7QngqBIVksZeHO4h5d4P0QU6hMkk
2DcUyYON5cyYQ+ra2zBOAu0NaJ+BWC2OvNToYvparTjq7KiwCXZWz6S0jnzY5uGlCrHfivEo5PR+
08VTs+Y/hyvkMDuuKuLDc691SMc+7fVvTBmIMqqsyha3QoVC8Pcsx7ytJ5QEoTCO/q//G100+teW
2VXKgg0YLdcvvYNV4z5ZvVw/Cvlv1BfK2x+dXiKZw0+dxPa94Tc+LuCx5zORPX06CEBCOnIUb6DA
rSVyWoGUqrYNkQnit/7HJi0bRgrElq2w3D0NZRitsP4oFsvs8wTzxeMb5kKeIiybeS4Df1BZ+sM2
1oC2Gl3g3v9K4nSRXvcHObJqW4y9jzopt7PMXP8ephD6LmsLfpIYRTPrGX+dAs2N/pLiA8UjWLd5
84Crh4wn+IkyaKuA8RODnmWqituukLDPr7UqELQuQxfn2pRCfTDgdFRphpaJSV4XX+cOZExzTKw0
y5YMzOE2LJZiaw6TEp5Jo7Tk/D384FdDykNzLdCPn1JA1Fw8PrS3pxbDuVj0QU5+HBN7bZsrYwUV
vzgVlwpdJeKZWVZj4mABsX+N9pS3gemdXtKlc8NgJirNIycBfWXX1wB1w+ShPkjInuLG6GwGZvmG
m211fgQ+dlLRl/BqYjd4AVL7StgeI9aaCthrlYdiIBa1AmI9kGML+MxUEYUsn38lpUDc5NtP/77z
mvYbuxBSMk7oIncvWjkhdoGepGLSQbBxy3D6Y7SlOZAAVRtPteoNEBDxFcs7Pjrgpr+AGZSP+Nww
d+hikroPHOmu+iywW1IZHDuf/XAroVgvPoSYOluaJfztHlrR1VkRhOPF6V6ETK5sSDOWouwaciZf
4C2NY9vs8mEpuXKaTWoWqidFJ8KrqkipcjpQHhLP2CVSk62OTkHzUDKDSU+040OFeMNJoY5dlY20
lyXwY6I3zt5kOucyOGmsoxoZDy4NrEirFv6o9tta20BlO66T/iGhN4SeOUhZ3bcItS+eoNkBzIhk
tC4M58UxMofVawG0kSVAt67E7QhBlMj5VeoDeNrh4xjQsCUHg6wSuQ4LNEkOShA4TnVZih4LL6II
nwWWgD/t54e0JwBOiaHpgEP2AmHaHhTZfDdnTedEfr1weG7EMxtN34qs5P/wxcle1KBgp+OYFjRJ
T+PQVero9vi32nDtIHDkM3QqWu+dZdp+9XwYnRqRWdY0a+Fz80KTHRu68P214hTANsD+xpWlokAh
iZqfC4oqSE8MATVzmqeI/IQChmkcU02FqooPG5UHUux984QsixM0ExN4qBSedsK73UCmTQ+YSHwY
2JiSs9c2stDRdCzBEa/wbTom+OBaMhKZzhTGGVd2YbJ/wk3ojoFnv8g6E8G8QN/ZqFosVqWd/KG/
iCvyRPdlAW2jOtASId05tuIdb3eD6U+D8l+buXYCzBVfjk5yEbvyA51xq6aELykIO0HSMx5qufkm
yTe/dMZLufwFfxYPLkrmtk27SqVOs2KZEcRPfir0wldkk6wOO8E5o7J9BkxgHiVx3Wa/1g6jxl/T
YL5fQDrtX3QsOL4RBk/s4A4dFrVxLYHzyvB8H9n50CrfieU45bfWKr/YlV13U15nPznHcKb4SO1w
KgiQe+dijuphJ+MWRpTHLm2W1LJVH5GyXiYwwQrTt4i01ws4QRasQ1wibYWIRTFKV60p7+N8qcLq
TL7feVxY5XCAF61XkoPTvkZjgX89IDg4VfS35wRATnHrsIVWrcUlud/UjVDXHKQvWYNUE4qmKHA6
Cd+pakOJ9SHh2412TiGuwj3zA9KpvOOiRobIdcUcD9xO6YJ63GvfrtYr3zTOfH6UpH42KRJA1wcX
tr6ZXBO7TlqBisFu//O2nG9cPXoIA616LLQB+mp7jefoES3SP6F8irqCxZn8Jqo4iVvA16hMYL9O
dNBSxC7ViqFQts2IkQdZxNRnTly0FetawTOHcI7oRKJf32cLLpUsaWTTQnifTsWUMFV1Efun7Ll7
BuBTyWEJ0l/NaNIlyW0ZhYapGknaH8v+oyGn5XR/2p7EGSx5lSgbEEDLPpIHsoELNbkPgAj6tVCa
kI8W09PJ6Ji1SoL7yQerQ2nnAyaQzU2GN2W8Ep9KNh29HuuzooYhtWJbpY7QTWAq4UihW+DPR/G6
0SmPOBmnwe5nAppfb9P+RTum3IcSaCawHPpqXBO3fwTVvIg2ahp3xkmW9MdxDB4PsQbpYs4IQuBp
7z4GhlTKKgpw3rm8QY6frfjoVyiVwGgxqfQP1dicOcxrEjXecHE/mKg+hB8QMgwUOGLAV+2gW72x
xVKFymzx9nWAoydzeimdVviAiUbQ5gFBPt+343w3O+Mx0/RikTClslU76RPbOyGme8vfEUOpnB3W
DPMSFuIrswt+xqiLeth2g5qS1xJ+qzug1d1EVp09uUCn/XRoabJSkmooTz+Zh27+VStzoHkJm2in
wU22ruuyweDjOuFNEwmB1hn57G6vacYNPKYgnHmsH4l4Tv6DpGyQWr/LG3A1g9gFalSWE5i8fEkJ
BbQgkSS3LrH/G+4ZhwqlJc1nW/qo4hJ7YTjNX9DTKYLs4CNaTRo/O5b6s9FyZVuM8tMsM0fbcvRd
z2mcHz9zGyMwgj0i7uC39UZxpDPU4ta1cTUpHL+eHQXaPh6tB2paln+w7RWMbYeLaQ/6En2t6N17
4GXP1qQJLRl4o7WPzgu2LTPoi33C0YxD9Op9watL79sOMp6uKoa26Hbm6R1RyU5ZHsTncKZoaCAm
i0JlIfOq2JhwzN8lOPay0ovWersx6UyCf25oPggS9ChcdsYjg5+KtzsFVjiKwK5GkTgR/8PeH0Ot
BCoSE+BMRgUjYzMTlE6UeDr8zudD4ZQ0rezt8N/E6nWvTYp0WkRxl72rUJDfHbCme9GoNZK3CLyR
Q8au5PVTlhrp7fhsg80jqrst2/yawOmQXjPhf5hUojZzyMSDs6gr/Zjs75Zs8dmpkxrWoWXYFalk
knX1iSP8JdFaN5ZIPT2+Ocv2umAFZd4vbpTpAEZ3GetZjlbWdjDlDx8BMSxdlqaG88zDRVEFNfZV
7OgG+XDlkuPcAiCNeeSsvDL001R+OCYJ/N2NUeKkpJhPpb8Db+la2+eTGug9YbiWrM9GLZGApX4X
VNT+qgHKm1yol9dhgj5aA8ittx3gz4J1CaKqe8wf80taPDxpmyZt84RJogEmQoRTM9OOXn2y0mp0
PbhjBue8CpYYAxLvXVSn1sQXWLjLmsU1ujHB/1fUGMABYTD2HCrjGlamX48YdH9zGLMEj3EWoNbe
Z2NXorN7kwMlajDfJTPxrh6xqR3GTXUIn1gKzgeKarIrWSWz9ITOIyPZJSwz435YM8AaOCuvsLF4
plIBQGJW2GT10IoIPs4bZA360BLCjCDU8jZ3qupW+l4qe8PeBOarsKY07DT4TC8umczG7FjfoCCq
RZ5ye0QhHQM02S9qPxrSucyxd94zQ3JZZPxfTInLEudP/XBW9/qdX3U1FDPMG9hGWeJWFQP1ZJ4H
QJo8iOEc/F+1DwdK465rHiT99eJSmRzHgJCPZ9RLGj6QCkoFNhdm2u56DVGk0eoC6IOlo5lHzXYq
LsO5f93HQNNda8mxz1deH5vDOnH3cJARZGWjd0IBjc5VpofxCewUBbT0ECobRTFcOBWl2WbjnYzE
Kw0xszsNJ3XC6G6QX3O63rl8cHaIOTtKxBLHBrXqeaWd7qs3rHHPNj5W/IKJpd2fWzKdyJqafVLV
1yIy7evX7Wjzl8LEO4aJB/oRTGxQAECUTHquTK8X0XwT015dZ0Xi6CV6+1rXgN+ONQ30/DQ/hbrd
mhxJTIvxXp6/lO/t9OwdMlooL5wTVwO3QWUUI+S6AsoZR/an2WAu9/aOKRfXuAyP2tfKnaeqTelq
0GEmC2xx44hlX93H8Lbctyf09zWwXH1LPAmV/V2rMKq13gqUnJBAbBHcoJbxoUKA49Y0FZDqb+LO
akGR7Aby7bH1Dqyd8lsxs+W5/Ao+SSMxQIIqFUpv9+KnUx+cbUHElHdPNtsR67gLO+zfQKgresMi
TgwwzPTRZFNDpDXfGBYC11VmyzcrKqwUMK8rafE4SBooWIRS4aYm24TeNn/SmXBXFawe0GuTmak+
P5Ce4YmDeV5uZPDsnpGr4eBLphQwm83GWAOR6SmSYn40HBNqBLGpwylB5RcgPomWbCDlsC5w3lL5
gJhSc4whx+cPqUjl61HEwRA8ca67h37nBOJUPO/wLvI/qp3NN3iVRygPq3zKq5MwfdGR5o+zCZ7n
tbYUMtMIDGPKKdvMPDcnbLijwGM9OXeTG/Gv1fxLxBZ77HTcxYDoxoT3Ofx15ZPdY0WMiXu63UNB
zB9o6N6vlD/qByS/X9FLNt2vWPCLDpQu48jDjaxtzn5gN1bRzHL7CwZ+2hrHxLgBubxymF0lTVgP
vc3R/zR0RNUGy9qLApw6I3MrRWCScH0fDgrragWA8XIWt7CbqSdbNhp2J5x6DmSpDDGnE1AhOjR8
JbPUbdnnG7r3nyBwHyuub1zhUdJCIt8OTMn7PadzqKEqaDudLPWQcJa7xnxmP2SEQHjUnrc1FcqA
dT2sRx9DCn8hjbDsekKU+c00yGc/MmJBA/5MIpXoR5jAkcOKiB/TNX93fcKCT0yePI27exGxEOJ7
d9y30fiWnd5s3syzd+nycFcyAufSOLc+hSdsdAZIkeg2hVG1coGHwvf9ObmcQfOHNitFrVTZdX/Z
Wly6l4VwCko5O3nmhMSTqX8yHjfcYGgJpQmkxK/0M8xZDthl9eaQ1/Kdrmu6+pATvVYHPtbu8Fst
vrg7LJUTZJIQ1Bu+6pZBuKj1/79sj5A4u0n35YHY1WTIVdu7SLzFPVtJG8s1eFKSj/P31zs1wVob
s6GQ030z5xlWZ0J2zoKtTCY/nwzxB8ED6K6X665+FbFusJ2/4Ew1GV27FHEVppCH9gUwsb9rznsq
TBSgL3ROIekC23/AVWPT3ALZKRVC8s77u8qnpgr8kyn3AolrpPyt2N/KGR5wgXMmcoT2pE0KDms2
2l1HCCJ2P5qQMx9w0rNQ/EiyIlks7eOnpIZ6euWDZMqWN86eh+sHYo1EGE4o7jBD/zlIqEZDAFdB
aUo3/airm+dhpOWR+WF3e8Iyl1EBdmFBMe7b7r88nymFDGj+r3tlxnWp/J9JymRgzV5w1N7oF3QO
3/8/feJo3Otzw/riTbd+FnZgUyNvFs/NiINz5tXe1cxmUJYwOj53cYm4Pqxs/imN0zwLFt2FqE69
ijF9WIEHQPNNyH4rueabL6JntUWkDzXKRvH67kq0lm6qd1ZJIe01/1wbBCItfFebkhPDso3fokyt
Er1fRNblVCpxImedOqR0Fk05gOfaHgiEna8gil0E68hyCBQXxD/tixcHpy56NiC7/04or+dheCpn
gllV2Rf/sQfffBr60BlPg2Xk3WikrBw5YKM8uq5YSd9GaEPSbpEBo3HAdWlSQoLoeOAvNzangwsd
2IDNeGOSd0PRwJng3re/hxwgj4w/qk+NCGep6H3CiYtUVCMTJE6BGszSKESG1xgzqYjgeeywoM+F
iwe06taoh1QPrNGXp1L5TX4DpNOpxb08E4SFVXiqsUfFPWoXGXogDlOtgsOMu6dUxN1xfQaCbYcB
ccRsfHuSbB9utk8h43XizWIPMjX3LJ2JKbftKOtv7FbTHWxfO4KH7idmVqGGDqXia+l9Ia3Z8e7m
+IfV4Zd/DAmz6kJ8io+OmfGbxJgUbF6dB7tS4abiFKiR1s0a7ud02KSCywbFUBC9aMfHUgazaoKV
syGTQ8uS4ucg2kXTPIweIQKP74eXZ6XJeuaa//3oUf+xMQ6ijznOmFgj1sSROpCK6PsaBUujW4Jq
pr3Ut2X4RKPy9cIZVfckLwLKCDHH5GybiB+ptdje2865fZiN5/A2K65dQjyJxrOwRrFsN6H3Z0A6
zhgOg1tQYFlaTp+oxEFbZhIDubLPS8pfsOHYTWS+9xhH+2eVBLk6eOlfPbVcuExXaioHrhEqAb4E
ThNJ1DdsBa1tNj+6PqgumXZJkqn65l4QTu0xz9pT7h5X5CZVnhqHpL8OxcCOI6OE72chZQ2zU+z2
Z6ZLL3EbKwcGrLCAa8N7fucTZpqSjS+7akYCFUMY9NGzL/b3cy01i2sJgDtqQiTtbZg4fLp4wimI
rEMlv99G+BeQ7w/lz9wPCXytGY/PHAb0Nga1Q0STAG/qe852Pm2ZAivAPwlyU6SLkupMmS1ZaCnI
Duk4vgT7BRjgjEFdqszty94rQuWm19hwMdDjxqqSHKu3EwvrM32nR2JOewyxaajTp6h4eoN8ganC
tdoALBpjO3oJbm2rT0qXovIpqiFtjAtCF4acK5qrqe7rW3CGdE0tb+bEqzlHI2oDe6a9Q0TGbKEF
ZnNGwog/7PkvIj41NqukGW7Uf/kRVoxAm9jD28OXchNwPLEKHJPczHHamgeE8OMcqdAS/mc+N+tb
/3LochAJ4x2Ja0cONUVr9QT6x869ENlwRPNWaQXmBz/HtM1fJCPyvH4w1MgX6OlmlW1dYzvs3jcq
z55Kxei0u2xR+QH25aTDKJRxTrtE5gB+AHxiKQBl9k9n79DgQyZRhBErgbKo5wQzTSNs5S3P9L6o
FLhc0xou3Q5l+mlXs8JX8pz2cgepbF2mOJpSkr1RQUNe7X/IS0O1OylUzwzoAUeG/J/XH66ExJ4O
ErNB7pXBLrFe+TnmYOCRhvs2tnfglQNC1ExMLjiMnb/B9ioePYMnC0AmC4douAax8NHt1D2f5hDj
b8R3xbHTcGJeDs51lnCGavb4ZWlWcOMyHnBH53+rSwVqjB6MT2ukcfkgt3e0HSNpOtTcSJKxWCQ3
xX5UERulFbhUx8l8tfiAbOzomXAMi2P8t9vhMtMA81St51BLArNfrzz3r6/Fc2xbZ6jUSVBxebp8
YFWPSlVr0ednkgcIX8sdHpLibL5QAV9RupIhRZtf+AUeTJ2xMTb+186kBep8n3jdXd0HmJNT8/gY
CHXCI58T8t3fGoAqeQCtKPHjzyAjCZcbmCgLQJNpQK/Io6rjxO1Z8VGq197TmWmJyh1mvM3e0vit
2Gmf9JwdySIFI7sQaHtpnz4Ii6bPT/ymafmHIIKSVFD4BdW0+ZmeFuPhmQHQHyTGtlwVyLebBXq8
ZdpyTiRLR48x0tUrvU6LWEIpXYq17oYbyl9LabRvCTLhTQBPe7qcfWVwXxwWvAvqoWWW4NFA+B6s
LoQCVhApJ/qcyNJo0VejjSTNVzGfxEEqF0I++DH7oG8tys/KNCq/j+FcTauen+6G7d3ftiU2SVl8
Un7QILFpXk9qapgIiI7zGfNUH8RCk71JuJTsDGP2f7GdSROdp4PRkAfEo35al7PsMop04OC84+0l
fAEU2zgb3pdthcTZr4C21HAybMMZjtFYS4haodwh0xIGAigvU89DRcgPawNlpShGqph/HUwbPRgO
ouJC/98bTELUIDwqrXo+qR4VAH7V9ipL3smONeuNrP6D5inwzDvlu3ALMF/HScRppaQKrPZ+UxoO
Y8SukfrRHG1iioesyG0EXweYEZu/StY6kR8s8ph7C+jyFCOtBlfvjnSVZ4MBzbbz9WHOiRZtu0rd
ut6lhnjovI7B8L5/sySjNhN9FbWQjagzadEFwtgjAsHbRY74x15zXd2venl2VwDcFWsrtm0jtbgF
pgEhhTPy/9jqvd7FiCC+tDIngQaqc5a1ttRdnxaDBIO3ymMekDHpmqeXYdsbR2Yq+s+Iu1+SAa6r
xc7MyvN0OR5FKH1Thbgv0OnF5zcv4TudAq7X0rwsq9lSQhRCw5I9iGuawIeD+OXPpVYdVPO8oNUL
p/er6+I0QobAXW+DP5XTcwx87dlsxs+P25QCCS8jMv0xZXAm7cCxTnXBd/9xW5H2OK0KmhOqRVCf
ISNHaQw+k77Pk7RIMoe+NBt/kVeH07lD/ws5SVbaFyfFXHE35ehNpDu1ssIC1Y+6gqWnkQq8EkJD
+jL726sU+3BpyazlUgOoGSHt5oLYpeJ3WVakOzNBVER49tbgGi6akitHdj2iJU17LXm6Bs1CITQ/
/lCuGssddTCty3ck59+bvaIHS0aUEUH6kUVg0GkpUmLKicCuHJKxRsHGqgd/7nf/Unx5Vu6MWuY1
VkpaTzNjoPml/ntmoq3/TOlO2KhL0Gri0UXGhBipdW2msVkBf/IUlls3rDgnnmWAQYWvwnvIqrIX
1OrYLl3D2lPC9fUqA4r472AYOTHoUjtdB+8Rn8BxhaFZ0JU4+/irM7VTmIgVAp9FR9H6NZ7ptqmd
9JU1m1W52ztu1YUwTXbPghC8jsw+Zy+VERCchtInavqk4W9PvrInS3bs411UFIbzXwtxN3xUqlEY
/28rKbYbsf1Jzb6ZlKjUlCASqyByORsThuokSc3o9QhOins8+ozlglHNV5r/aEDm//Xt7brP2W1V
BfGwZCoJ1iuYlKIMPfiaGK5nNCpR4xH2a1WP8f5UDKYKOgJ0Cap+PQ72wFwjMxUxBuVkazC0Dwhl
A9rmdQE5Kj4FRQ+Y7GWYUO8aa9XVdGm8rlx3eNiYmXrx850CRNevHR3TDej2Pv18BraFQnCAB0us
ieR7BwighFKGJtI3Tk0FqrUAD3sJEHjnsjGymtgX5TkO8K5El8eVUo5px2KpmjT2HjpPcYsFtXat
1ajDetbGan/FUu8AdhwgHUgPbDRmOx/yGGy3IcTXELAoLH+P5eHt2leVvDQs/GtFNpOUukjkKBbC
YjnYTLEF+N24xf2qh9zQRufB640ojdRVz3dqD3V2wkmCtfMbavMKOlsb6dSE68IQB4R3l1GIElYp
mw8slaOqLXYwlphLeCFa4kkqzgxEJBngAaR1Ct+xmApapYr8xESm4jfw2iTFWThxWyJcntzJhVLR
oAztYqpQqFyBs+riGzcED530GYkCZiLVjrurWilBm0wUTvjTUGecXftepO8c1xHodPHBdI+yzZpi
rTaVB4BAoCT5MxhrxAr6XLJREO0z8b68pGt1VD0qLLAC+DSVoVi9xPZtYSI9K7+hKiC+I/IiSFZ9
A7svGGAlvdOiQaIoDcDghKfjq933mLhut7C4s+O2G4BGHQLNo7Z647QsLoKWdlm0U3t4C1yHJl6l
zx2477AKy6kFd1Emy66uHVkl3qaL5WS6Zm6SfVztdeQ4khvzzBZ2+w9E6G7yC6uHuqGwc4IXdZoO
mw1z+pMQQ31K3hNIV6J7zqURvTH4FfNfYxlJD5QRESuW772RDcVOYyFYeB+VP20ZpMBM2OJbtHGG
7zyGU49XlKUuQE58+5SratQV/sRFA0y5j2NuS1HMrJQD8vhcijtKJlcSCTNeYUXup2fcWOpYGXWI
ROz+joU6Ry42F6yMFdsZvI4qgQgiN232sR19G1//w/dbbJjzDVVDUgJaYCXvZKu7aGdHcdExgyLb
9KwhWoKfjAUgJAT2881LEb6dTbfe7ls0I53J1dHQcnGxZcq2R6wpHYqEEVCFmKzDFshT8A4XLaLL
YVQkwH0MoB45FT7mdwrRVkYnnMgznn8gAYs9aPWym6Fs/T5Yy+Ph1Pz7rhaIOvqRP9mtxhPWfcFk
BhvKc1+qEG+fGs85iBaq1sDEZjutCSkF87dvyjGyfmuiNuwdKhUyDELTrukbj3QfbrhyJkyIoJrt
STVUF0djuqV/auC1iVPdLqekhFKuRG6Fvd/5fnoirymMjV7wg0L3d1Rk/lBT5fmcnz5/1i1SmRnO
F0QaQaQ1pm+zt74ednCe+qLO5Qk4QGfeN3V6HlZuZ+8mfzGrywVm6/WCRvOJNe+pgIBWIgxtCqdJ
4iGWpSfVwFoTV8/TNVVwdbnBt0Qr6/e0buKNjMkL5qGalqC1iGWU30XRaWaOAb0j0g7xiAPcBbPS
3x9LFFAi9qhXv9hmYLrRuOcOvZoLrLV1F7DS/mPxfhsW4KAFoxzsCg4as1dyQO5JEHXOksEpYy2o
4ZFFmoQIHLMwfsXBESe5/kNfELJWkxhbgQeY+7kedJNysx1y2npU4xE0N+PM0i158Qj3gU9iK8Gq
Z5y7tc34SN+7oy9kHM3hLK5VW0wh5CyC2GC6q5Ns3y4D4YqVMMRF9/ad2eoK1xzKVFv5CRDmpmjk
XnsrRahZDmM281IQHl1zFz57UOKkmsxVOK6T+QwqvrRU/tA22cewoAhjYwX5grA7D3cVRlX7ydsi
gW6HTd1APBuwPAW2TznAmlnXv8muu4S/PcrNLg0O9GLOevzI8GUN9ppnoEcnA8BpQFK5jdRwlPIe
E/2awh9BctgmzQ7eG1HU6XwGF7PQ+EO2NuzENQTuiM4jtRH1jJClGhL/wESVyfIDeq/OcCKnUYe9
wWTXq1BC3X23zwycVr/K0ofcuv1Nt3kUMnBJDjc9pX7kEt1lTxNoQvMReXlx924NeMSM2P3JxFez
TcHvm3E/0i4gwNi42G9PFHxmjp0/YCnrMsB1w7o77+uSN9zUIkjFXQb1uumhc9bnQ/UMerQWCgHN
Z1gnxHttJShrOyjY7G+aFUdEBokJ1KSOBd1TNm8yW/ZgorwQQQVi5QrCfFmUv5U84FD1eNXUnEXy
sfYrTiD6iBE1gkUuR/7hOWeC3YO3gRNTKJNyu4jM3y+1FBIX21Fuhrix09Yc0c0+IxtIiiwGUFHg
G+kbyyy/poZsCdSTrYzy0eXKAN1afahC7z60ZyPSLmK9cr4IPOm5OnB6Gvnaqn4kXslTIyXCLN2I
AWEfIsMY2I6/dSrxBKbUZI9wU48/KuulFrs47875e1duN/p42GmZFyn2FjIXwo+Vb2yCXMF91fkP
54qWj5y9D2nCBPrnslBkHGeaMFeGm0wQCDjFEYh9zdWLfEhgQNpj6M4JU/OQGGAqo0ojEf44tZmX
ywIqGJcHmlkpZZOj8Wd9L6LS0LnvsLvH4b8IZffC92voz11yVXoIclXrBpbGLnZcMBx0adr5/5Ia
L5xUuuo3Z/+x9TEGDqvmmIHWKhAB23nIOgQydUeypLevp38m15X/34F2SI14cXdac3WeAt5lJelt
9bJ5VgTqpTNO2bcARPfqMft/6uaxYs7j/mTBdyzTsEZp+/LpPKnlrRT+GeOaSwATIP4TXa4/omV2
oIfR3nDNKdY/g9YVKCXHDaizeZdIwzOvA4TlPZWT2ztewHJPL7ml3r0Kd0OD0XgpVM+w/7Td+fRa
mGPJvH9qeoNIeLyYMg7RQVFUnyt13xXP1U8Uw2qRFUvjy8xTveal8LuKzM44Qp2QgAypPqaaBT9k
Vf5eQ79h8JpuP6+YbO3opFuYiCbfSajAqnjNa4g5ypnLiLjOe+emGFz3mo8s4J2Jon8B3Tl20kBm
0e4ojQR9VRA/YFZmuDdFoApAQwn0Ev/uOOpNktNR1+z1aoO1ayGiPhTS6Jvs55vofyllmxuh/tn2
QMh+d8wsbUFKI6nO6NQ7Rj0B8Ye+6KHLZ5EcBghjKGTCiozwNYYDgrMrrVuFXVHmfh0JgODiVFsA
OWUsH8NKOifQRmmXJZwIc0HY7WW9vJP2h/AC0uXM3xtKkTZ5S42Z+ccnFE2C96SanS6FCIl2jpA+
1O90UqTpgfP4IDPr3KaALrYTudQdfD2tocPkC+ZTmej6RjU2CyCeS96YXzUbs8PgdXkl9cG4UnwV
1NH3vzkD3ub/6VNEzzV9xttStDsIE+TMHRvlkgzzkwqUBdsu6E+H3iwBBCDbTtLvQIkA5Tiqt97R
kG2IMsawQNoMfREUErQO25rPLA4RnPH/fYlgM0RJRS9yjq4mCr9QuxEhkwPb/Ewcz9np+/aKscem
8qX3zk/2CIKhcXCjnZ3R6Ml81XaRrwZAZ1sMNesMAH0vGDghBije1ZS1d0igMqj6ycDuWVHjKZ2E
4y8fbgvKtro8pvDmKyEoCrKEbdl0CvlyixI7hF7KcX1Yq8Lr4qPiXxI7JxOHY7pvXhc/mugomLDo
oTH+jUg42zSbOBK6yf2Vnsq8oSOjUkU7fv87ED05xZpx0SARg36zhfU9rw8vYRlRFxs/hiFffu+I
FBnQx48FUQfP3mnkDVmvgd8cvS1OW4LC+/S7w9heVF6pG4liTCDCbC0O+VxCDFDUGIPm73+rf4i9
YjA+bocTzhB5PaSivun95Xh8ucoQFxFevp+XvZdmwJYU+UMJAdAMmarLssG8Qc5GCOfdu00wzEBC
sVW8ZYI9Rn2PwH1PcSKxTfP5DdkzKksm1xAv6Zq5UfN3OBO8D5MqGju2dldYGPhpTvPPdYxH1nc1
rN+qBzWwgstHGMQlwEcs2Auad9pTMDzVqScB8ghuEL3sx7Wq9FjYWgo5UOAo3C4FAPswVZf4TW0v
LghMo4LIKYVgfMCyp7bbFT04tkrqY8cF/e87jMswAoPd4dndyxPtSzHwf9HFGJjyDk0kXAFCwC7R
/LzdoS7N8QjRrqGN86oDKEjpLv3ksr20A+SZsjzpd/5+Nmir88LP3FjgYUhGUpSoRa15/ub2ZdP0
e/WTlm/sRy9ApcA4LDLt+dhkW/QbtSBdnM8LxCkRvTZqE8zvRpp41Cs+Tna3AOYKrYTB9puV7xrC
S6shVHzyX9HvgXgI65xIqz6yF7OB6h7XLHf3eNsrnBALSEGOh2Tm9AIHDIlsQYM4tXJFu+KAuq2I
b8B47K/06b59wYa+/vX3xN4carorHYsMfLVzA+gDmZOXnSN+u6KHo3I8chXTyu7yCUR8i4hAriUB
Cwo5ntCnawNdX4cHe2k8HP4Y5D03ErbjYO3AHmeQm/kRBmkBr+9vrjS9vPoGSlJCP1mQYdhV/ET/
V6O2uV7xMrWp5s1M0H3LL4NvFc0jGfpDjr82VpPz1SjGwAVfraO8QPMSaVokfYj2OT+L5syphsHM
bpIP1Y1nZOhGE58grtvqLgb8gf6lqAMrJ8aG+C4Gs05vLE5RsvskKZ5lqpegvL/eFaEt9ZMVDlL1
w+idInXCXKII3rF3Rj6utK/CjzjbPKZyy0InJcY2sUeof5Nvq5zJfECtiGN4lLSYNDrNYva2bi2d
xYmIucXdMQP016M8FFrvcLUT89jUtMj1X1iaeneHwau+qJDixNLuCAr0lSm5DJJuyAwQ245vBaTq
Mr0wltvFvGNc1pjVEvCnuTBYz4r5dZK9v8bwWqn3lLGjtz3gADFi/Pv11RgdjyuNjS5lu7nszVQU
4fMI9yj6VNvVsZf1lD7EAn/Vf2gnNUAQNCRcAiG9aNS8HXz5A0Zwpf6RImiiBLQARfi+g+lRqE2E
9BAh8ET+iXBde/LeNtx/YX2YyBuOFqF0WVO1+Nxws9cDO06dQGU2507t6ZVSurZ0zwjFm0qGGgFN
in9WUiqLE2DjjQxt3GF/T9kpgiAvoLnjbVjSqm7klBVH6T040j4xeY3OQWFHwD2m5lWsU+/XMyCT
BNwpanFGZmdPVgL0OMIbzUvYGJw+DJEMPfxWXYDt0g4kFP0MCOFUlL5e0dvFrYZGbxTb5rfXf76X
ayp/DstDpXVeJBOc3ZEftfiQQdoP4XcBkl4OxpQUIqXeMD4yk9Od0JwHQXS7fHcvcbWw63RqtQzU
zQzCBgPqF2kZA9/EPeUzTCY/hafEZehWLOwryUm59p2+76IIHr3KQpNc/YyYMULT8Id5ZTer6eYV
69vmhg8PyWi3t655E7bW0Y4MfBbuPxq68pcpEQopsTev9ktPiGNtn2AlqgH6SxnTW6c4J2Uz5LcZ
KxjTl/CT9ymC1d6DgomehTA24nTFUAgnzyt8K2XCsemGy2FX3GEhbM/8jOxfY1pmVOaJd2muynK+
Qf/0b4LfYl+nTBf9mfRhIcMGBCtAKjIDKJhRa1P0TX2lFcTnOh5fMPVffxVDXyDKOsoxPtpbbCsm
JMGeGB5W47oa70N49qRslyMLvmoqDYx7RXvNT7lcjHIgX6shSBdhZYeMSXa/TZhJmMPFvqjnAwxM
pSmRq8AChp7GKnIIdd2MFrF0VIIRjQ6YdfqJJmTScNAkvoz5vCb3i268WIg2kETGYbY2N4P8Xb3v
Zl17gDyht22YUtV1cDZP8Mx22ItuCIMhRUH4gafZ99hyNwmYUXYJ9COo4fsjwA5fXf9BDbXulgfb
Cr5XZxisSta8XwTFhYsGMgwS2hBfmP2p6J/uelDsbKxW9IU8CgWgcF3QojHBbSA/1UjRG1aAZMiK
gOnAWMvJvjUSY5BFFt85plMvbrlq1hUAaXIRlRgM13fsxXufHcnSTyWoEBKF9FtMCh/llSSiIoL3
PW4UvPT3pazJ1XJFBOWfkGpzj2oJKAco29t8gFRV9AReUk/1VNJunPG+McsCzOsGVQEZrayEd/gF
3KV8XQYxCMQn7ZPr/3N5JCWMMW4EqTynaNAQ5D3+1I7MgKcYuOi852QoNUNF+RBMfOT79ACyNgB8
RQQ8RrYxfa4D7/BDo79wzGIoGbkCvTLoe0qoNhoXiTc+JYVljBQzQLxVSIM1vfoXFqKQOIk6T7zS
ekfceeu/nZKSk99WFbSPecbZrST3shEd/sOZdlphdXOEMi3sFHT5aZtLX1uU4INaZtuOPtSdg7VR
Rdh2/METNtcgrhS8XPPAIJDn37XMheq/eyzSz6fdf2zNgRH6TCEUSCyDokSD1275sCXKVfLi+azW
Exm8u9vNfyrwZR9XAhHEUODlG/ovQzJmdCAaaUii52Z+5k1NZyM1b4LW1j0D7v0MdJ4+3Tavi1Vc
2GrA/9+RNqHEMFIgcLk3cAscbXdPcrthk3+Kiq6w22tB/6LYTTRi2UAYTBEXykXTBlVT4l2qP8DL
h8bKxxQo98Zc3e1vzP7LsL7wbfBd7oSt/3m9yyKkmdnfq142Dh28UR4L8fSlxatU/NGQwEe7ES2Z
D2rV2Sz5Cjwu/Hn3UylcxJUi9jaDn/796Gu5BwCMZ8po17R3CUcHQo2virLMPwLLGTRnReVWwJEh
Gi/AMRUUnJFkHCBFo3gAieSVEpJnKPPowcgasw7HcQVN9O6OZxX8zJ+jJyNoJJaLOdInM9Xh6OEX
C5GwNqB76S6fuN8Z0BxuY5c2GIFImIyhoxstVuV7i4jU4d4ToDlA0fkCNIvtif/DK3WWuzliHMkN
qwYsZSg42kF6UjBUF9sl+w7wOB8PBD434r5V9v0JwAeYk/yjhJHtsm+LI1BhQSKpXpnu7ODTu13c
+X0utx3//v/X5F7ueXjtPtHIvskWemHjHifaWhQkDRH7h1wmMsauo64NOQsIU2E+qV0yp87Npk0C
oqt1F0qrw5Xaks/uPruXrIjEqTMEESYF7SFtt7Js3tRjSPakFtxuwQTgVSWMaI+IciYXuDGEcqfv
uyXsgk/KHUQFwKYXVKDodoj32gSvnHKQHLDOeV8wU080Zk3NeS8t5Rz4RNqO9uld8g04tG3lbcwd
KsleTK6GodwtPSqmQr5Yg4a7ez7evrvT0xVGopDG2gYeclYK9lbG1PWpIcGseHsvTVU1G1b342gl
7TlertSoXGSK1MX0lg4Txkhr2afZQRi+WbPjmNoPX+gMuuv3zPK8gnz0VngkoYp8PLs3oc1LpRnC
YbvlAB0Lwa0oh7hj9yB8BvWD+KnEQMMvPE1f+Ba6X63y2ARYfVVn2EoobQPmP2KyFUzeMwLcTrUB
73VVG9fOamh3E65YnsiRaDPBo9yLIkYKVhzFBIj1qMolHlHWyjHvpMNumX/5gz6O+7FqX4kPlIYy
2k0FDCDBpLYXgbUIWaT8RPRX9n7NTa/gfKXYWil9cBx0UhOs/dISN81Dg7FThN1wbVLxDJr1Zq5l
Yfp9pbwKjfi1aXxwGPio4GTgKGaXWb/a/qMLA3qXl0T7SSXs6W3kk0a/EtMZ11stUxZ17yrfxI/W
rLvCVxm7itlZ6IZuyBSD9A7gbGJ4Za0+fT12JXO+rDJRgJ808dQ5IVWDpVh1hindo4Y//T7xw6fh
9SIxQI3qXwV/OZNJqnoQ2ew5Nhy1Sak1N04gkzwu6ezHvxbzn4/lneMQK3110W4eXRrTQJgbAxce
k26LA5/xfjkUG81D7YdhK46XuapyZhe2jg014FoO11psx1HdCTOoFJZxIiGHQW7dFKbiOc3Q3xuP
H9XDGpMCet73t+mnLhFOx07RejupZipq9G9PXsXbRRxCWUm/2dE2167E0U6HMSmmveU4mIxD1U+t
W3anogDo6vK6BJ3nYex1KtnuhWruhCCBMtrWzkvuPSPwPD7+Nn6KpJeR6VHcZJ0Z3uXeBveI74xp
2LXD3BwX+xqkT+EkmuGvSwN2pqazmiamepi5hDKrMS+S274krpTt+0W3MiMnZcu8DhxqpWLVzSmj
APO4qp6u1FBlnMVzb2K4vy7SPXKsL5uk+iX/vmqsgbrmShmugIOgz5zJon6NdIKa7/q0gZpE/6XE
TeEdoivnEfNCWw5zm9vPb4xR3tdWXMSrDvzeObL7h6nGqdGn3FkYrZAPq1vkcwx6LXNZ0OPk3ouU
WydjbX5f0oCKwzIqzBiPXYxIwtAN/X5lbFLJXZA5yLInOreAULwExA6nIJVF8qL7yfNUGsTmNZNi
5Wqhv3A17B0twMw/h3t+AHtbb/nKDcvQVzkfvoqqgx54pr0lzFBeUfFgZtiYRPY+tqm80al53Enc
ATnl5SnzkbKVBC94tThKnu7qsajfJ6hcwtPuIpXgGXIhFh9N+6xJYPS1FHqe0Je0EhKS4dZGwKCV
rsvkVHve2DeER2G/tlJyrC0bp46zl80UzLr5H4cfaIAQRGUATvWyJ54TYo3RXWJXdwwAd9jgzh3/
3kWAy0gTrx30/OO0iquU7fnCX1gVmSREYxw42FotS4L3prou+HbsH6im3+MyYotk/urJk3cWPNzE
1wJZFFCRIeyBs+o2rBztog2CnH5DEdLDt0MBxTLYzJEPvzmToXJycodYR3YBkfPbirxgDFfZDuE+
O9hI60vC/H356aDHtBuXZOMYNBHh2IVu2pkbF7pMThFxUBz56hoZgqSmVYcrQ3xbbPTTtAZ5NVYD
fETWW118BpTJcaKTmJWzCL0rqr8Tz8smTPaJnD/jbI73/mp98y0vAlCj/8IIVU5gxQ8mmhQALit5
aI8/gqWPmR5Pvmku7F8Eh2BF5o+wwURVQSZbl5xepMjx7ZbTK/YqTW7maj/yRA/fxmBut1m5p4N0
i66EbHHI0ZulWcbWDI1JNG8kpSKGJZPpPtHFpGiQ6ySIi55L6RtsT0/bVJKGWYhbjTUH+/w0Boha
49md2oT+g7cIl4+25x8+EdZD4HRNvScbXL4IzBp+ZMHs1eq7Tlx551h+P7wL1AyOkls4sVeCIaxl
hnlA4rdwjneZ+Q/6+BhsTmjpLPAaZ/vDireY91BD9jXsLOyN0evm1puYGXw6hq6KnBONdKpaGjnN
pu7uEw5TMMv7S25ZqhSpArtwVMIfrPNgFGXHstcDeJ/ht5Y38jtuHm3Z31gfPhLt5wLy/YNJImfE
IdtZAPSmpc8Mk0XEUu1j3+LjvhqjcSX3DaCH7SRCagXMG3K4S8oii30RHaJaeHQJyNvQSyKtpXIA
34O09utWahY4gKHArlJ6TRDEYJaqnWQRCR+k+4flnmCR9B5HLjiyC2B71VszlhIR0WiHV/h689mh
c3c9kwmk8AcdegGcbIHeTyMV/gsK5+8vTMsVZNCue4jUyUbXKHwcahqKLXPtKI8Keoxng+lGwq5E
ni2xq1PcyaVsdxu25xxwTbcOWp3UjG2rsxA1txozKxz79g7tbNsniRaQzNa5O9J4aZQD+OiYr7bj
Pq1Qp23hA2l02brYc6NyW7XwfZbc+kFwwLMrGSWf19mi7+k2a1a/ylOcsONHqgNvNNHThvN2ie2L
qiS1qktIjk7ldVRkBb4FhyRYeRG8IbvBj/toxp5h9/nmsSoVG9qE/HtBVT+VZOR7mHF38BW1tcGV
TLAz2+wlzHhVaTg+dJoMVQceOQVADWPHk9/jmBwQ8TRPjCf2EIWD9hlfi+wRn+sWPV6vZEmCel16
ZOh66cJu2BEFYpbm80IIZ4qbdhDT/VlfDv/AjA8/am0HEa8uHCmPYKM0Lgm7Ug7nFH5RbyFx+7IE
WN4jCs3ORb9El+6v3R+4xZIZ3VUUfI/AAehjg0ELQRpt3OYZe9c+fURHjw4DXaZyK1BtN9CchSUN
cjlO3b8RpbdWOCfZZs1f5K0S5uAWNPNrJEUmLbecDOr6+LNTJw8+eF5d7LezWqcQaMJToV+GP4Ga
5Wcue5TuQR1QGRLD5wKDIwkR65OhA5M5di543WupjoR7pu/jvOyEdZOGiI+/ptFTRRJuZvfxiFQq
5KFZGe56yRIW2VHvznoX8DphKrOKumcNgu3bFvEquitPeLMxylERNL8AepAn4YaBY+FXk7VTMvlo
LXlH7MhA1UihfaN8rpH8AEJ9+PNBqfOIPZfWnE+AA/yiICCtD3ptpR7VGXCHukjD6ifeVlFpxkbT
gtEWcD4UIdXVHHVXSSxTvJLXTFEzpbQ1+OtgQIGIP7IhCmoDAJhd6J76l0m/zS1vADzX+KQrf+9e
qMCSZeCoSgSttH4eFK4ZuntOrO0DkC9s4XJoiAigmT5A5BESU0n38Fe7J1I316H3q0GU2z7Gt5tH
xRuSO5yFTPE3RVRIp3Fe2+r5cVW/Fv9bBXblJ2r02tl2FDAbktGV5N4IXgX2JfU3IvDeBit822On
jF+fLfR7HO3bk9SNz6mdSkxyiUqlshvnqe4zLkPxDRUfztsHCgbHGwNp0bX058RQP0r9Kk3UEcRs
5//Wm9TRfKcr2bBO2GLtzf+4FPxuv+OuJhK9d9URbC5sSa8r+rgCYEQvz94fhR4ZuehWzlCdVJ3y
wTWv5yVVCWBZ3gQmfo9b+95V45tIR6OdezKoSj63ll3u2CEmn4qgC9ngMfBxjBhhcDmmUqvlLw+q
xqELE8LpIoV7g1U8lPYwOckYATdS9QlQAizy3RP/oOu88xmBmDf9PSPaLinS9pNHlpjGVLnZ6+It
HMRq/Gq+rumjASSOPqBsGDuYtDchi1+xanI/073j5VFZ0gr+bwLDXwzeFAnssdnmIMvp1beahjxZ
v9swx1cejLv2mE37lGsi5pcanaKjzVVuXKuMWnyhVPSpL5VZ3Rr7v8hgnCWZj8tq+04Nt0QjchqY
whgoZOKelA23bTzdMyTnmBFjWRRBXaAp0/wtdZn2S8IEDTpFK2VLjYQ/pIrrFBkFF3nqfOk+Kv8K
5+12QgsdnDKNcpR9wKMWrpO5avctJpena4kDbJY8WE8wpairkH6h5XSIMApUD8AjrgykMHpH4oIo
l1xwO90bSp43KAZZpqPzgzv67P1OumXy0MYdDLjHK4o/WSKQCZfyd3cpSovzHKy+AI4cXl7waLoZ
kkPk1G8HXjU1gpks2C+79aYjDxVDz3a6aee+YJ4wf9RVwdmGenu4jgY/Sw5qYq5Io0IVSGKT+8nG
6VznOi8kTK4PTxU9rtRstdArhqxxnOgubDvBILgkDm+zwclkXjKck1ivDU6JsMkJMrUacWwEFDUB
J6rq2mykqfEwaSlA8qYFJbOLoilZQ7gsirTI3/xopJgOhjX6BZGsjkUnckDO5GHrt1/GIgkk0ETH
DiyqX6y3Th/YwwpRDEWOxtQltTyGEVsXnH1QsJnyVcIE+gFwgrun4vUjL4RzpoGsPHIKooKWvumK
R9qxnWviiogjTYvfDjO1gaCSFFc2S1MLNTtR05bOg6oTbR39wt9yb0EvyQsHPcPvr47P7ih2GXnG
3RS/kixwam+VLpd1uC1ayyfYpMpAWkdYJKvIvMyYz6qYgvcRXPt2fuXfuaifFk+yCBJoLGdD+mF6
RlJKMqpxk/mB0y7RXE94DE6p1YrcRF8a+Nhjiv0jmRLp9vMELZRP7nn92BdUS4EFRQXKCK78Dn7E
PcQBxUJQkvLOtOSfkzqOvhZEBeBX+cl7rufUwhh1HksWLWkzQbAQP7JZrRXIZw/DhMwkUGCDz7wZ
+MgQbq4DqxHtN5pQZnYyS1TIaq1nvwWMV9IrRnQmrLM//kmiAMVwcMv7Y0zTCJ04ZTxQV7GSu7w9
dM9jKWUZICAFjlo/AcPTgeMOmDm81aYe7L8KgSl28my5wd9PSw5WtRZR4J3xAjnncMNG7n2p/u4y
pqm2RQEP0wfBSOpH7yaxQ8z1EjjdEjrYQtUteKOfZxqL3eC10M5GUF4Zm2ETxADPggHO4OaRj1p/
w42n2S1SpKPfdTtDCkHhGcSkGWQ70hRC2XU6worBA+8PH7J9PA14tFpONFkaf1je5k/a5HUX4iW7
4ZLuknfkRnaa+ZHdeeIjkDa5djC4IZFrrr8HePTClAzjkHCRvONXanU02TOTDJhfBr2RL00eJU3U
STxYQxBX/fvLMttS6qRKgGtew+wW22nYerU3POHObVfqkcSqG9/NV08DgDQ7MG2CSqu9+NPUSReT
yV2G2nmgWqxeNI+T8X2QGbe6P7BHJsfZqAwcON27lw5xFHGSwxmtYdbRMwUIQA5e+t2huOb4Ukb7
2imFnOP4b53yNUy/e9Y1XMCBDE+RNNCX7cBKf6GV/Fy6ihwIuGJzVDRjcTGrTD2t3uMuf6urGT8V
VTubh/GhRpjNQbCTqq3XL3pp7maWCo8rhdTzdhYGlk0UlrlaxvpA9wlS4Pj0LHSXFHegEZzOWo/6
x1lOBCnw5auR8z4noA4RzcyzPKPp0Mu+ZJrakYLp2WVBHdfwbsBA83opnovCeuXQxEZGvWPUkbI4
REDljPUjYI+pX8JTV5Qz4f+cy65cmlZRHtbmHp4xr6VkRi3vkTDWqaxDZCgOn0G9NwEH3Kgp3RH5
eN/iaJsTTjFPmOQru0nfFKLDGIgSJkMlhBhma7SNKl+ZKITaOewAhP4enQbQ180XjhGaPV5edNvl
7fGe5tk6QO+LZVLuqpetgskjgLemdnT/I/sW++Z2Kag/ndPWqu8+915zwjlLeTn5b7W1hwkd5Dno
BwBLxfEtAtw8q5o+5ApINb5OtN9Ohgp+H29rAG1svDOX7ZDk+BErU53bbYRIHGqXRi5l8hXofuMl
h7aNliVZ/VKDjUwKEociUwG2ulw7yNz63Y/FQpFiLt7d4Ua8cN6rYSwUHTVxH7J5pORZYIE6+xxl
qGEj8w9ak/mRWzNr1V2XfzUUg/6iwG9RDHep4RvE9nWo4bv+ypTNKDIgEzfUneGqls0PaBpWz3hh
xa6kplpt8MvQ4U0TKMmutYKVWNTstBhYsblHz34zN7zuObzF0TcqBetb+atn7I6nWYV+A4NyoBry
R0Kh12eUIUnmmp6GRxfGTbH0yFYpyzsW9Kh8XJDoJ+yrCSHNhuC4wnXiJHd73SnYJBEqvnNd+Zy6
u4prJKL6y14nRJE2tUNc87p0nSOjTcMfZt4+jSJScc4i2e+nm0++VXdIz96MWIDSnDKsF5ZALhyH
paF0sz+3mviLdNA8WX8xrWuizAP3N4Q9OXG6WAw6VDj77GRnRveawQ6Q+4XtMyosq3uMxFIkwhxC
cK3+MotFZlDjIysDZOnzAATgoHv/OPOz5l+W1fKRvN7I5zFutdi42S2tv9ab3Df+fiiLmchYvYRj
eRC2J/V1/qUpS3xSMeqTW46sB9u+nmusFNFATJgt80Mb9QEJyiBzGLCAHiZShoWzQwcIioeOJ025
1R071Ih74FriKa38cGHVPLYM4BopSKeJ9Q9W2ILmN0a6uA+3x/wh2hkbdzq5PQQgZC1JsOWbGTlc
nvK08PappII5H5IYb0WOY4j4lf90cgqsWLUPP+FaaS8C+RSSMdEFMl1trnFHDwPG6q+EboBZaIha
CH26MBunaSJvHOjqT6e6pNQJqo7odZR29zkuVcEvJZEZuXRtzgwcyLs1VPfSUAo93FEyx65oUpHc
feGn7p/ERhy9RwRik4r1PcsCnCzYZAXHHFLTW6nUkqHbHZpm/YPMGscgLv43vWRAgqZPP67gknI3
E9mLeJviGgUEKlq9DIt6KmlqG35yP2144+CKZYPU8qCTtAtcBNA6VGUbyuBjZn+rL5B223JHUdJX
Vdp17cVk7qcnRvg/DwQg6THHckUGf8zQ8E0a26aM/TUVhDwB01KgdtbBfbsjmS9ubfC04OWpvdt2
XBRx1klmOsBRbax6OJ4RkERYIsxqaUO0Apy6QpZUVKI091xJ/d1HWyorjyBLXLeOId8P05ieFDn3
hwkMX0b9VpXJ3FyLVHSc+Wo4VJW1zjlxjxRobdfhF29NOjhmF0/SFYI1jve0H88DGNeSDEQzC4yN
Hlk84MqW+b6hWHpHOeo3OZjU/C6loEMibmNihy8KBHTuR1sBpltae3X7rC6cbaDA0udP3rIOySh8
iNmBpg3eQ5YuRgHuEXK4AudVYfDoRKgUWVxoo64zcKtlz2nKS3UiP01tkZfpJ9UG4RF6YHZD3+pL
X0t0fBe/40zoFW5yrleE7XxsZhE1iXsXCYaxjTNqmxa7d8u0blC3wlJNuzlvR3vndTQ9rC94WR5b
JWpcj2tSITzAmnv/BnJ/S9xzW9yxALllFf7CfINkweB9RbnwaI+KmtayvUK6m+5ANbBKqifq6bxj
xygRyhXVQtfDgE2wVWx36pjKRW+nkGQoTRtgkma6UK04cwbp4swMZ84Beg23Bv+6MJSLzg9XNt21
aGOqEB7+uDkWHQ7WLYwGrgjlD1HFim0fccsa8hWUmoKLLO9kem7AjKag7nfIT2mb7aMZUA424pam
PDcyAzohFXpSTHeTfpXW7E6TmbHkzdU2/zEI0UwyWbe+wysVHl191v5P2vM8Z3VTV8KFai3nT/xn
iYz9bkhxGnKmi/L4C0Z8SwrUBNYvx3cfTPdtTbXXWTfjHANNBjkpN6pVkQbvElBB++HPONIaEHR+
9hOi9l1YQfWF8Hc6NrXVuhsgwQmsnJeXwn47OTWe1UYECRBqJpjnSD65FcRR2GFqmcoYyTeZQW3N
b3o4c/MmKJL631Csr8TFEY4RZpLnk5f9SHr2fXP3QqJTVwyNyCzo7/FyPY6ys2Z87T6TnIUceba5
6XqzNbxN2NJIh7o427iZZ8FsPP4apTJBZBnPNWK3e/jqezlmjbKTTwB2RYgjertb8nfWES8v+r1V
lDTrwNPYSgWXidTRnbUIGe6es9zTpyo9QW/eEbgVOeOvARZPOLlfKvl/JS51ZTXty5l4YWtU5OM9
X7fdm0l8kfIS1CWQGVK6F4a/aUQLOFZJSzqlgDbDnAAWdUcMLTNRxnWLoI7b5fiKKUvc8qPMwo1L
J6pWlVU6z8DEf+PrHX56En/XT0Y5f717z6CBra9qqgM+5ShhNu78w3oSlTp9YU6DuZf740e/OuVV
1JErBPwBSeWhvtaQVuKqGwAj3QDXEMRhN06NektK4uYI3BoAGvz5mxuC6iF7iCszjYr1RhDPPGTX
/XD1/PzkYIu8bmZ9y8v120FUDtASmGorhHhEu2jdpM+HtEgehhsSkwFs4SvTo7dKAIiIB8iIywmr
K5qlnkF7GFzsxsI2H6SHfVQAYL4h+p2Fhnx0Mx/wB9UugjQONEbO7GGAiGc8OUs56CWj0Hjhn1nn
QgPjPqrBPytNvG/57uuukPRY6etCnMc8jrJn3NrR0Yrb/umfbnDuJmOfGPqY3nGH5ySV6RLOnx4k
HSjs74Y5WaRmrf5MnIOnsTtPYWonTWpu9xe3PzEKB2iCJdK9g+GSrMSoTnYdh7gYSfFW9A2vA3XD
fMZ0o2Qzij/PMSXWo03oaqGZ62ezrXxn90lsZ9pZ9dTwbk4hDk71O0LLqdT8kM2Mvu4UUXIQNPCi
YtnJptP7/sjBDl7dTbSv2qIA3FyTzXBuIM8jq/k6LKjrEEi0cpeY2hqu+kbZa7dKJwO0Tgcis272
FWLnXlaZLj4Rw8v5FLUUQ4FWQ4uQ9lmPJDQm12c9qp4/mU59kEwbZjSZZwOvlB151dvw47fV2hWT
NCebP94vjIZt59jy6AH99c0yJojDUbQ2ciolSyHNZ3VLL6slyBw3cbtJmOTum+kFsYle31YP5qrs
ZY2WHnlosAXiXtN7zZMJyNMW8p92o7JrG2EAWU67YPhjmyh8QVDglqdcrpvnhY/o2PeEh2ob4P78
mbPfeG+I98xPwHOe04WIAsEjeW8lztTG9GH7EekAtYKNooefYX3Y3ccwb5Xvyp3U9Kt76262XyYh
eLsOLVpGVShUvqdJAypdKyPSJ1HO3Z8MfwmxkpcdWasKs8DCHYtEUoJrtdJmg2fnlUmrva4OG0Rb
7P0filg1dOTeTqOB9ydvxdd/P6A5lSE9+qUUbQSnrh7SCliC+lootJ5Qugt3Yln7KbaHX6LpmdXz
JBv8Z2vT67+cini5dGUxQXCBjmQU/CK7JIvGCLLCaVmHUaRxSoL7PPXlr8EjKYQ7zJBOr9AtruMx
WbtZL1lDlwCfNNM/vVdrFJcKmJlfo719cGiC2S21y0oMAOFCTgpDFnEDm04e9KjYlUuhqW7c7lQm
25fgG++eGvUxs7PSUjyNAC5/cBJ178FD6Y07zDKVQZTOStec9E8yqlpnAE9uuqE5DiU78D0lFd9/
HuBM36tGA/U7CGP8t3PO4spCfIBxzCoecoIlvuXeOZBD1VPax5PIotWIabfKtj2ycY9z+ibi51ff
lw2sy2OiI5HbQgpUEbmJZw8JOcxLxjYjD3gAkOqMXnYr6/VK9IYC/W5FjMeMtl6avLBsy2d9sHe+
zRCNIKkBEhXpaW22D49/vF9bhEgY0SO4ZXM5uGfvM105eX1AHVWmdRQ/9iQxPZKa5iSjuHa0Lk21
OGL8vA+G3N78LIozPpZj2z2Pq8qbfvdWrDVMMmxfqhSu8Fu8Ob1nnQ5nElul3SdoMuJGKng715zQ
DN9yeu5NzlwAd9WxBJ+JLSgADCNtq+BVGE/T6NDGzIHr94+5xvVCRgLVJClIFsX8tEvA1jqMPHzU
Qws84CMCgWyHHaqqNMvwRaQz+VGa2XH2J/xhvgxk4varAeP9Z8kerAt1XYgvnC6tU36qndr14Qu+
CaAlutpcVgps8i8OK4dLz0u5poSuh+knVRdmmIIreN3I3YFb61uW9g0IwsiCav++zBx0a8hcB0CJ
UBKt0UDA4TOSb5qjZbi0Avg/lSQiWivEB5EP7dTjlpp/gaGVgGl25lNzVUWUAi/0ZD1UOdb59lAD
LYRQROuYbKnOPH6kRY8AzE8yhWgbig+v9G2nJpB6vGXYfmIID1DiF9WmghrVOaU6ccByuAdB5HrH
8x8k0It0rcvsCMLf+0dfsBkZ8QHBnPfirwrl4j/NKDJUhyOysn6+TdmJ8dpPmYkba+RbdhS4sLFv
4qCxmyeORiUonideamEGotP4fHjDleupvnIUDCnqwUvZ6ck1HiNQQOXgVPAO0nzCzOEQKXyOddDy
2W2JKK4XdY5GnXvBpmAz5sU/43W6r7V5x06vtYnlYASM/icxGTy1R4hI/0/vAg/p0BeHPY1z1C1/
f/EuAJkrqJWcRCUmBl7y8wOezN5YCqtsra0Zjsb++hoyF+VFBPkQ5vArKeqrathhZORZZCcvhOe9
P8LChQ/QiBvQvCnKpgN7duIa9phLABoj87aRLDkE+WoN0b0pG4VD/+cN6/7OC/My2KIm6ytXshTr
hZ+cjTpt2oqHyTAsU7h6dn3L+G8N608z0X1fdS2C/Z700bTk8coMVLsY5qQ06wqnhEsQYZ4qTP9Y
JzEbX3HKNLp7ruYZ+dNZNw/35AO3KE4CcKdRhl4qiHS9rbo5L4II0ow3RS3nSXZmZNLK29QYV2WW
4zc8RvpYevv14v5V/+Qr/HMiStoEIAty0CdoAD1XhalShVLaW9xexvvaET0vujcJ4aifzZMVgP39
XVtW85tiSSrgX4t+/V6Fp0DSY8geAfIWpTg2mscPXtsDamSILrk29IOocbD52WXAmbMLBzglYGD+
jz6P90PeyOtG8W4+PD8wpg1BZG8fBSjQoF3U/D8fPIPCn5GFZ6sA3feB2nFgXNU/hrNYWuXyAWem
+Ei1QOOZYvx8AEbJ9JMD50zx8f3D+YuFLPTs+FVTntlzPttUn9mryPhyYBXwmD/AnxSBJ5K+iPjj
uILYf3NCaIWTGXqoI8oTUFgIfMYUKSi0wFT64j3IYSmyrUpsqJ6Nxaa9DZQGM+lM2wo4Hz2xWhCo
9BU2r1P7GQNn0dJSoSLsUBMtvsVbieymGExRBR+9K5+iooy/Gfq7Puh9+3IjLdIaNwuUXXmLEDp1
PjDh5aMOgxHit25Hi1qOD+zonvX+9dYPNWYfhCW1EDRN0at9/4capyUfYLq4teICe4wVWSa8Hz+Q
gxQWtm8ifmzqOl0CK2rqqJFXxhfh3QpCdWVW9A760Fzsd6wVdinD9RoN9xN3W05z6S47qqbO5rXT
m5hO6Bked3zjKLFkW3NqJVC4DHJA7s2iepL9Jwbm+5OqCU0yKtpNzzPYFj/7n7D7uFACGRbEUKMF
UeQ25n2XygBLuZrjY1qYKGghyn/z9KRQAAV9msljhTEJioeGiKrx5j6dXqhgbw3yIQOJxPaNuz2Q
J4YMB5vP62dJ2LKGUeLtKq/Z6iU3v17FKg9F+0vtLvaVW5jN9MUVNM6QF95NIhtuJxd7k1FJ/THJ
PbRhDK8h6098cw1wmEMrAx657Xi4CaDsSXL+in1vSE3+9yNY0rELAz1fUS1dMK8lx5CU2EQNVz+l
vk3EqKkFthgADDLRx8aDmQEJYLoXSWT053RjfK3DT+4JDwF/ZsU/9JESYDvcvvRpKFNKTIKm/tC8
j9wTjwGgOe2vZJNlof4mN61QxKGKldGjAZ5dv+vXslgmc7+mK52RZsP1gkcd0dktU3AC/yuPI6Ct
dfHh290YZxXxIWShTHMx3qetXqACn+yarMSjn+lBmZYuGcwrkGUHah+Tpgru5/JLFrqNh7jotvZz
9Y0C1VZcybHzI2osPtyLCUNjHSjnTCwOTjqxlRVtPbAiFMS5RK7LNbJxHUJ4BCFT+dQkZn5XRSCS
kcetaOqkMcJY1tFIIQlNWBKKtJyGq7VepZUQWNPSgX6BIGDstdlneNCpVMAKh9/jpLmzVGLd22ur
TVN+ENNcNavEif56//IUahLr7tR3j9Y+8jgDCQPsXBh6V5II+pK+A4V7n62060+3ry8lz+CeBB/0
L/63FHX3lsZeNZy6Yhdr7fj06tSZccrJmOHBNEaH7QsB8RNwATb7JvP8yShq1QWFzH/thxFMiKtE
6YvFL7LwvNy7dEbWqFB3flxKQ24w85wKn5Gmcgy4Z7IpQJCFmTdFbTEtFMFoUmfmig5TwjboG7vd
L2V5UVyjC5FNvd3NLDraYNOncMiSt5WF9r40L7HHjOFqw7hMPXzS2IsiLzJl0fRRcDK/cca2o/4W
x1/+H5+vZ3I/8p7yuSEWn0mtMG4gUumV+dXa6Wdjnl8hz5WrZ6ROsxaI/NUaAF9kBTLCUoHcxAKz
XjF6oRjbMekIvn4wzM1MoN/7Vb1+UG0CHyAOEzR7QrtVCgRbactotnXBpvah4izDf4OBbqrTFbsM
S+tBArJPK6bnIkceDFYcBL6pnoga3YHq5uwtfFTiaMDixb4A7xje6GvvZPbUfQ1wsfegnkpDjHdN
sHPAoAce+k4peTUF9FskHfnAPMEbvualVuujk/Tt5EoCK8nn/uUqmbQWE7qFJ+I4EglTTezJKgUd
TMYR9P99KKBWfK0F+EJnY6ILnUp4N0YXCUHlMI8jMrwC3We1GGyMDdWFGzxcKgES9iab/8Sf5zTv
SIsBWZ13y0M+M0WNiIVyfRNwVz52wpnCbPh4SGy5oEB6p0v0CQqZxIm4ZvklZyhCrKPckQbONMPz
uOYTigMpw8CRIe/KI2ZDSh8LZ9AaXZmwXpZhgxf6ekoCD1i9U/JwAd5IKUC+qy5CDfnVNHZzgFtD
a6Pnuvtl+MlroYeqP4q8x7ZyTRFyXxBuflJoBe96NF5LgJx/fd8UJiEb6vE/+zoVHHGhyCD1Xe0d
FWHL5ibaLB4W4/xsZk7BbP1BGJQEFEwN1B/QjW5cABf5lNiqLVTwNf0dBNX40rDgOQDqMbnjtGj9
AQoXCcg6fCAb1ZS4bF3NKTv4WmwLfpiF3fJH7z8J4CID8McjKZlulSaeAVyYFt3D7XavQ3KzQ+5L
mK8E4J5i0LCD7qdzKxvdqN7MdUJ7S6oOmPf2LzH1rckdh7E2FIe+y3BWj2fTxuUvz/KSxrH6jAue
bhX3l2J8Cu/NOX+UxZPwxsH69j7YpOhb0KU9pFSA4UD8yredA+VCPtvRKgjRQRLSueU5053qAqK8
Id1JOXObuZrR5uhMzzAbLZmiITEJxraI9fp/WK9P8KHua/1LbkhEpZN9lsdhnSMUSV4raA1dRDOT
0fsmXDlj2is94n83+nCx0dodPz5D0IvlvczbxsFIaybQWtrc4Pb5+9OaOT/nYk5Pkc2RsLZAaPQV
gtbccKf6OhPtbCxfgEwq+53NDpbp+8I5YrRhHwCw+HjHLmDW/5Vxt0npT47VUcErFcICnijU1tH1
2TsPIHU/+cQJjjGNp62Z7X6X80NfloYRPXrISt7uGVkJNLIHXePmaWx8hmh0l1e+Z9eDGCt5/j4F
rqePJ1pkNEDbr6RnqQzNrE5Q1pglrBEuCoxMgAE3lr2ZO/emAVd3xKUBiJgi9yTZ+vPlDHDD803S
taGnmZdQSkngtLJFZnQ9wll7vlIrywyWI/E/PESne1QlnCiMoXLkXzBfkKeku2mLdLJ6osEthOaN
Yp1oFGHS/LHiC24hjP90zORZ/9GGtF840sRaf/mp1h0LYe7fm46xKgPEF/4KX5NgROipJhLOlVzR
tS5wd9FTXprsam/ltPkypz36iQvnzrkfp6MaD04uvB7TFFXZneeJyQMuSYFcOzE61b48kX7uHN50
6uZ+yIyGpsH8S5ghE2S5XNLL1hBxLQCcOPJJO+OQnBzW/VJTo8ZzhqXfElGe42zGZERgkxSSLrHX
gUMY0hO2LIh0LuFCONYwlOM2MdJ6tOSvULRdQ6eheAp941+uSE39UJonYq105iEKJuJC97bKz+Ym
dPcyMqJKzkBmXDsDJ4xK1VUq0oTl6bcTV0MuZGUQW1oEpaQ5aah8L3v1P20Lk8gDDBVmOYZM/ZzY
4bKt4KKmBYhKZMb+J5idYL/IbtPtNUBRv0wLCEdGk6/F0U2czLlVTBNZTRzP3ifrW5T9GcC/C2Bh
HT5fOvfzPE8hp59cniqlOjXUbG1EUYGSWMQ6IFRKPnSxSnZHGmNaFOfhd3/Nz9pSyE8tVkXQUHBg
p9CaORVoCbS9rA3ZfXpUDMCRGpu6d/qx7T+C//J/KmZARDesQ3kXo7WFaWRF9pXq5ZbjTkJZZ/pQ
zzqbNbyaOLIjV7zKrMTu23+3AwKjr8rV5u/uqDx7jjUSrGSg4W/UEhT4z1ealsevxR2mdfYUBiu2
QJAYijDaLjhiC8qMhh7TVhM+mFlSZtvRwLyBhRWp5n+upsVQUR4L+GDBecjiK/Qol9WZqV0IIK6B
J/8t5qQfh8m//MAp/J+qZmJw5inICt6TTLjaWChOHFkG2M6YOUUfWUICxYgjxiwQYG5ujVmeiMco
S5NvYi39OGW/CJVe0IKV4pFp4Thqbn8NeFc7+cGcBiPaWnMC5tTBxtE2zPcd/o2yYNtgqR4xOQ7R
FkFTGqYgDswx/Bv5LG9g++B3S+hfwVsrrEbk88S2bB3j3xFaHgxoxr1HihvbZNvoj/lrgaCsKHyT
+ZZWNAUHVZ94+A0CvaysopRGb4nyNciekM46c9gjQ8/IFJgbIHhgP0+j7FHN9xCIHkS0Kg/rcmeA
mN/eY2ANHOhHdlJJkX7iuVEKTZVbwCUIYL2toLS9SBF466gEXCURUOj+w6/46zU+E+iU4k1XAIkA
f9f17IDYlOgtAGThSnVndLtNNH+v449r98VSITkY2O4Rqv6myh+RSqNQzbm8/65dBZuAp5hD2buQ
HlBs0sanvsrThYJpf3DLrXDICRAsczMi+DmjaSoJxgeT+0EAWraNMKvSeu3e9kInhXJlDuFUR2im
ut6YJhrwmeJGgqoajl04jIchOWDgf8TnW1k7zh/Q1Ee/4bqLonaIrCgc7lyXLEQFKIjFsEmDOlnE
/mtjh8097eJVUudOYwzwKjnTTaLpBZwRifFNVlVGK4WmjWDlwtkcUypEs43YD3oFJ1NMMZcCdgly
TAy/2or21Jdl2AfZl+xnmkk03rGonyYvNmpECKN/7ODK9hU4GrT/M4BLKncittNYEcxUqvg7Qxdd
asSf5dpZnInJOXC5sdZszGGf1AtqTivBpmcVt+sWkSJViPaTLAWCfuw5GwlzN4jDkIRHJmyRaV6H
n7wtIoj/OJ4XN6c/x/I6Oefub49rcD3caZIB6Moq4YadZtcN7e8m6+Q1cxJKdjFIb0CSvvmqobDS
yEAWORoHWJ1tSAbIHzQ2e8NOZ1QFcvOSMB9QhK8ElFkFiWa6d7Lf0oeJXx+eTb3lDgxXdVeMxjrf
I1v8p6o6JWKR1HbqRvlpe/M0WUhRReoEF9B2PAsuwa436HZqLQA8/0DS4zjnhtyGG5Ma7tzKX6lK
yrFC7Ctya8jtM+WGva2xNqo/McQejw4BB1XdNB//HZqiwkuZqjFy8ygevA/mUuy/Ns+ybgYlFOuZ
nsNHHoiUA0NaW692DXjFG71o+wM6h2jCEyzAMSnudZ4y7YIqirY0ZCijfJOeXS8SP/Tbud4ApsYZ
uOn4RpG+aTMgsXPNQlzXwvieVPoFFmeQiBYdSfnyJc2pO3NLyMNTINqsUMIiNWIM8X/0j0hC9BhT
jYWTzYSbQ/41Mi/jE7/MStRQ+eQiLfCYFoBb7KdqeGaAKfd2iwkn2HT4iCaCPC46QHCvWcfsRv9y
Yv7qUJf3YjmMktFGrD38jqUdW+6OcM64bmq787YyVCsB+QSlbFZVD7w8mtN7WVjYxnCYo1Jxg1h8
kUNmsqLK684Ef1uiza8eRrm48VVFwbX+Vytl0MMdBmBNnFeMr/9Uzwg+YuwfhanOF9JVP2G/IlZt
tnshWsEWqVwFcMKt13FPriD5yN2pWYHbtwJgx1wNACueeUygsfbWxXgqFekYYDCBhST0lNFX3lTb
cVCczQxMVXW/k9O0WdUnkQNqN3mp8x2BgZO3ZPis4TxDrCuIQfs2YC3CcbLgVIY3kes9n/CAAMla
kv3Dgy70aMIM6bP40ij/1bPRIC1eAQBcOt02ScVFnNHhtySP2xvbjLKzsIq02DmIWQl4bNkambkr
Qjz4Ak/IYW6ZR5BYGa5UwYr0ZHp8+NE0Rco8OdaMCDWXtzcT5F183cmFEPEtU9ZECzCyZYAWnYF+
Yu9EhHh1RBIbrNWVEYBYmDDazXFcwIxlaPvZgpAcDTOFH2vRRfFEhWcxKSG0pnQeEUYTwnPRqBxR
or8X64X/BNfZP/sU5pGf/8sZWb/HMxxA/apGxtiky34ddmIybYHFCFsInzoUZHGKJUAHGdHjwK6Z
i5726gYiA2jPkBoJTwG+WMUkE+5e7o8LyfCTXuPFoSZCU/lFyqg9WgHxk2HjoF8p2chF+58HWYYc
hmVsCIueHnO1tWK7y7NYCLax6kR0KvMYuNUri8e0PApBN1hkIMi8wj0ZrLllQfycONByvaNSZXj4
pXFZlJY/HDkVO+bHeniF7Fv6k5OyEVeyJuXNWocwp8m4LUMnIB5FSeL3OhfMLl05SAvwn14KZjlg
ZGfXgItu66/0P0StCg5Tyf3GQGmzNEUBgnpukuRyTz83qc1xgPrgRA5W4M20b29OfDCKQmit0TaP
fcj5sroVBL9KW6MxKl1dH5e+FlCh0sDg0AlRiWWDJvnSpDB8o+3qb0MlUVq/pFqrmscX3WIKHGDt
J6AM0jDzBBnHe7BtfQcZS57axipXZzIGqGPvqjwaHpLI159XSYhZSoW55jO7pPutZJMIfAyXbx55
FNCKGYPQQIW2GnCZsA9GvaW3jMA7Go9zRWtgFogte7j2GXcOBPrN09VyzWK+3P8U/W+9saeCfc/p
92XjWoXSbZBJZFzHvIw0aNc4tdTPKKWLNvEdUcba+3n2wJn2VrbcLy51AlDg0bSF4U/GIyL98wj4
egqbBRnSVmk+iykJtK+zIfsQNDr2ViFdaC7LLYojBrGNEocZjY0QgPOHP1bv3Xcui/Zq+tcs7puA
aY8rnsjpgFkqewEaf9Mn8S0umEe4uMWjUdMuYiLXOt4GunFdCKmT2CPN4DR03TGwclBAa4ycNY9O
v+EOCH5jx65P/psyqhZjR6xKF/nL96vj7K51GGwAj5zuaoS1xesPPV2HXHgHGniyAFVo410ApTX+
h9hzSF5C7vQHYaf9Gtdz6/9Mb/+0VDHUimZlo4YrcwEQMcMJ52evj3qoB2PqplWNUDui+FaM718o
kLj72S/rsYGspjZcjX2naB4QkMCcA5XaHlIH7cGFm2EVWCv2GDm+w1SfqfpMzz/5GBpDMn9cob+m
e4Fa9stGzbMesN1D/lIYJ0ab+tgentew6bq2bWbdpojiCa9e9LXKY4eqeeBkMdUFztTJXW6nY2Wz
YXRCJaLEUnGymnYucAhXuc8rKTYcNGsR/DxXqDE7rvP5W6I0EnJHAOO6PmBRS06hIqsUeUiUoWRC
A+CSGQAFf5KFo7KK60pAQZsEnpP+4/lpxhMZ3BJ2bEcmkDz1ubfgsWuWHRW1J1zVFWoftzLJqYjz
7i5Gn4HXMxWFV2ixrwwhiNIm9d8Js/uuQ1y4KIFVC6wN+yEwSSWz4pBjaxGxFZZJ8ge1KP0SmpPz
Xiy5ZR4Cd3pq3JNoo3NL8q5seZ4yY8qwFt38riYhE96MnekPRMeFw97oWr+8xtWVd/11zKS3aN6R
JrdWS7SDLuskX3pql9fJq7olAtDLGZHQfjfLsK5BSVaDyRc5oqOCYpHsXKQDMYqybCWwZ9UNdtEC
eP9+EL1TlCBb5L91WZ5vLVq7O7c2OeFC5XplivAYwEHTSUdJSa0EQbtwH/QecGYMTxcnzZqBI6gN
QEefbBrUC6X/IRybiHGzuU0NOD0sWs0GsyHbNM30Hn3kmd+Almgf5X97/N6cksODSWz7R2b4JFo9
6hxKZQY++02vF+wKPLSNvH2F4X/yBEQACjnVvfdxo3usyfgi8ooJFpetruER5QkC9WmQ7wDM2/BY
mnmjUpGa857Mnc6BQELzuTgPpAvgfyxeivAsdnWCm8OWtavXUHBMCdvwGPRUcOOyKHIca/o8T2gG
Y07m47bPFtCXjjqVsJoFV5cDHPzJX8FJAF3jnPT+qX7d9bTj2ZLQ6+2aratY3zqeilf2UMAr9WZ+
7xnhihAR2Jd4Zla9RM1uQ+EwuQSsZ2IWxGp9QbabpVUjnPKN3DnNVSJgf4FcML7gJu3EsOVi5Vjx
YsTxvK5t/XcWa9SaYe2I7av+lm//PSJbXt3TtLw9YwZSNl+L0128fpF8KZeH0QwVlC/uGTW1X6ss
PqdhQsWCTxgkK7+4rvAhMZzDXere9s7F2qTZFjRnrH9aBZ8BTsoRxA6VB6L6YYuJs7/Xz9k5AZdu
2p1MgaveuT7RCFBTcfFc4ojPsQFJ+Wr8DldPGhM0YAyQAShDECEBEKy4XBqazgHYduPMTtOTOty6
uJhTHj70d3kzbMjmNOC4ca7sX2Kch79uhqBDG+gMW2xcDhqkrfZkKxRrV9YML9KiLy6MNdHE6glz
tnKIk6Xh1g940cacvkAnzgyM4PC6KUbWk+fMyp+6U6ThzsogZj6fD/hgwnXV88zRL+LTfoCrr1r8
gtHmFQ1C/c1GUdAQ8kecxwuncUcT2TIasxXcmdhcOV1l+Xh5Ynr3LG5U6Pq62g2RZKawGhvOgGk1
6Razhu2Mja5RjXcLS+PGYBofsbzvGWxWPSso87aPzQwVoh+qzVmRqYlbLNQMOLR62nZMdyEVuPao
kRJ4ILnFNhQ5awN+fKaDnSnFDl6rcMJHwOdzus4ylG+lWXH2I9GWJ7SzamzKAHxVQTg5d3q+HcMh
SanPXpEHn1T9JsAdGvzhPvSNT07l6JTUWMAdLI8DqY2hC+WbbLXbm54dG/q2cVpyOdOgeRdBtc0w
X8qnHKNnzRbkYNMhM61bNDkEDP4q19znNGf9dPeLqu1VN1Yn8ohGeW3dc58t/9rbZ2gwVnEbVXfJ
FSzqpBgDgiA+5tR1uduCJsk5/9F2rm1v2Wag9G8KGCE6N/FzOJQFvgd+XbjCKSA4weHGib9R6iAC
Hcx4RfvCCIJMgErEJy89MSITmeIVlE4YtfYuS2Cq1zdUb+4PMJH6/ZyYk/BNCkiPi+uXSiA7xsUQ
o5D5mPy+euOzBbIdDvbO9ODu0hNmHtqmq1mzRdCTjdJyUKgKTDNcFiymZ/2SCv6IyqhkNGJmAwBI
LwUSBoI4ht1xynDK6RJRrzpRYd+yHTGaeF2raSSXiq50MA5mTUGHfhjQbOSujL0wyLcvARLPI7Bt
roJdJ4YEIr8ppFD0z38n6L87iQP0MsGb9ki9g6ek7iL1rriBHU771xDQwmHZ4B0Z2IZHohI4BTWo
lRU36eRyN3kCMnL890VZwx5eADTXfZuCjDGgpNo8XhOLIdFVTHdOj6gDEsyf/+f16dr4TaK5TrL4
OP8UrC8wA5cq87pOXiqlNO0xf680xLNT4rryX4l9YdHE0ve43zjXK/EX/D7eNQphfQc8WuNy5PKX
Oja5psIN+JvKX1zrtNLH3jJeEPyFNS60qGw2LRVDzYjiEVajdNOMK/U8Ed7KxSrR8s1QHXuicLXx
OXtddzfvUr2yPbCTspJ12FgR8+BulQaFLtnHuOrEUc4aTHkVoxWQToLuDVNG8FSZXHqyuWckZZR9
xl966jjQDYTwbVa6xFAIns8S0fBH1c2VK4TRuNbXQKKqvIIBOSRKYrlkPfJoPsACqEe+6j7WR295
cW/0r+s8AR2aavTAbGZ9ToiovXi7tabiGPQxl4/SGpZCAhCCxGkBH3az37W7T9NWqbawPTn4pPM5
MRuhVbzYPGH6EdYUh8efxz6q60dFDNVGjlV1HBuz5GK7c3IN4yeQJ7IDgTHsaD/FLuRdfCwKlHT3
1LO8SYQ5Mq/qmLCHW9+Pg7WHfcb0pkJCN3pmw46bjnZJBhPD0cplGBMTwFATQ/aiXfZx9DeLED1D
isC0DE4s4H/6fOi04GE64jiw1xrJ+812jbqSsNmvwigoOSLavHQcxSNqs147+4zUSid8j03w3s5a
KUkGCztKLlC1aAnjM7qYFQ/2taU3u/ZXnxsAfgNEx28vYbtz4Fo7IUEqm2o1hCWy5o2AQRQeyMTg
QKhJhAbw2TGUMub9OZs5msbsR+cQf8rfRy5MzW92FwJ8+TvHJRzsFcFmA8F5Jv1IRP3ncoVnsoAQ
x/Lq7t8MP5GMk8j1R3GG2Hr6VeCpVCU8abplnQ1G/QA3C52jrPEQ7ExsveMlABf5pN2xo1dffxCW
8qVXAoEg0Ixlh7N+evdT8YnUeXWPiH/WWbQLkzRX/0xBxTr6FWNIVd3DbjB2/RH8Q8lojf0I0Qz8
KS9z9f2ktyt8lTylj6cFn23q5Ow1TMZeuPDpK7FOXrxpX+3nc1X1si4mM7r6Dtz8KOCx66V/pjA3
fNSLU6LoyGInvYnpDzFWpGRD3LiAzl+zUE+7Jf9SpLivXUnG1Pq+Aa7ylQVVl4saMtXQ2FmAL2TI
OC5Qk/xzRn7fptEN6Oje6h6oeohrqe/RKhkcsHaUXRmZSMA/9CFUyRTYO6vof3hLp86VhqCov1pW
uIkoIXSarixrEMsXr7R2Y5BM+aWIV1ptfucPATGnc6frM5MtsVcFpb18uD7D8/gwyEvzBrMxxfjf
myYSazNBX3Vll8vwd7zWqhe3moOzXNCrd2nOcTFImfY4s6mcyQm5RAjAiSM1GlGwb9Sjko8WsHe5
rNTbbhQH6vmTj8FM4haWZAC/jb2kPVaUlM+v5qcXMeIj9izhHKc6asQS0F5nCgjOYWTBIWPCPBbI
8PSUUyP4rnjpc+LCQyOy5Dw4v5PcTwIQ9V0c0K5bQyBgC3OkxFMIoKBMBKxQ656w3b89vkZtMWJe
FYu9bTlloq0brQ13uh9NaXcf1pKs+Zo2PxFRVQa+Qmb20CuRYfD1jlxE8YwoVIxtUU3F7U7eap+4
MQAetphGjxdx81XB6SQqfiQY2DAk3uVyyNO6ZlDDWtTyXQJC08IGRsX33bvpQ//Ti19GyFImJF/D
D5YSWH9FD0kPvZVYmx18npv2BlVH6f6+fvHn6m6B1aCtjA+OFuOCyEv8DgGv5Mi7IDFOM4YyseN/
RQaHrfrx4PL3A8Q/2DZM90lNMBKxqLRvxckTQzIloR6ysS7TnowlkoXNXLxAFBEGnGNZ/4k3IxY9
3xvngNXO3sKeTpWBoOM+5+A7rO1mMJFH1iRkgHQ8q45z4H4yggaOx2Izy3714SJRe/cpiazE4MuY
kC1UDkX4zBsNmM1PTYL9UhzbzIY/0nfFjECM5vJ2XENhlpY2pUNwDVmbMb0333zOfM06p44Ica+/
eVTeW38OfEOn8xOAO2urQDrCV/+pMi9RLDT2vn6yz/GN13R9weOLRuFT51ilREJwmDP60nYZg1jM
7unT0vLPeMYVzK9m66NvtcPtJKYzcTDzcLZ0lkC/BTqgZLDspnyOvc5fH7szcit/nnjfgtC/oenF
X54WAxP8kK/g31qW1EEpLH6u3guTSVTvSyk6OW03X2+q+fWL1vgjEgvMFg10qZCzNb4ock3HooSz
swli6AdlzceyJ15Qj4gCCK289+NdxkPPdjNkoJolt5OBAGwm0vKP6d2ftY+gBmNoQ50d81A4AtOl
qTjfus0Sdfog8Hw4uVrmkJwb9V6KpWaKb9fTK60Yo0w5n7MlVE5KDaMz32rDjBpSTKeTkkK2Hg8A
opX/SI4Yea+v6mKJYJdh33Ahtkxsoyr3pPwf9cukTF2594JQ0yzNv4Nj8P+ujRUL7zdNC7rYXQxC
RUV/T+nQjjYIKzlOdPhODsZhBNWLAjTF1qjAcoUGmnNRHu1G2o8EQvncbjJtglfAlwMjkICWi/Pb
RUDtznS0QR6sCJZ4GWKeY4IUErvfnXPaKLkrHpQcGYNpLqO2yCZMbEbf+bHP8/UHWSfBW1PWGELW
Axqzxv8tH0m6pp1Lb+4hwgeWLZ7TdrrmI2tKB6yLmELtzImUcP7BvnaMmNg7UrokuNQTGTgkTEYg
gTbqWIsEerDH3dnjKvbQQTei1LMEee1UTmvyaObu6A1MAs2Rp+/AzSILYeW14HtrOayAAXpfr0kh
a8vX51TWUH7EhGqkz+0mO/5epY9oxvx60Ievytt9HFcXqsrHDJ4y1RLIm6xcVmbjkaLHZB6CEw0o
qcUOPG3lmrpm9sbfmySjrXrwAbMBXyJUTaOyNAu6rPoJHjRbdFayjmfiwZsXmDOcKmrKjNxzw9vI
SsHvisVj/PYf3Irojry9rUb28gqz9oMJeumwsMIGAwksKjy04rVZqo8UlCx/3hiGPFaCzt2lxRag
mREGyoOmS7kDmGvuuIbP4H0TMaXtIKHterzkSGj46hHqUEjvFtHszHV20zNcg226+ZMRdlltWvu7
N6MvTAn1p4lTa3/+ClZQm8RJuihPjU9E8tYdyCTYvCOyZUgrJPFmMYpWktjlpf2WNY+qIveTXIVc
VT4rA3jVuKiA9hMInHZSXyQGKLLRRVfiK2wOqB0+FH2RPgcvewZnIDsn5S2hi2KZNvgc1T7N1sRl
1pDkvNz+JLvNYnMGvUdk08LoO/MSPNn0fN4ODnKZL7fDkx5uNsEhc04uJnVnAStlwlJUcwbNVLfl
lbkbhVgfOPBEd52SMsJoKPP+Rk08jwZSYqIyGSZN+TfLxjwJ3rSv8yBoHrejzk/nwX18UZ2HVv3E
3RsBGPMdD9RTOPgniFcF4mvVaZSD5Hv2D4QOzLsCkUgSfwWRq0lbDV8xxzuWcSeObPSnLtqTYouT
aINCoYfSdl+Odg1xGeJHMmWxP6f1M+w5pgS+ZvUOjLyHxj2jRNbXB6eztIyqzTE/bO5uLWePHZ6L
A5SEUnT+pC+YtcfUSLXJWJ/Epg9yEpyeTqJqd6iH6Ivx6GwXe4kZXwV33fgcsjbQdt6awlja/HEb
UrxAPyOvAvTb9DqQzYyOoFIksEAmuhFTTZs6ViD525ulKOoZN8gHlh9E2jzzf4BRmywNsZ3JmlGq
MIHWD8EjY5c0xYJpWN/Vz8hiAni6QkXYMpScNdjYct1yqPrdYtxGU+nU2AQjO+VaFcQCdX1ap16U
HO802/dqOOgNUOmb09JXfiHvoQ15Egn7E99Ijuc6emW8SB1VEwnGC6JAe0N1RCnAwmU+EOj2pRE8
3mDZTJDAKm9qJdpQ030fAk7f56YOrRp8c+U7VSe4PjdcM6k4JoMJ9mbihlNT2oU59EVrl/xAOznR
exnfeNo36iewPr9EuHRjAyJ0yFjVL7CeFUaj3LyCD7V9sdts3mihYXCycbpgCIi5Mi+jUqECzQsd
LAwDq1u2/vEgCqCQk6JFl5Nxato7GVY0qhVH94ryiB7ygKwlwhLIWhoxDG4HXcEXE3VKdaAMfNVi
prBS5mQPeaLJT0pb20eW4Y9EHnZ9V9n41bZduILBwOm9jS1aBdItJfnJGYtr59Q+qgybt1RSlRMQ
GVHCKNf4idgPGWuxAP9vkNC3+Ci2KJ5ifb/3pa3NiwoxHtDHNGLJtCdNA22XoRuveB81Rj8Jt/lT
KUE6276WOefzpksyiAhfkb+raUUxH/0hF84WRtBiL2kiXThNWZK6I+XnHL8DYvC5N2urAffJ93vI
FmiRLthd6WzcKpZB4oTDzGZfF+yZ7dqt2p+EsZIdfxtNzIoqQ2L8BU4xaYdBEj7kWLiehyTJ98Hv
M6HuGpneZdkXOhjfak2LntjcvuRV42ExioeOHjPJ0XWTo4OgcC0ATfwgmy7BzCFC/UVJLu+OCow5
OUYEgksYo8tZ4Ji+tzpjB0pDvdO0XdrV2soVkZVy0KNKCvRviYvka9qvYWEmz1foMzeRc6vHp9PJ
GsFywLr+ETyDNt+dCehu0AKs7qZhLQ9AQ1o4ojSMAWxahmq7wUgwyCcjiXewAIfMxxUtBU8nvuh5
zwB1atdOSL0BlZ7LepKmYsjzRHsbcjFevPL3Sta0RkWw1HNpfI4Je6JNV+v6UZkU313RwYpm4HKC
V4C+uXa7Kz859GauMKZjQDwC8INYnEGXeVhxSSFad+0/bklny5ISYKDhH/tk9QOIVqThnMNGovX7
d94JyaAFP1fOMUz0bMfwe05IJUTG53KjMdM+znJaWgYbb5br8g4PMA2yWAnqS8CFQUDXuxPJ/wQL
W9784gOfecXJ7yyhh0u+4tWQRUdHnn+CNGYjzd2akzjP7SFL3993wBQ3O+d2DZWjjmNZtSgyWh6m
fMNHe4Ur/O9MHLVA+Muq2Y6cmeapOzpXhq3hl93JQddHCnqn+/cNuLnW7XvGDRdLq123pbw4Vvdl
BMigdNUBZD5zRqSpxrcPB7W22CgyYGjlf8TpFk/gPdabG0sDCRwFmj6e+gEfRPQX2ux7ON3lXpBW
8xtgkzLruBOZOFbGYVhusuYwA2f/8EVJTjAlJ+mCW7g7HNj+Dh8ICryopUEmxzH18Qq9TgqHJb5C
DpbB5zgAgOfVuRhUT9sAQj7pWAJTy8L+7H5RKyeOhybyKoJpj8iAnlECzqLQmIdO0b48WLLfqTJy
PmNSCJORd/b1zU2nib26Nac0Og4WJ66o6v0kHlZ24NKQKIcPInoy4pYr9Wx3LRHlNzhb1p0NOQkv
USRNbW+sHUmRazW9/t/oTWThuECyvuG+p04bcGgqQq96Fqgv96TmsjH+NmxSEFkGJfQ2rdrCp+Bd
fpgcMoLYjolqmX7qWCkBb4SvDAJs77jHtZvE84RIZILkni1+Ta57x6H0SDorolVMfk3Go3t6YD1k
K6DKTaxUqUCRJqso7Ufi4Ul02q7lwVWC+OpjNd9k6zp/hD4qHvwl2IaTj6XbP3zMReFwkD2hVK1u
XLp7RkVHSFYFc232ubfvKa55c7GSFQlONQDb99WNWSCq2cIzOPlXW+9y7uX98ZqbNVwxtd9OdbmA
s/3I25qO7BumlSqq9mPfpKvUqv/5VrdsSY7IOqYexKI14lonVKssZviTnEeu9jpDzo773nAOYLr7
DR0vj0QASC/8fPrgSObldRd/ZXIJlURsYkpXZqaa57+H59vtCSbhc66KKp2B29iwn8Y/TxU3pPrH
TUAsqsrBs8CjigVpxBIh7fJu1htaQxbIQoVpSKvSnYSiDYkA8eupLpBjOLmh6v/EvLT/0JNMTfA4
0tjb/kCepqFRqh0T6MVi/nmDqqnLb3IhTOVrgPYaYJoe7RiTvdpNI9Gy7961j3ipdWJNPu9kMLlT
B3Slc9tyDnXmbQ8aSJgXfByVcOs79hOygkBlxrX0nzuCAEjF0KsseKTqpr1tCOMsdxeinY/NUSWP
R7J4JaZZPqYWwCLxrkqaByk7URFWHc4/SKs754XKo+JLH6LPPQChTEU22BnIr9zogV1DHT8tASNi
T8aVSFSdZvXUZBiftnkcM6mYk0LaHy843FI4GGP8QJzYWNugbiJTtCK9AkgOhMCpCEp6ndX5CZar
53DyJntdsekbfy8GS7SOXcau+4KyIxpYxKfN2rVJ35u0d+4p+h6VtFbbzmPPpXd3vbw4KSwRcyyY
rOr9OOeYCoENL0SCW8xRFrZ1GVoLbm3n5/DxboE/X7qeYnfdrZaZTk4bjZRFp0cnO+OOiHHC8foJ
R2gaYHdYUPd2lG+cgFBgHGcmWfns6qKH/wK9wYzWQdwH8Vl665IODrGywW5nfJ4oaB5U+dxfoUPW
49F8s0NgHjvTpoRbOYK7wrPzo328gvQ9zCKMeWZSYGC02g2lD89DmRisoljgnLSbG+Kg3NtphDs4
JiJcOaWFnIVcz6A/4DODStSpeHUdLVbQED/+cYN1DUVeCm7LPA0Ah5ZIILhctRgYfJyuIekh4On5
HXGLrGenPKR74ErQvsgLzdKvTUINNlQ+4iRDRfXB39+6rhr28CLYbNNcf/15W8M5hjuqMClCD64T
Wm3MaDf2ufcwEp9qOBKd1f51t+RQNAIlknx5Zb137ii/wAqb+6VUUAUwQGrIsf2fwyujqjI/XKyx
FqUxyP864UjXzYY9+aKg59ybgxub7V/rPAgnNeaeY4Hwr5Ll5LxZW5CnOmnMul1bDT/Sh5vaHPj5
TUT1wMcic4eB6wqjUX/gVT8xuSNjufphq4ONtSp5CfvVmByooP4iW80RZEkQw+uMa7KvaewXWRYJ
QTOqzjbcHCges9EUmvCdYkJwYmDyE+OU23Bv3Uvx1O/2pAn9A/caVrFUti8IYdKHP9Fkj1Hm2g4D
gIVPE9kuhhkdwZg86ZfaT5EXVVwIV1/Nlpx2zK0yYSmdSX8tzajOF0PWmAM0APmzQkbBKbv8BKJJ
Aij/ncs25KG0HjJEE1RgQFRqwl7nO/evJfQ+nOOYea3Ng+9oFqZaaEDlYe0QQKpDlrppfqaYTgZB
h6d4+26IGf3CPfV7NTKweN/XwrsZS/8MtaXm+UT+hqQqXIkYxNdpiPeniFFz4+8qDgjpjzQfudsO
jg68WHxfr/VDyRGYIS0gK3H+rVPaLVIdRKjuPjJFiqPsWAIa7FL8PltyCEHWvGiq7sYMHXugL++Q
QcX73EIcC7EKHX8rLtKVgmqlTGm1LO+JnniKOqDqpCGF7y49Wb2n3ZcHZ6vWjf4t4XniAKpEaGiH
2ETRQ/gSgvmwA+Ph0qNWIYmybXy4n6q+DdtUr5ydA/rN1HRXMQUe4gIgSl2dBgn4vkQHSQDzlfJW
7KNOqFOTUxKNnJhUAQb1kRfaQXlgw2B3mayulbMbF4CQJqvLUztLIYSnQBqTPZQTX9U77X9oK60W
PIsmQEqtEIrF1XfZSPbkpolkR9JI+YHeM93DXkA9QT0K4yUCtx0HfwwlxRoTYW/sV14t+XXF/PPq
yEg4eGiMpPK4fxdeWguDGCen3hgm5in6YRyGIE8gxxP8bKcAWn57yGt1Ov2k3+f89fto333OtT4O
ZNcgQgFLk8HLoArjm5nBXNmLxRn2VN+qUyhdNHGKCu91TKMWjraSVv7+xDCUu8cPYQ82HKrqFnJ+
dNl2JSuJFCdPqtAtJoWZLblvZ2pHt3B3SS6y2wsO11XTKIX273SUcbHNl3kFrGh6uO/g6S10dfy2
FQ7eLmVUPB2yeEWjXxFSy9lZi/p7YIMpRRg9J9gR3HRxHm4vJeo/oQUibf5JMxsXnuRyzJ6txeRX
IjflmnqcEqfVDN5B8pxx4tjZF7Muyzgk6aKub/Wh3aAkbckhAZPiJiBU6Pg2FZ6puAKTYNxM888N
RuB+nlxBkgkn9fV0GynfWflozSU3wVXrolC20hU58FDxT9+5Yc63TwLkNd4pF+7255OGwNVeMH6w
x4HcT2sj5jcOdwuasXVKw/5v6PGV1PEEAVa9pHFu/WYTFD+4L2Pzh8jHp9znPfwU1FemHoIT2hPW
+gZhV3pgoO3DBgC28SpvQ3xjjKknLf9firbcfGLjrisoryOEHyMfIgw8U+woI4g9K6Ob+8b4mq3n
WUpA1+qkRAHpDJjxFwz7jSzu/ZwsnsiGCFpExnW34vnvLRU+RpCEsGdkvawoxmBHLd93afjd6Cx3
lU7ZL5IPDdL5yyrlxAzFBXQ8mnJ0/poShAEv3KuKMy0hQZHJABJGVWQRPC0XTdjW4BbDslXhVC7G
Xf+Ol/KOenB72Hg5faN59wMtbGFAYePOTBw/MzDSlRXczk1h5e6wqY9cci+6lzz7w8bO67Bj8wXS
nz39cA66pUB6oJ/Wis/GNxQ4lajJDqY2DVCpkHl1x03CM/u0r1jejMWGIr1eOErvaDzO2xehr53e
UB8zK4GHuYftRTng7IZd9B3GTgbV5jIPORfMBx0suQBDyzhfXyHE1X0b3ikP1ZoAcr6/vCwPdkWT
FzRc4kSM/Zid3Oz30GiAX+ek8dAAvS/63J6O/WA+FoSpWx9w5NFvBW4PVO7TEeGHE4kGRCZp8g7r
22b8hoTP+qoQeYvz9LhBZkU1/l5/KsyC1GPnNLDgjTAnNiwkYb4kC3XFDqRaa3j2TU2BBNw+gyny
IMOan4Pai7sDjs4/FalCSOMCDWrPBMWXpKMIR08JoMS41hozGvOd1F6Kb+aqHauvYL5BOwM6NQ/Q
54JGU3bfiIWC0veW6ClwKrQvnzfMX93NPB/bMtMzPThjYmdEPVIVX42ciApDY6+jjTwD3gTTtNQ+
cDoU066TqMsbXT/P2tAQFWbHJVaIQJsPa9Pr0mfQr9XKuidM8fn8+BrDGtRw0I2ZcSOew44U4fMy
zVe84jeGAskykz9OqEFOHUxevaAfkBnLSfhTg6nC/FEa+i/UUZZNN6yvvCRJBSSwrUdZQy0wx4MG
TAngD/ecBKdH4FU9XhbTkxeWSkOO6YbCHV07jMOcxAS1lEAJuHf14WNK/nIB3T7LyFHjFA0WgNb+
hrMN63zmvUq7c1b7Bgbatv1MMSBWLbbDAKwWq4IuBk7GFmjmx0/6D0TAwna5ILe2K+Hqwt8zCgUC
B1dht+AVZCLzlw/XPSqzpSZQoxB3GQIC9SgaSvChnX86cK2Npe9HrGtkyiJkxzbOGvJcaLHxme2c
AnJa0UaA+fcifc2DLzvitoag2yri+O9WxZMy3t5xdIY3nCulGDiakTOju/3Y4c1Jj6Gdsf63A4Mm
28B5sFSURf7tlRJ+KJiJ+pnHWbqcdLCCB6RfYKyVnQQ+byM/XDaNvFE+kTRcT5fk3uAUI/goPNXl
MLOKoWvo0xtZ5I+1t8dkIPIO/p3sgSkOUpVFCJUC7jyPtfYMLgOUUxGRPaOR4Kdg58syOgbarpac
xEmgGVf0dp3XDM+2zYlPQ5Y+Im57943sAKVsalpw7+kMug0EVyIM6zPCXdAWUd/GBZO4IenoQ8sF
PsA4/o7ALrBy8wnq7HDw+ujxq2Xm/a3wQSrayzYu8dYsGi7fj9TiP5ranGhupGqpa7u2pJ0bbxSm
QintYYJ2B/jzJDWW4rNOjVt20mb7IBuklhLMBF6vkog22/ns/J9ecYrYuFkVbpMU8rOQHWi+J+9f
UiluMyWc8E1VX5S+DhB5FT0gw2fPuX9Dt6/OZ/uNeWATcqVMt56i1vANXOVFm2HFDBkA8r5OgXL/
17L1aM1uOmGHjjVqL5gjBApfqJJ+fOYmODJK3TvWAT7Kf/AzVC1QxZHenXoeKZo3u8dPi4o5dpZt
AcQf8FseXmnXBIqLNXOS3nTnbC68v9/Wk34lSsOzLOWdDhuKixVxTojxiRD70iZXHT4E4nOaJpB+
9rP/DkHEbtaUJg3AhkEPZTzkAnUGhWTrOls/adzXdmESG4nDYcWuju1Um2SSUsF7P5QZ3//WZ5PY
ubdJWlDCAOtICibBsYxLA2WmqUUANxSd+taXtgS3mvF/A4oVIRIdHoHatXSTj26L14SEnw3S9Q1t
8Lg/1U+hRwQOA5xYAVpSlQNpbXKgqeABKB6QcqKOAppZHbwXwwnFLJF/XrMgEtVK/T5h8wY9a+p3
nVm7Rma2fbRD8MezwOT3GsikClTMSITx8YFu+nXH2mBBmFNeuJAw+QpCstBetC6BuX8lF3679HLW
Yby9nSFWBYLN299sGPdhlzOtZ3s+NzxZ0mdIL8zCujv5MWjSR/TGsmqQrn9QrgD4k4V5A1ekZ/Wc
jjFM2qVk5QA2YnX7wzPK73YOX3InqdY5rx67fsyTifmlPeHDYZKpy7WNn8ywzCeQ3EJemeWu+sv4
64ZxkyM/Ai8e/Gat6Ufc9G+LTBeoFOBsXxD2im6dqNGXW55ABfFt4pLgzdaauZscqezhtFAjaFjs
66tsGxH9UXfbC9iLw9nx6xphvBl/OlYHq4LR64KOeFYszuDcmSIrQ2lCJKgQ/d1VgZUoC+uBS0Fp
64W7PUFQjr+TiKlH7VfAli0AqBrqIq3fapvysi482TkTvVGLhhHCzWBzMVDGu2zX1yuWHYfYbACk
5S0mNmQyN61SQeXkqWOutY/tWiCSrZqqn0em7IsLPv4d8jfH6Gny7i5w9C2ulTdPkQfqpXbKEg0n
mWjWjFQTZXHBNcDRToQDHo7ZeRU2ss40L55Bmp/TeA6rJaCh2LeMCOwiqj1kkt6jPphUzm0kj0R7
Ioi5Pakpr19/Gt7r26tjIN49+ZyP8s0RYBvlFXfRFJzwaNXRJgzTlIX8UiosK7x9mJ0VuyTi3T6g
GgN2bc0DhnlBVusNlTz6VqRTCFijJG3jO8mfNod51qSZfWBcoIXNQUkyQaVDCIut3SoRFkVWQZnk
Pk3pCc2Je/8mtigXPUX5EocK+jhGVdzD4uKL7hsFSAttnggWE8e/SbLdKeC7+gHzaQstjzVJGjsv
rEmb73XwzVqK6nc5X6qDgPpxpaqlcjlva3TpHSED75pc0Ndcq71Z4b5yTA2F4gE15MDV0W6iPFmT
VmClcjnOz9Sc8j09Nxex69//K2Ju+QIpAz6WDfBAZaPtOXwttn5dhUw9QN65SsNXZaM+hCIERyuT
QjoFB+GnOAK2PNoCjTCpAIXeBIY/iXTq0miz8txv2Z5nkG4WJqrEBVhNtWOSWQ9P5n8lKBluA7p9
SMzwd9hF5wFMgWnN31qe1/MVG9UKPsyVtBHn9hmEOq6cU68gaM4/LHLl5Q908o9acv2mzI9OEqow
6dUhNDLF9+iboZdkPQEfZEpl12NYKo9bBvslYPvuMkdCxKs4fYWoa49HC7pMZLfuQBLWvZef9sYh
+oWNRdPsXQKE7bZErfbIi7ShYFQAgMI2ldtyuY7tzhNHG3LOgV1Icme3KNaZILXfBDDc5Q4NGCEP
BIdyZNLvtFxEKu7EMzuULmuaLpcEbzjBJlsnhVBTnahw+ZyXP8JxPBE2c2yFyDSRIP/XqopOHwVC
CTTv+d6AupKNIBTB62GL0t+XwvXJ+gQvB/2HV//Az75E+GCKsSu6X+G4xKwzzbJdCIjmYnN9Wmg+
kRZIP6JTB+eIvhzxxwQUc0jxQRkSmed87nvyWBEXTfpC271aBPHIWKZyVzsQOREBYLwm2GnSapei
YU1ahJBJKZIdlWfCnWqXw/YUw5crOF/18Ww24M34BqPfiyPYf32PO2pGDCDyOsetXDKJsgzkdUGT
GWgzcaThf/LGrk/bO4Kz9RljLe08dpvNcOXevRFtKKFCIwQUjfmpi/7UzL+RrnVgUwn/sz+zWF48
AI3Mm2i8r8+I2XrKl+BkZgy0ep0IBXivbQrpreuCUvw/F82Ih++hRTeA347yXGYqjjda8jz629F0
dLI9ao8+clNo1C2gdMWGEVezckk0nu4TeaPGva/QeTxxAWgBorMXBsgp1d1M8WOaLzmuWZ2prR4D
r3cIwOuG3p9Xd+Ti4qQgA2JIakv/Eh3H5oF3KfQIbBjN67I5+KuIK6gp5Qg+oWpoJYjJ4E6NHS0f
TRgcAqFDw1z/g2OejzUgFxPSJNwXqnRHzLe3h886C0abLuSfkVBV0nItSuhBp4jxxAsJYXEVCgGI
MAn831McSFvzX73gMnUF8iFXWgOiQ7LTLQ+5bQ05OdEtUWaozanbyX/gDt6lwb58tKfgeFq4F5N1
2K3+1cVy/UNzwMgDXeQUMQjkezk9+izf8uscySyQyNapnOEJkbDVg21YDen8lR2DgUhdgoDnPSbp
edtFcKKUl3Ea6NQm30lovTz2bLTEtRJYsbPaC+QbvUjlgeoFrWIho4mQ8sHiY8YQxIeblUxnM4Ep
FffYxEwYFOm230Qs1HbG4M6G4LA4aj9BVQkTzsBb/xq6ShOl/dSMRPHSEzeWwSPd+sMDFYVoj/xV
A+ClHKcVeJEdqywc3bJrgYUYcM0ragkHuimkJgrkeCD6IfI5o2nolLHQrge91juZ1ZM3qZEyqL69
iDfXQTaE+tv2zlmMqW9NLhnUF9S9qQFIQ4xx8DdKetWczvBbwqGAD2N5/eksj+3IdzPk5Hbbg+ia
YlXlCt3rLzzeXCtodVlszq5+nqV2+3lpL1K8VmhM9Ochj1dxFphJC7EkrNzU6JQ5+zzGOeLMwp+v
tAGTvEcQjJ2OTPoZc50qZnguvCFkjQPh7jJeIZSepmu1/sDjmMU/BDga8KG9aua2n5wlQv3VF+sN
FC2N4AJAvE45D1F7xiq1SA/ai1PqDCg0MEK2191h/VeOeXlUA69lyAVIMPFNNnHzEYAL6jOIbAhK
UofyLWWfzqQzpUnexxGuFUbWiX2LQseaWMF3KQbVuWmFrn36BbnwyvE5wdjwG2CrpIWv3Xo2z68A
1gjNDHZAqXIXtls8krWzJriuf7zEndHXeRXhzHOB5uUAaER+o3qP1CDn7/wTRdkdxxHeVaa58Iiy
A3cd4UlhmfwI/3+x8qsnEguDGYMTJ9M6CEFaEeksSLHmCM02w4ptgQU4Q9wUzHLCd7V3MkHiryZM
b98bvdqaajrTuDBG8ZRlVhZDGxnOFXyhA4P1Tmy6K/mH6nWpp/z386XdLGNxjEWUzW2bgDFA5zU1
z3XE2G9X/EFdIxd6OVxWqFwoa5sBYs8ELI8XpXU72Lpe5PoW4u5Gl6eTNvIo0YDNQuvvmCYhNy9A
8q0h4L4scBRLMt5ACKQHX3A2KTxlQw/2NpFpbPDDTmK4OIBP7MrPFnf11fExkXm2R5t50oNbXJar
Fo2dT3eHqwRfxKYIdKb8b/6j2YboPYYmA4Um/8DQpHSBvBldxKT6DWViK8V8uxFQMDq27BR0Bv0p
yc1f6+5WRp5pASe6pX6W3GWdYL1rMEx4+RfFT+Lk+wf4x5avtntmfw7c8naOtv2ZmpM3Ooy8CExY
jaE+yJOeJFO9FJqwmy207CgqzFbgTinRy9gNAqY9oxxVJ5sRT3uWWWIU02uojJp5IYOeI65Ye9Wh
UMLkruSQxYaXG/7HFLuErs9i1D/NtwNJWSqlPJMkpPXLf6WgMAfp3vn7qEes3/wGFYJL4ROchFAt
2gloGk2OjKHZb5wkfWXaaY42gOo3Oqta0vVCKdYevaHUI7lmYaCVFwCsvoU3F21OG/mDWZJX+8LA
z7yPkgY0Ed3c3sKX7T4XhwvSaJQZkcgnmNTM2T8ze6kstkkaqh45xe8yIARxqHWh7C7MhLJ6h6cm
S8zSuPxfhiCX+N8cuoFQ1ZuyMT/nEwQXbkeBDONRucQq33H8YYRgpPzQwHZ/o//jms5zb2o1lLxq
cecEplsaEnH0lV9awQz5E+LV1bL+Pwfv3lG09lta5l3pDyNJTnJtrejDGsuIVSo64sqDtEhwj2bg
9MiW4da8TYE865yuzeZwU5k6V4w0VumGqDQqMhbIX5Huwai8568kqGKjewvWN+o+PAWS+sLEV7Eh
n7VFCo3lO2jxOIMZJw/u5vPrwikscmB1jzHfD8utiqEwP7QipgXOEJVdVaEkCtO5cikiZK5OLkyK
YX4t1VcSNJcp/HZrw2QCDsC+ENQb8QVRHWmpZfTZvznjhaqeLTCR0aPVvezpLkS/uQLBKGHKKlLe
zAvuF8iDG9o3dhbrvigCdY/ai90CI7/8Nqo1CQVdJx15/dm21h2pWAVdeat3PDTBKERtmtV/DO5P
4tGPtMK/5iYkxBITM6VgsvEevjbaYrQCkShU51g4Z4ggEhNwHCsr/wadFSXQOZZe9dH5khb7sVEn
AFGOccblZXYDGY3f3YErWJCPODSwrc2MsYKyMdfEw/C9SVrPVgOXoaB5a/hUx+RAqNj01ZqIUev0
rPaRdu24bA4oNJAjRWlriqLGOS+sbEQ597bipmTx7OmTEO8/67k7pYsKXdErmpM5s8CHoXoVvs2b
w/e+FXq6j8zNXGhLGU/nPH1DvFB+j+s2auNP+IBZtHxCvIqxaSzYvAEFWd59Py/RjPSCniVx8b0b
SZaCTM+0kdnpZ28r9j9DpwIdBNf9so2820PaGX6kHTijkyGy+MvL0BRQTJ1Mw8xAMIN869EMjxky
mgT9wtaiYpZOkbPXHe3vuU2IAEJUhm737z6PfLgYQXNPXA4R5xBzw/ovmjsniLryWpatnTfBrn/K
ia5FrNdadrDZfPyz/63dbGsg0RW6CPtTEsgYKWp8M/QrPVOYVUuTETgkRSvd/sPmaPqXp8tKT4nQ
uNmqLuGqLYlO3Bm8mAexwT5Lx8k2pU6jBrd0w5vLBnLwcDl6f37z01Ug1YiaVduTObIpR9VVaBbC
1HEw9m2oaJS02Ikcc4JPi9hKNPrU4eK/c8qEbdQFXhIUpqqhQYMpWHkPS8zBAl8ILyHRhZWM/O+V
vBTuy/n+eeHmtV7/2SAdBR/Hz9Gs8YJwHtD+0sKZPtCab7bz9f7DNlN4jM2v9BrGmGb33Wsic/CO
NwhaA7HcfOCp/gLjaP2BQkbdRYJHAgvn2FOaSp8fHI+ASLY/z/GHOeY18HfKb14lmlipAjSpD3ug
w2ri6SE0cow81uiCh3pdTp2VhV5Fdw/3LtC+zcCaIeLn7x4Wg6KVkHh3qck3w3Sd5xU5cLBt4QOl
gVUNTsGgkk+cDSZRbRNH4g+42NuM0vHirnW1znCRL8WTt8iL7mIhQZd/MtH+p4shxNtqVQue1+jl
hAbyN+Ag40QcVx3qUIJEt+LMpuJakUZzgLhS9D1+19WxiKu6bYPtcq3KiX29eyGDhmhgpfumrU2g
8qljTBiIVJsz2QEkVPI05j1PXHyDs8Ae3vTbe5BwGqSku7xkot6GJ5Kee7Zme+xdAOBzoxJYt6w6
x4XV4ZQyq3ENG9MdVeUoLdPLJMW/qbaAi1lt6IttKNfkKVkHoR5cVGD9AdolgJCYVJl0w2vCf7TW
HcHrYO6r56rjh6AZW78IDNLoKpC3ffGsnfCOxAjA3+M3v0s6b0lX7Hvnjy1GK0hbQeQqoMmMrS+W
BVn8O00Kc3yvcL1rvNCwsqKvaBvNuDkYMwZCwkIqkurAkfX8X9VbXHkkwKEEhrEP8pAmWCVNJzGD
3/qpib5OGvr7DxfNLIuJYInK8/eGtYTxuI6pdK/jmgMt1118aaNfMfWdsS6mnEr6O+ohTCSspnvQ
xzoreT5L8mRRCTTo+9N0/eCM5pMs3pfx2J6oS5Tj288aoDzb3qIlNYvN0n37ZVo8xT6piyC1XJV5
VgppoNdpb80o9pPxjJB1VFmwh/aLyoXxIiSCcgWhVbxF330InuTzSxYjgJRm81C0h0kQBaJ+DS6k
bFYeKTdJCB3wfakTHHJST1T7WQr4/TEQC5kaLpxeVIgg0603pxa3WIENoZNXYZJKMWanA6j1ZYoa
yTH8l9R8zfH5LyT4pJSevdH12dm7CKYQZRLSU1HEFa3X6G33bJSW267+Wd4ODRH3BiYL0SoQJVdm
1glvqTUHYR9PMDj6LxK5t+Oj0c4JztupbjFwBhNxhWE3LujBEs7zJdRINJajVeOP8YQVJ7+2Pckz
0VoMui/VVvMMZPHxdaLWnh8hPvvucyl8MbEPOb7iWrp1k0frYcH1NeARul4jsEG5/yApW/o5Ncc0
3QKIY78LRXp4xJnjor4ZVcCzSUNRCAsvDJ3Lt48YZes8gjrGb5sc3bE5dTqtTzXKRTG+jxYOXnZu
WrUudkCmrXKeyxhA8wsURSkig8jY0xs45jI8UAboU7DMduDTahrHoVIhVFdPWxVxsqhOZ/BrZd1h
UZnEP2Q8xFCyK/G1OtdCXshxKOltlvX65PgsOl8qPAuu+ZBMmcEU8BEp9o/cZYF8EzQzPWQ0maxm
P+RFMgKK5x+bCt52U1RQYmzn7S9D7D7LxdS8NTnrQdnZgqv/3sySl311XHyCYB+r1Q1Ay6I82CMd
UTcE43JUGQT9Io+aBPaGkgDEg4RLBo4G+u6NpoNj+x1U6Wjh/09XqQkWLr2QZFr+XyX96TTzimVy
ysy9XQeTUUUJN6VaE4vQRebEnT/NVvN8BE9sHZp6Z2e9kRtS49hiAaclVd2DQ4i1ifarCRhkhn5E
j42b8yGsFI2RdM/45jvqzkQOqABkCacUscYrCfCbgNzoL+sWcEbhCLG9gU1FgLB9lUIACKhR+pQZ
xZyyZZxIIcdjwrmtwlEsTfWabhOGVrf1TB/gRtJbGuCi9kRa3q2fvjVbSqEm5OdZcezGg6jENvVL
/GbeshgHZGVKhIr/OPn1WMiIoEoZGR3eb28WRhhVvt0YETqNiznidDOu4UD93fSViNwoSoondsyg
dRO2BTg9d4V9/vU6paPWeLcK95uaqkgdHc0j7wl8L9KZLo/AEtoOp8sC4AQSNu/MjUTJDY15shny
gDSibsUN0Wzbm/rwwCzAvimnhtfXoV4NDbOf/RmwZDtND9OW2vIExnU8EyNtbdBqzygA5aQgIbUP
ZeHQPwUAuFTVPIGrylsUU5vAIZFBVgzcY2LqkWjdKQixSV4MPm3+7XJRwKQokFdGNbbc14Vmj8cy
R07+p75Ns6IrYQ4rkBwAzzJMLO63UuXRj23ZbgAqB9AAUD6TvFQWD9EKwpmaeuK1TuhEfrT5o3JY
h5xgnNJrTvuSc8b29+EqNYVnLwft5VPYN1kRRatWezseo1a2xUbxDEmPiAxCGXWXWGXXUlwjpq8S
PdyKo3hSbc59PaDZCDveA+Zbj1hMQMMBgzpOpXRVkjEoHKsI8FENJ4QXhjTGfqOxNpEhfF+twfpz
ISZxQZ3LqXwMPab+qq9Rq4/+/OJv4IQfAh4f8DUUo1yLqe63Sfk56h1V6hW+O61VlL1VLahmqbQT
CK1lCKcG9QzhbQb9YxxJz9I1v+1cbd4thaymax/UUHvej4g/+nih9yfLX7wVWGGZKgZlOEypHyTd
0Yr/kYjYddrKo3d1ozWHyZR4/7MB9rXRPjVPKRbOZlL/I2zmRHz2o5qbnYjfFARqD7+kLqILxCPm
guMrIo0n1Xxg9aVlXTKpDoq1xkXElInCr0eIa2MyddeVuqAXUNZRuSvwNBqFvUOmmj4rdQgLeTou
8rasf+8FKZcbAbI2VH7ie5u9v5TMAPJt+RC9zCcZLpMr0b1NVzKlX7cIcyS6z0zaZBTmYxbAH3Hu
yKlRngw386Xv/UzJtTJTPasdTz4/30K76BGA/lhYyp50Gh+eBOHWpr90S2c/eOlvGSLANX+sAaKZ
C7pMQxZEWXkIALzbllVO0X4bn2ElciuewD6jfb6OdwRGf+du1hdQyLI3YrCTWyiHsxU8QupcUU2Y
WuBhtjqY7APrRyqx+vhw7S7n2CpQNqipMtm90E7/1LzwSZUYV4mgx1jI3UsZk7Z3ZFADqFrsRL0s
h6rjbJFgtXduC/ltQ0kolajrlNPRqLnz7R9ehsvvI+/U1ttP75QomGYOlC3xhtRdCX/2sYmNuGv5
OXQWr1R2PboTEDKvzakKpOznYohir1u6lbz7bpWLeJyLVrHdgpnPVcamwIrAWDXx5Z2LQp7Ei3+r
M7gg0pFN8OeWUp1Vkr3OTuu3RGoSVl1Nd4o+0tFWS5g7sxsuDeANYYHCKL6rrLGExFpU3Foq7D/N
yDkwRRS5jDXGMD16+dMMg/Mkur3GXjpIL3qReXZ3zgktLSGUqNJZ/igdp2iHYPlJ4ML+M2Z51zRw
3PyCCPa54r3n9XIzyaEuOxXCYwawDw+v+gl/Uh1BebehawQ9V5D2etljDOsHWp6/6CwTfl7GwJ9m
9IyvN6KszNO000yNDoAEW1npG3EyceCtXRN1tBKBMtKI+1D5MdB78qKQhJKwotXm4ac33ogDwAKe
SN2KZKoQPdSQlYlV6dPNUE1158QfBS8dggsxdX+WL4qnVZCycovc/28+HQE6E7KZ4wDuv0h4fDOT
qfcKiTF7/Fj6PbyCoJ0go3nxcM3M+YVdzVi1xpJ+C80wIa5KWlsK6Ar/BVs0yS+1ya5NyEeChXiY
RYFZnCLmD9QGVQszAIDovKsSwq1AD9Id+oXLxrx4arcEIC+oAgqDt4OJGhy/apXrjbgX6GfVXOpT
CxjkZaTILUBT1lnKf7J9W3owvqq/WxtNpxbLLZ6p+vbRV/XbdtUlXpNbRbJ0SwoUxVdsg1puNjsa
fPCt9EMDgGiuz6u6DtUHPOQ6mT/hW9pOMm1uMcPbiqgYoiLeQLxt+nkY+dsmS2FvxFav9VWR2PlW
KxaFw6na7raYEr6isAXqicthq6eI08Bslso3BtDARJTcgCjyLT3eBYmEmprfQMzQa1gptBbvTB9x
8UKloHQ3I6NeFy7euo+4OngL9PjwFNy7SEy5nney6PoXv6xsOHLBtZmqGWuvF94C01Aek6oqGUwN
9KszTWI1gqbUXS/f28kix+5G1AkiymLf+fp4WchTM6A3F7iYEgX6OHa4Duw3vlZfrP7cIzhUfT2O
BcsSnfrofYCywOCoeW7JScO1A7XKkP3DLofIuqlHv11J4aOdYOjwJYYqlmOcprABXD9EfpVXnfiR
yhSPYJ7x3naCNnsZYBIYJXBwj7L3xiJ7k0ymjy/TaTuBh94k9Yl2Y+VsMXJzlpEV+lgHmjjX7Pdj
10JJZClyeNP9yzIfa7RgVr+ymGJAsVItyggXKtojlgq/Hu1YfyLWwzyqp0y9Yoq3VVMojFRmpq7c
dYZ+312tlYMzSw4NDghk+g35hwrpJL5KTUCCBeZRoNkLx1BmW7WNe8qtwldGXzQBWavGy7eMJpt4
s17ZDm/xxZVIHIe2iQOqPUPDXz+0YznhXg40LO5kkco5S11PL8YXKE6NfHS0FSfTNn2AgokU4YjC
UFhY1uSiKgYR/uFDb3hVjJnzrckJ/oyRdCv6qtMf46TvuCpSYF0FmUfgyPdoD4vkvHQlyzUrUvfD
VBGxgWL48MqETfLHySSZDZoKwya8DinL/WrvlYAdZFlefukAu7UN0wC2LNAUTvM4oJa/WSwvMiPg
8aDbFVi+sbSuDgZ4LXAJKY6VzojheKQji7lGsxZieVe8WMQQGBzAmoPLYZGJwYTLis8ipPUBrOX2
1bXp9rwAYcre4PLqZRLJldcB6lhGaN0/w8fSKFeGdnd7W+82g5HtaO8uXGrRYhW7Y0j7HIysukvH
mTJe23AR8QCv3MLcIvtSyE9elfDIx5rUXXUHzmNZVDIXCfiI+sNk9m4ITV6+/n3W7DDG+KeROQsw
Pf5VPQiyyPocnX9CB4zORm0I2pG5htGmjj3VPMqe5oVNFF7a9bai45Fb42YKOiJs4j5LLE2sY72R
PSIHMCm4D8dFgf34RdRXs+N9S+935p+wH7lInX6TfSdKlimZTqZ4V8ohSOlstW3GxWpbOzkO52wG
Ky1JqFNE+HALDxEacWulopUBaujaeT/Vm3ESR97z/8ukGWioIQlGsramXs/Vjfb4FUc73bVoKuH+
rvWlXfNw0ibwM5knERyRgZdbs938LWFQmqDmd8B5/6wuL/C+6dB+70H5vki4v9SDYpNniA/nsUoO
PRVt7FQ+B1Z+HDEPGN7SBZOJeHLnz20KYzio8GC4Ygshtzz6zqB10DvtbGZS3uYpg1G2uheb8/XA
YojzVc36N9SCHHBcqR7V3aoarvZ+aNWS5+t/9U1ZKd8P90tVkbosxbvBOD7KR5Xe01FVP+//3o+K
bbO0vdohZPAk8pHIOAHVHFOt1P2LzcEZwJ24iXS4FHGqDlvXxHZEF4SpjsQMuCbAF2ky8mLkKUcW
0Owri/+F89nNFwc5HEJimtU6qB+Z7rS7fBU2KmdU2pbVfzm9Zr6L/RWoaOjJc9/vfVq20nLMbfNn
YZmKGiSIV7e/Yto/a8yyffDNliBS+74SJoPGIcwmRRvTmoDJZiF64ccajiNMD3CLBCUKbO0E34Kk
mWiGLtGtxS8Zk/qqI2EZaM9KkwqEVnTBEWXx4eT2AmjqGwoOiEGag1KgUQQQOeKP8isV8T4+CvQg
LAUf9pKpF8wqYeMGVWVzebtVs5xoUNJCL33zlKBB74t/U560u0IeANMGhhjOHFb8CnN9dJa/dK8G
u98GG8RKV3Irbt+zhKjLc/IFF7umz0hgS3d36qrt4H06YcVoVJ3LPXUoiRGPffVRR+7a314egh2D
Z/3bB4tiJ/+ncAgTQP7mad2DTAOSyGfQw/qoW5vOi5m9IMfMfo77a/PFZKkLONZ/oCPAqkCDuX67
9Hcp81CXD+nuHN95eXMezQRcugnuIXejNfTUUmV4/ls8Lk5myBaLaSQxo4iuAdXkgWBy+mAmXBmQ
qMiHi0yP+2XbAoqWGpgdJaTiZd8U6f02YxZ7gSTYSJvNH8QjXlQ6CKxR69mHh+pUkSuJ3b5YAHCx
cJjRRxxXcLjbXNW/McVw5NoRZD9jo3t/NIXgoFE+2g5pyUTb5vYBzgnpUUFJCAm74MAsmxAXKpdb
Kz8DaDKM+XjpeaHVeRn2IIOCqansx8kDXZ7kGTWRHcsL2XTy4IgUKqvlXkD9Az0Whf4iOJd/vSiH
PqoRqv55XIxZedsKNRsDBzucWoYTaamczFZgPCIbolWSHAwqteOAEw/mNFhhis6kS4fDMB3NmLWN
iq2Bh2G1+gHX6s+CBdmnnqYuB5WhkCnAuDOQp/7LUXeNgC6dJR1PvMhSPP6F68ulHZ5WnANnNdyM
iaI5fsW0qm3HETH9yDCbq6HVdrJu6CSrnEFysJVyOW4S0dt0m34NNsUyF1oQI9PGmuVcyt8GBZhV
FD3MN7JkwH1NVgw5+yXsgNMbv5ja3cdNREvPPPAcCYFMJr4ec0YN6iI+pLxVK7xWrvUTRW8bZSfr
MJsqjuDOisSzL0gbaEsxCKX5iDw9ttwV3dSZl+0gSZ/SvIF8comg+Yv/cjYxMKnbiXA/jhWJ5JtI
bXty6R0QoxhgHF7JeWzKSaAubSyBP0AVhD8g41YJ260LDvWi/01fh5V/Ywx9JhxE7nbILPJVhtaP
7KZWM6VfF//toaC1TwNiH6tQcnbcRg2OmNmzSchbfwF6rkCF8HdxdRrgysDkwj5YulGBp1sUh5hk
uF/kgG3bi/2kEi/sMKQB7t8Ct8zmpjYzTcOYUmfjOCdAIvRr9xXZyE+0XNQzMbYdZAV4wJpwrGUJ
puYWTnCA3J/ZwT5uWpFqgtCrwBHjWzLHQ7YIBWg+bf9h7IbqrY0WPQowwD+mNQ+JFY6yf28PWVvV
3jk1rty8+J5PBGw2BqD3qWE9CwCKewm7QpaUvbRp3jpc6ajFErMJOk8xdDNkLMWy7QH0R5q5eRur
03XAAByP7bon0xDFnYs6894ridakLjo3OSkHFewbYYI/QelVjmRFNLhzgmCbk+naZRJ+QxJa7oWi
Ain5PrdXUGt3fTTpRKiRgR5GZ5ZX+DpOiU9+2BxtCMlt5xyOxttDcwDi/9q9wDUDsZQeVAqglfN9
x2xFocsgmW5I9Q7M805fZqX7TFmlsWDZFgKXdUrjtAs4H0EXha1catELgX7PFwbyHZxpmbvKpUp5
FE47tfnJTrdc4xyD7++WIH4nNitXy/8jQjUVj886S54Ef8Mojb4i4HLv+0hfPNnIcegGwRWRtgeQ
tvjHW48haAMx0bwtAC4xNYjvUMAM06fvQ9O3mB9UKLY6OSfOuGmnBanQo7UkkGjKm3vd9utXd6Y3
u0tUoczYXquMbhQesDyCLfd78l1ODRAIdtVZrJTKb1Etk72OiKRKr4uc4XImW/5CWY7aB4OJe4T8
xkfHRB6AganycWtUj5sHeB9xvRF9sV7RhAVx6JkJTW1wWNOMDNuqJhYjFtVeArsleTaI/QLVMTft
8P6iaf9LSCRD4nOmgzfHM0ttusq3knshC0EsQcSsMfVcayHF8I81yl+Q3rusv5k9tRPimSAZnH36
qpUoc0O7iUyAiv7wQw7s0fB0O+8IWCVrmLqMDaaJRJn5Cbn8pEp53lA2qz939+FS1tYaBHYgR/Xb
BpdNwbyiwPJQd9zhKtL6+GmRZ4FEL2/i0CgnxA+yAxFDCcgFlF5Pg5bAdBzSocc8U86FRyGTEomt
MoOHJtnu2EUwh8uGdmGZtG2pe+Y1gBUPP86NT4W5JjEk6UbLHbHHuhTq42qtNlS1xc0Nwb+5Klwn
eXfPF+Ik/wP8/HQ0PY+bMmC4ddZ4leXOuPbex7LqtQmaBryzJrzXjiBucX3L2S3zO0bGoKaphiJa
D9LVOTILwqEANR9A5QjNQ43R+jkKnBS7NiEHw7ZPt6YwTCJjVDayUcwkT3SKyZV31maUjbPOnf57
uQQUwV2n5VR0w0cYTdeyCanlHfpnfo9Ioffwfi8y4kkCcb6iz73RNigOFWNeGhNyx0OTwzSbaJrk
p2vQO2nn3/lTXPmzRChlj1avkse6GNu+q9Bav3eZiHPVSH6Q2tJ9ngN6Xm5CEFmfR7T/r/BSkHDH
mVecLj6yyY88CUH9ZteO7OLZaM7Ivi6NT/JczwSNySqoUNMlLCi4I72sunZEF/W8Wxe09PaYWWAN
q3TGRqWZnjUX4+/c8QzhHV8lqYNqpxysQJ/HvueLk+tzqyEtNSP6f1llMyzVq0h6m8J5lXUzfJ4w
0U0TQKif6yUVsH+gaBxRq1GI/1X05UG4elcOc6TuiqggIjpakRBj03J/8aU1mgIWtZfbjKSU2g+g
GyclXwC7qB/Buo3etVs8x3tG4eDoZv8igMlRAL72v7BRGhPNch1ZQROqZJklg9bBnye4ek8389VQ
42PbcLdC9LeuU57P5TDqf4Z3bxRuduljxo7eqwKtkc0sRWoaATeaWU/BaG08jHSO8lRUNN9Jiou/
Rxg0tvLepopjq74+5c5kU3pGKyxugJjgWdbE65TLQDHpp6Er3QbVPvflPgDre+UVN0OU8VQD86h0
azhlAoBmDnYDTNibqA2B5VCMZDgv4woMZNbdDyp2wEoq4f262wc1A3H47FzYL7T7Y74NABsfAp6i
n5SIWT1FEI+PZRTuOQEZVT/YjEfijl5Vgmt6+n8B5thfZWMDwvWhHblPrWZFwWZUHDoeTY9yX8ba
OFE377uJDlIw7XzAsXgTcdq/ztYtqMzUDR8/4mIP+RGCVzG8Y7b0TZTZk4dbpO5bwbc2KSL+jpVf
Pz2qC62Yl4qRVKkqh6X7d0nO+E5TL8yV3MSTVEj0CikgGp7BPyGkUeFSUyibS03O2CHlNB1ElQJp
uoA4/g8aZwffHV7XmpPoEBUUyNUyZb9n951u3zisgoAZRLwJSXkuYE5sfe3VAY7IobXMKpjpyDOS
xGXdEjPsvbo8NkE+w0iWj1f5Wn7kSOo+rKw5yFdf4up631R0kE3XLkLNHjRTamGBhe93vIZLWKcH
w7mzFfUDsjP3GUQIOQ2FDvptpmTYjCdUYoSAKvgLOL1v+Ku2NkZh/K9CezWilCSUmlV77PfkVwfr
WeSgQNf02dfTSHZ7pqGC0ZXYaPDQVIYjpJoRCIRCC33kZMQKTu3HVr/h5M3qcfAfypUx3zMhZDO8
iZn2h2+7mkYFzaT37o7grU12tQdLzvzm1uWBxcUK4hF6dRD9U4Bc0We8EYOToGh97VMuogeKq8Y+
0X2WIQvkzHDXY2wogbE0d4DN9VZiB/w/xUXh/DzguJTMs+6rRnddos03hNZ27Sc7O8RRGY6TW/CT
9x8S/tiFV21cW4Wcp8NokYkExUnVSW/Bu+ly01AFA5eL8DMsrM67xAy3Izf9rAL0PD61UDcMIf41
iraun7s8Dmg4cP5GrDoLmIwyL/PUu76VNEdHa4MRIx/J2S50sNYON+wjJM+YY49S16wBtusAO5ti
ht8e2Q4KhI0thYT9UrA0D7D9zxjltSmuoY8BwQSVOzxjNtngHnJWoAB6OQKNdu9c0CUmYxyBqeRC
qhzTJS0EAnoxor88LVqtv8xkvUtHrQEbH8ZLyiOqgR/+531TibHEMLejo2sJYiSQpELY7WH1MA1H
glAMK56uQipCJMtn7H9CJnF+MhWdbOwReht3bfyPF0FhXD0Ui+HLpXi5QAEQ4+hxpQgd32m2ciea
ZPaUmO4d8RF1Q3ND9RvVMTHEmB1pUNFYXDERjCODgbi9LItN4WIfpJKHVD5oWYxkmp0tJys/y7Iy
OU5YoiyroJSMxiHH+ZmDdfZ4VBDpReBUxR/7Uo6IBRS1bRu5jWTbOl2gFpm4vTREJjAPVCm6AjR8
9Rj7CXrtcqcpt+EokGJZAcefjgSKQVShv8Jwg68P/IGmTpBayrgtzY12D1CQUU6l+xM4HKnrAO4y
BnqXHeGlUcGOdtrhkudg8gNaE9JJwvaw1GMLdnZp8eaFCmV0dvM4FvmQii+NJt4QzEzWULRPY6rY
SUeQEw6GCmlrwQ75RNYV9SI9f2ScjpDQle34N069u4MWL4nC/NNDWQ4CTJcvil9MKYX1DFD13iaH
9r7xwFwD1Vrc0ckUZk/QV10BjoWeKP+VKS49p1W8dyxhd2ZJ2RKdF8alNFZIR12L1HX6g5Oadfsh
a9PryaJma47pz8grcCAVXl+kv1/2g0siiD1PUlCnWJFufbcEPUyZcFEecRZok1Xqc/vdE0e3Nec5
lSh04OgRQkDR8n22BcKjk3K1hQ7Olte+Nx7V64jQGQ8jkv1l38/0QPkudyQkSQGqyNvGIw0pqAQo
gyMT5opbe5WywqGbiBEsq55yZeMOeF26rm/DOw+ikWMLY9fnA4qGy+AZACn0ZcujkvIK6uVNqyW3
fVTTMfVT5dx5phyYqARR0djCoZ7aC0zuwcKeBE0Xwqy1PqxwOU4VGgrPcLlljIQZeCOoGu4LlC6C
d3ivXTltzkPRzxfG2n7fTa5oiB8OUQinAR8tzYfrHEkoRZ3nP/6t0FgkEpLuyx9lx30kmqIQzucL
O2w5fuzmqaQWQAyH62Hu+LnXIKFjLUxnaJED/3UneE7GhvSvFxro5NuaBfi5fSvq5sIk6R/5SOQH
bfwjF+6/6QhJ/5/VEy9/hasVFF4JVUaIpm0q6aunaWh3wqt+QPHL+sBNVeXP4P5BKYdJW6CYAElH
C7iGpxG5e+PUHCzGgfA7U6ZiN7DhzUjU9Gz59RAaXGj0UoYUzOcLwWlsznfHoIGbW8UjV57phCgS
94p7wXLzLeJ/X3PTw5HZWZSIlZIoQ+oCmm5ffKSMWlDnO9PsTvoJQlrz69+3EJUs8aYoR5mKf43L
U14P4/DDsbXqLbKIB4qcDh6rKeb1FiNKXpKTBJJ8VfEpqzOUJxCl09nA2ltGl2VgETbeJ+/S4Mo7
m0SB5juXGtNwXBbDWh8EOf2K3rU9EynQuEXJO+XHIO3WEFDFAa7CZqNp5Voo8sw1GwulFEGipxGo
80/Sa4sw58IKDWt5jIdmozEMtVAlfz7Ag6sFuonP9lCOWwCt/jbLt0kapze9q3Cdp+G7P+voYaeI
JuT1/3ctWfbCw1WIJ/aMifj8GUATDcj9G2nGB4PTM5UXs9vCPSVSq/DdnVGkEVY9nVve+1yHZwT2
4Yz6GkadhLXuiDLu2eFVfdaVaYsKR+4vrL1hn2EfKv5Mf5ceqSu19CgyX+EJjROuJmGuZL4NM7QO
rLNF9r8Uz6TNnGMiH15bwv3lYEtqohdXFLbxPWJL6nNzyJS9MVa+sdwlMnu9McaVpII85wiBixAf
UeDXW8ZTJLJow8BkkpEshtl6h/rr3KN+IrsPam7wEw794rn5dRiMotOWm1NiTEHvc997BqT8onG8
OF/ViGDf+0i5nzf0Dv9chUTeNMKb6mXrT043WmnNYj0YUKO1yTY4QXQ4rAYRCPaIATBWGjNhnuny
jzE+E+Iib/9lgQ+bzS0ykIIZ4Eyg14Wxdc3bZT04BUXMgMgsFNroT9goSqsjlSz8gj+baQ/JLJJh
MW4WP7kkFENQR8ucroHHYS80HPhab46EqwX6KoTe0cwFB1PgzvTc5zktErlOCNDktoZnyBr3ojCE
52969UjNec4MHyzQ53acEdAH4FdCC7LWm5mK3oadAwlrnHlVaLsas96p/OyQQSYOyeTfByOTwJR+
SMA0apYk/IJUI6dip9axxXA9TMjGZTnepVsPDIQiQ5DqhC3I/tMmJjxL9oPYkqsBq3xXrAqtMFYs
MK3Uu5kGJL72/uz94brOph+E5aqdma+C3pNkhw7f7g66nBtPTNctZ4KuXACu531t2Ft8ShsTFJot
aPs083BM8ksWXzgE3yutcYsS8uv1GQHOdYrZmWRjLT8xANcJ4LiowNH/p/5nyhSG7QZ0MkWvyZ9A
MlDCCc6eVxXU8FFpGw59H6L1Psm/kj1AssqNEJ4xMi9v7vYZf4KQnJvRW5h0OwIud8dqPZswmvKf
JYjnul4+XNn0pGMoJnJPweTRrAYHFGo5eS9lKUGCCLovw8R030KEcsn6sgImCnEl80vXi9Wmiq7P
sA+DG0EwrEdxXGw/DGHIzPfQiJ9hqM5TDBC0rjiOvXwNpdFKsOyPMjDqt7FeeDZ0VCMquX39V/or
nvpsX/fhTa5mFrCzwaIPUSKn/1/cKu7ivBfn1dwkSs6N5Kx1Ml6nGsDHM8T1DA6oFbWG9e43bdo4
0ISyv15FPCqPALqpgFziahPyi8D+pZ05jMP2C0+chqveWi9+hKRV+wzsxInpXrlH1A76kcF7Hrdx
pPKOWMSQJZL0TppJZn5j9WRLv0N4r23AFHPAC61+nvbBsfaPwfBLz42+/IjLJOeD3sLMkm0UfhHq
UpUhf2Rhk9iNJJrjw/DAfOM/Gu5tCunJgPyuVHOFXMEJjxm5SnARnS2YGaoN23LP4H/1pNr8p9Hb
llpA6tghe5PlUjxnIFut6w97o+npX7TZyE1pO82IXNrWWLgR4pfj6k53qgqU5eFAQi9CtQowXs1b
SDluEu3adfKeFskn3eNLAzJJZZTFARZsWyVcoi+eaI16J2yjjZSGisqTYEVOewvwnKFiBl8eyBiL
VyiiLwWtADKcESMXq0AR5zMMSRZF1M4FM9ViBCB6IA4urpGc2gM5cEfv7a4PG8YFieinmkwoI/tu
OPmPROsKanyDDIz6XykfZ7Aki/311MCET4OECmq1L5wvb+VYLnlv7eJNn5bnImL8HxLfLf3hnL6H
niHtCuBiEhz0y9pI7DuD00+U9kEcEN/+rEawz2KeyJpIxYztrORvojXYpWk6aQDbbafrQys+eroD
TfxlDCMku/4FUIyyP/OVFBOj/vqbc6peDyqlIbdOWwGDMa4einajtlkLUnslSfpbTLogdKfa3ETO
Ng/dK0Fos+bYe5ZexDnZFeqBmzC7MHnLJ6gkKof/ILU+LjzJPhBWoRYi2vDJrp/QQhM4yGTo0xz4
Zscrt7b1oukzZb4/MTRbLVXeOwczb+VUTxrGkUbbOEnXX77Yhyi7TxhTG3wrY02vWuhioIJ0VuvN
TXjd3rd8MDrUUSIxuGvkoVaJnkl8ozgDf9cHNQTYhmq/gawLGtTZhgyqwPeeEZZpugPWrpNrGiip
AyFwTdPeROvRcx+8q3d2fe2plF/novi+QKNshkphlF8/BSIsgRBv1BDKr4BINLdpvnMmuE8EsPy/
Taw/yl6n+vux7jfqoaIxyB+sSs4BLnp+2m5pH0/KRYQxE11ADu6XFR5zA4765IWd5TpWOKoputGr
yNTq5dvXh9enAr6/MUKNPY54fv2cv/hM3or3uY3pG4zW+HulbIxzL7Az1X/uF/610IvB3wn7NjTh
fQo6Djyp3zvFG7UJvvGWdnl5FUrSyLYZuvj86JiFsuVvOgQl7FVmRMrawdwg1qKFecANXKaC2Ixy
7PQLOk2S/EqV5IDJhLx4WtvTBf1DcLbevSYLIo4mDJ0jXsoVCarwaCtPeLl5zX+XCDXlVO0XYXOt
KRIBK6dy4+Wh4+hgitOlnTqdXFbCThJb35HyZ7Zum5ZwU+AQWIH1S/YQT1sZsTVnyD6vtWG/QJAL
NcHWkbx71WHbKleHkuB+MF3e/Rq9fP9OceRyyzlYxmckapAbWYyPL4hExb2RpFhWfACD1d8L9Ol1
L/mqo/Ys21/Tu4GqabpagvPs+Nhy7YGO3IYod22xiLQ2tX36I8d86YBPiIZAyMh3Hpvk8mSIhkOV
SW7O53VXN3Rm0X93ANvSMtzf0+LNXPTectjkihcNn5QMl69uANSSfnVAwFQXRj3m5U5xzBIwOiY9
5LB7wd7tMUHLrJ3rRBABCJ2y3M+ybghixSyUr8HL8y/ec2mnvm/stM1E0CdpF/4iizMobmiJephs
jXlgR+lGf39QktdKRmnIXkTAdfbFAupJPXDcUmuvu5+qkUvY80tnAbUjwJmkbURTVggBD1ObokZP
u91NgrBsAGekZwkDSvnrq+xYKwaFOcQwDWplIWICKx+ZmrdMoxoxS6Isz+aqwKPwzw99+MeY1abi
3AuLI7eGVXMa8WaqEcFcDyBg1VkOdAoPj3ZWFduQlDmswL743fVNZRZ2HwMKkjYC7ZQq8knjz0OD
LcsitIUnKVducBkvS5qb6oE594F8GobxwOKPUSd1fRO/P00cN/1Culs5gp7CapsbJy3erTKZFMRu
W51SOQj/pZOsh8a+A7GKsx7fOvY300rovLTJseiT7NSn9ktCGGZpx7yH7PL3Qn6v1ZeCEmYGgVXm
aE825dZ63VlRlL8XReVCIesvWXEaAGqCAcyznAg3ZhiF9WDQOfQ9ZbhFb2OYcNJ0RpCbhAaNlTo7
h1IXYJpVTp5T1umHgqtQ1yBMGQr3mvSq7UB7tIfbwKhsnm1uiMzchXU1XZrpY5d2HRoIb2uoIzuI
SKdQlF8FAHJl48sHCGkL7JOGR5B/Z8I0LaY62slyrApjArRQbURdCXpcoJlHV4mH/qyNgneOE00t
oVENSzAYW4xQoIsVoNm5dFsklPcfELsglHGqGXTuKq3bViCfzNz8v7kxfRx3oa4dMbt+WCRj5sgD
V8LdoyX+6oMuYPYYwmJPaZXyOt3FrwpaEJP50RykIVIwOVObpFNyyqrX6aU0A8KX1C//EvJiD8Zd
thvGmhZueC3CuaLiOT+KQhmS1u42vBkrzTC7fTufcbH2I5RVb1b+1wkEUrkkkj1SCEN6mcfDCBJ2
8unVDw0FiTuL74LgvTGbW2czwvYdVfIUGxb4AkkEDG9JpuFiMsJb+KSNfYVeFPiGdKnU9deemNoM
Q/r3oeqfd8uHTqZGDBZNQd7iyGO8UrALf7IhNGJTPqPlT+OiapRZLWzdFxkAkPULtWo6jzeauFUV
LGTHP9VVsGJOapoVMlG70WM7/kEgHykRY20BMbTAYI027OflxWjCliaHSTMFbpFYVwzHQgOeT+tF
wYTN1HihdF4UUCkrAwtL6XrhoaUJWgsvEV2vKJ1ID0QElIqIUANfL+EYswmwam/bbloOvOY9I/7Z
EzyzzJr8MtN68zvCK8E0B7qGJWTt0SnIvJ4qF2A3Y3LI+Mkp+6n7ZnyiwZ+aefgP6hUac2AOskDc
v4fFf6wwvvBu6DGLtY8AeZInMTt/uTzSjxURT1iAOLScHnAaaLtfpvwc/AvZ6oIcrhk+ANVlsd/I
W29JCQkEk7y+/LChOSyNaOxSl78MplbP1Jx1nSMIYQOWU2nXdu6pnNDNby9KEurBRpBM0Wv2FPna
CxhiB22FBzjjr0BtPZbxPftV/Gd00E2E5S3NSwkw7AuVSm0TZOoNUZnqFunfTlGawzKUzPofwRQs
lJTZY8hAsGHjdmccb94d9FviUrBtK2oC8DdtS6iUStHKCE6CfNHyCbiveyhSoKStISel/EvlmxIO
5z69Nj3gudEItA8A63IOp5OSXy8jcLCtkwLLj+awsz6YsXRcmRZS/qpk7cLA73SiMADvHWxGzW/F
MrpytV95AN04JUU5RFe/P9QfK1sbIQuJyyzMs8SxoBZU9zb8sv5AYOkvm5Dkg41wfMjyZgORMGVQ
dhQWaHfFodKWjOjEi2/NfpZjkHaHKNaZXYPDZCfkmJkAm92N7Vu/AIle/F1kXv2RAK09f8FS1hfu
jR+D/N+SO41duEtUhT7hc+87TYcfjlDQhLFCbgJ0ToECM853N0mFChwk20iRKtW8Owfd9I/zCCnK
gIkMyTzpKMbkCBAJXCHBcg94uNafshQ47gJ5R16i01DUGfctQDPvRqkWQW9u66HTYclINaOfhlja
oydOESQWjWHWaw4LM7mfDnRyNzj2rWUi68WtxzXsHisrJKS3yijE+oJ0n2y252SghloXjp4LgzUe
2Zzif1JEdaJ3phVgWcd3J3Klbx/8sMTQR5oa7GGoVKEZy1tj9Grp+N06yzw7WMHIkj2aNaJOc1lf
WQKFYt+1w5SZJf7gP/LF817dDh7lrY7f6AG7XuPEoQZjv7FSSpedo43DlcpjdkZL+6WJRICKKdmB
VWfyGoWlkdzvs6vG2+nM5sLEMR3Ti0BQjHmflTM6otN/sLWc1gSEZhaOTzfvGbmvVChleHI5LSgY
7NhLtSH7E1k/lzUVWsLjz1Wf1eTU9ViwW+3NXrrBjsJ56DaGzruz9LyjKRp88PDnt4St3lZl+XDt
btM4EQT9O9SCh9cGSU1GdRbPoWlQhqIYBFfmQQVN1LVzot7vCxdFGLQ/7U1gG2X1Ey8DW0Md9PMx
nJZic9R+RKCfFXeuvlnFFKkVnifHhO/UFJitYK9V9222e8+MnM0lv+yhWyb6++gM3HZik69jeOjj
FHNX7A2ZKymQi3fLcq3ePTGMiNNgXaZiaS8bxLgS5f3LRk7bZb0fyjZ5spGHUioa4NllVW4Z6mPt
A1QlOgkQ0u6/M9qZfuaG+CipR/a/sf/7fYUNeDCdwB1fKgcyrsAZ0pQ/ShQbzHeIqDP4IPajmP7d
hhVhJm+RJ3ciGxvzkhfVyCQmbIMFt7ig9pRBf4M3bMK+yBPQsA19Cybib2OlcaKIr2ktjBfWQGw2
wa8E2ctzV1KccCz7gX50Dim3A4Z8ll4b55aVgw9AuxhilGTGAq8YLPl7112Hk7XII6nKLpH70xTx
FJNhCVvpidmAG4yCU5HxQ9qMIQ/N2LAzPj7GcuLQHp1iEAjtoGZsEAAQDfUOfHucO0dsJV8FQvZu
MVfc1eJoBPkOxKy8EukNsHTsBsM1tLw9O+GDPSvdEXwu5emhn2Bv8JqwIPpkNddcXbkOb/bfS1ad
Un/32Zt4qZP9JsCe/WjBjZq2LE4+T9o+b/5rBPh04wJWLYqTk7qTMG/cot8ALijBCs7pl7NBYm9F
UKdsA+pYiJg0vduqbDO9g6wsuMZgUSGwjMTfzl6LuHjngeqRXjReRLCGf9NTxk2eT+lwj2rVbwa5
j3RBp+ld+qn4AUwQuteBaGl0IU/EMN+B7tZEnoP4JwrYEa8MDEVYgVkbdjgB3G1yw/balD7RInbC
CHgbfYuUM2D47IeZDGLbx8P9zw9M/fwQloiZztRxn3MaPjOSAx8fCghXsgxnDsdojkC3sb2l8VWI
FklWCkl2uf9h6IzBhvp48gKT/3kraVwRJjL1UB4yVXXlsqxBCc1SRfncQNIU18si4QVSZv2FEx73
x6tjS0DOXy8qDO2sTGPju59/CC1vAvd3IMr0a/wRgBTkJkXNAH/y54WjG+kjB5+tlxqW6DBRayZw
KTKxmyLbDE9qbyTzL5O2VymyMrFsTAMxYJQ61e7eTg6T73ZHYzq5rGDnzA2YhXrczDRurR+tRmRk
MHqeM7XBshUCOi9Zj10eviYsYlCEdl3kFyIi6IJ2d4DDUNiusIyd7h5p8ORbbE8E7j+Q+a4PpOvS
B/IQ46G3L5bDuUmExvM0H96JQimEqMepdGCn0xYeWzO4pW6Cp6INVuUpm9q7Se1dCIqJTlY3bdQh
eMdZbQLPT4CpcnBzCUhkPNZ0rOiqH8YripLbV1LlkgHQlnji+iVGcbQAxefIkzJQXeqZz4hO+m/2
wF6jgbWR2Frh5+byMX+pNdtTp/53vsyom3Vnw2jXPUou1oPh02V/4uY3AW7Z4KzIzk4owHmUxma4
nFcXZf/4FtCZjnuZE9OR8c+3/z983lwf9ABGIrEkktzbkxNPwnHtMT8uoKmOvxPLeFiB/j2J+rZS
icQcTTdJC2BSVDHJjkfu04CC6Ss3vKJDLfLwjXppOuPTA1xG2hcZzg53zofabH5uYLpeWz23RJ/y
ASnoTsnZOcbliVXXWLfIwvC8XDyJrNPop92biaqd2+hjJyXYA1tqzsjV+dgSRHNrJjRh0XiubPp6
0bzI08NOJHe/UCPi9My5EH4Hc94Ib3r1AJ0JaoJU60JVrOVwqVHR2n6iSLDhkh558d6v97eHUoV4
2e3t0q/91lQtQmB6+byuYay6HeRbSrR1EQWd3UUAYhTlfImc30v+CE4Jo6rCu0QVXXTtHOyqsvWc
eGhviQlS+iZ7fekue04FQExvyCQBKYc4z5NgLz90Hg93NWrs1CeX2aYr59yEH2Hbju0bvDa0bhSR
bNcidXuXep1F/LEFTz79fQ9A6X6MKPdPqsC7MJPhHnJY9vs8I9+Gz9h9m1Bp3sWLMVufc7aXSie6
7N75BY2cem39TrBUloTa/zhf0/e9AxxfiPBCAb4EwgIm9LOKQRe57uV6htkfgXgv048fASLwV8Fi
guLq5+5kk2JoHc34M7nmlsCB1EXi4uzaHv0DDjXrhbHuXt1Ber16TNs5YgyALBWK6Xdb+pAF2IKg
ahdKlkn/5wgCMWBiFbEac7WeovDh/whxiU0Q3vB67UmqsCu4tnyAPnuU1WYYTAeIu10SWH3w76L8
EGbNVtufiAeqUkZRQCCVGcfe7pbinsUbo+lq4a4QsM8z6dla2OvHFPy3QT7Nd6LHdTrK+udZ96bF
ypH0D57WOz5aUb97EqzDXyO+iSVnreuIz/76xInaces50DAeN+f10o5EEdxgcmjaeo7mHUcfR05d
gfNqFpFCWp9rEG+7YrZc/WC7o9j/W6Nzbs8bjD0/oLNHU3W8nYjCnCwmEMJo9mLmvyfUzQnr8s0n
V02z0Nkam3RHTHkOONIOQXpjadH3+IfylfKcAUMO20l27gdDqzCWi4qrEGqtPRsU4MP2oWTWv2D4
i6bHgrmKrBEiaLFtwmOM8WYYFqYclFil4qmvh7C7sp65ILliPJvDG+KlT3JAP5qXimrpd1vT2RYr
oVzMMVAtaacHRiy5KFwMVkLhy+8H9ZljYOP4tdSbDQt5yeyLxjUQj2KjPT2fCJkAFPUgYISzBmU3
rMtYmXVJgSkir6giTTAQPuto2FaZStG4TBEl7i2c7OGxV9L83IpK5jR+p0a0khTahXT6bjdDtmLT
hHxigofg2q3T0rMv2s94v94Q8gGxoi58FJSbf9zXw1CqvhNcIwkxgLvxliVRrhdYTxW19t//mUaz
0c4epYKgVCiU6g4ZxYeToqnZEsFy8ot0vOZ6/HBks+RZ7bsrweHXKmviQum0Wn7bSy2fGSwYUTF0
vsTkYBrrej1fWWRliWsVABKQLKjn6ZCVWQPNyduvc4NW5n/D4yIne9BPVKhWSpS2DXpgsmYvjxBP
orW0ld+BzG0tOEK+c6OXhKalQ3/nrKlY+rdVU3GMUKPBrznup3owZH23s+g0rsdups0Ndpaj9ScN
uievEcofac9rZt4ryOXIJ2XiqpRPtuMUoORrnFi8xg1tgPhzAmhLFmyWDMfMLv6+UwlFpP5ba24G
MxUfA0290r9tUg9KT60dUfO9g2NF5r7MeugMJDiJhm17J8MyiGPi6K93L94ZfwVH4Uir6j1p1iel
+lKpnqorC3fgdXnUGuFuWs7IDkPbUG1QnY4KsdWlZcoLkIpGPypsqGEqxpz/f+T0mAedPlH9LpYn
ANOv500qBFiMUxjzUUu3Dqnj1uVUMPJ/rLsW9KVHTLI6G1tUfXx9/eF2Fqyuu6xl9WP1LoVSYUfh
mdjnPr8OajmTxxCLWuLYXXAM3IBe4agmMmtK5InNr2FIULOm/Mua2uS6F4W6X0IpiUAxu/IP83s8
RtIpdUMt8eQDxLxc9QLjr71TPVFTlAqt/eDiROTzoFsnjIZ0NCJ2OxmGTGHUwR7faNT1EQCkD8V5
lOncyW7JG6M5RZq4nPMae6AhpBRshK06QJc4ClQcz7o0R8bP92n6oJvQrxKTDMgRc6NtVNNtTPhg
S8Hh8fL+ht8m3N8eYJrUWOQj/WJ2o+Mf2jN6s6sfXQ9ZMpx47p36wNxy0QtQ1fKyZmQ7kntz3V0I
iAxFcfR8Y2Hh8lEganngSaO4niBPUZFabzDJJVIwe1kPFdHjIXeURPmGK077tumKo92IRK+njsv9
Sm3mLRliqkoTaFRX3Fjw7bmQlPRw585Q+gBHYTzwZ5VQ6Fs9riJIKKIijv7dEub4Ay5p/trx5UQO
UWGzdFaaeW5nGAtRqWnzcdMhQM2Qr606YneLDCXU3IQ5a0ompfkJSCj6CKbUjgnrbTIsA0GGrWX0
fIP1raAMxYk+u2DljCJWiau20d0qN8bUlFIBqYANRfmEDIUoHfKUbIqJhvgTIG22RRvoHKv6JSyU
6KLFg91ZT5c65hHL9gEZq1jUMVOa1kluF7ilnLzaVHYODCgMnHiGK7Z5QSXcNCWLxpnmptABFVPr
kgkAstaP7oyVMMl15xoeVuc2Fl2svb3uxeWVyI6LfzIf6GB1XYXdKurasOTIJuK+XlJGubD2rI6t
3r5yJ2JKBU2YGQ6HOuHcx61su41CceyPuYjrqZa/tdHrbHp9s/BxJPgkqEZ8tYZJGi8x31NHEwuC
R9ZzvCRNpWOcT4mW7i2hJ3nySK0zdVwnSQLjcjfO+aWC/EjX1Wfuop1zEynISHTq9RhqamS5fWiW
xNTRAWxPcdoDtwUDU05OkaJmkXYzykyEL4NtcmERWtCuJx/mDq0zPoueI+I6DBN4YLLU7LppqCp3
BFE8K8tAZtzBw/TNQx5v7ZCxtEhF8SAATONI8kX85sPcPsPK77Qx2vZabjzJkRoW1dM2IuBUTbLT
X/J6pMA14AYdNEHi2HQinRct5d98R3cxNX2pKiGBQIeRMrV/cz/Lij+OcUoW1O7eprZvDF+FuSMG
avbwyToXrGQnqj7fHam9/M0Bl4+jx44cjvkVOH8FwdVkwgpeGGYpSKatNgtvtdJmoVMc34r3WAuJ
j6J913X0Z3OjG/kt3dKqHkfF+8sMGULcsImrA8DHmFLWbuPMfNUnMXEXk+b7Vhk69NsollwaFErz
NmfZUOd7QgYqMtMFTqEULkglDiKqXoUa01404CDT0pF+JlQgT4T85TMlEZJS7OcFSoP5z9R+UxJY
5NaLiDgxrX1VV/Ol4yeMIL0XHpi0PbPGJi+rrRGKo3gb786/mif+Evrx2MAcUiwDcAb1J7EjHg6p
OjXX5+eF37Ypj0QSqtCzOviCEIpY4fosikHyUaVbXSQ6SFSvDkc5Np1LBpxrV5FDn7uNaaXQ8INe
RCRUg8ovFBgdFzggHJWTrnH3h74vK6v6YG25HjUO2ZDJrWbuTVLCcKw/1OK1dvb2dawDZFNZhAND
wyuDsGWaMSACaasJY8yq4h3PY/SicZgHHpvUzRI8Zxjy6aSS/qfBpxwPwhDlJ+HqNG+kNPK6U5HK
iBp1KOwmYPldGpvj99QL8rSnGZky/f7zI8vKlQLuZ/pprmIIuD2p75qtrTqKuiJixh4RaheIrf7i
zYgUVxH7RRDEJ5LUlVisqXQD1qj4SMvd/YM9jpctq35XbcWDmuEAqgOni4z4iuS3eHrJnnmBpZuJ
GeiARsBUCOtj4SLicOg1MxUbr4USSV1ip16RxdTXVmOsg9crCggiSYefQLaXwcJ5C3VfFZZTV99M
OLNTEwHk1TShhYtKEzR7tIiaUCwAk8oxl6FH9y7sMf+xnr2EahqIH99EqxQEq7jc6LwgvE+h2Efb
edCvY2E7RCUfng/lMBzN3L3vPtmOxqZ0hhyrvkLZoZKsH3n2PW13fLd+xnJ+GQGZ9Op82zH6LsPp
3EZ+5JBonlelw3S5sgTj8t8RMSeYKmAdKx4aS2wmBKoSQ2wtZ9rL2W022xxYHIZegorhEnuXfPZu
j33QSmtYpkW0mmEfn2VF3Q3FfzkFtOWpCoC+IL2g2siXano41xzmnlgzgvM7lZZ27f9q7Mgq0JKJ
Ie6x1U6IYx8lswDp2Pyua+WTc8ENm8y1kVNyc2k0Yl1w/d8vnLzsqzZdImStJBzXpHeQEPyiVzGe
xBv0aZRE1jJ0KkDttI+ofUceJKjXGLBPTlx5uDx7mUfXIsuzrzKMgJs0uoGjJvu8LMfvnJI4/lD9
bxlEUp9mfVph7XM22Akjx+xvrhhFWbwKsI63VFhJ480FOW/HssuolH7yvXTm6+WERa1xx2PDvXY+
CkhZrTN91WNhjmKb6f5rPN48ppr7pX+RaV5olwcmZcU+zahe08enisVpipscjNEdw5/UDQJLbcQf
Zq/GxlBWy/OmTkVhn71Rf0G6DjEjut9sT/QgCkAGRKkdoyTCY1SUuG4X/q3piBrr01LZyz3yPcyK
5Qxqzk3yh6Pv8XqgrU7OvBcm4nPx6gMmhHvydZyx++nIM/teOoUM+HHL/fjsf3dZ/QAh+lxvGu4D
H0mD7zUx635GdYe7LSnNcOb6a14Ga8ODq+w9V6JnOQSl9q+U3hBS7hbSmUFq/OkK5lqr8hRJc5Sd
E6PwK+0ayF+bHsQKZ35/RtyX/mT8PZ5hNbJZ53XAj5ENtRFTaHmoP0Ql/BOdbf5VBZlkYKZmXlOq
8S6l2gAVvdfu4Oxf1TD25+o0PmhxZMwOIFrhXnGmVgc7LDwjtZTgTgZnUbPgYAOnlYmeh+zKP5qP
lFoMX3ngfk63djYX+GMXp+sazY+Yc8OqeI+5XQmqEaxBJcy6DQWOJk0+0kI2KUdlL8eCIZxSBfbk
PkJ3xRXaes4Aw4mDNs5YOJdZHWxVWKQJg7OGRj8W5XaddU5RiZLoldEe9SUpIQ+d0mZb20qv2mQS
VzntHQjFrfpQnW+/45eFJ1X4+uOkxtE8lkDbzfMYewLqdNBTfleF4ExqVkuXZRT+EC7KCkSP7Ucy
zHxXLr2bbB5iWx66xX8iWKMEn+MMZqOgESFfUuSTO53OETKnTDrLa9Lw57cjKpuiVI53Dd5nwhJw
LMdL3CLXp/tShuFf0xSUYZXZ0DbIkjORv1XOm9vxa1XTP/fl6/av7hUN58Ud0aluCNgZ+pOBqBPQ
uIhZmmsUNc0TXFH+H1/ZVw9FQ/FDwFuLNjpzOQP4mKszurxguRlORfFH0j5rciJ4adDLuiN34Q5k
GejGi1P2yihBGzqpCyPkuSydWWhvjN0F77wa3Gro51gj1iMoX90XJOCp3ad4l6gvwB2Copn8i638
pV7YaYZEun2YFDhYA9z62noQTOi63pUXEnIw5Ea0YksDAX7+lfEe7hL+GuFvwMyGYujacx3aBC2l
en5Mf18g1R4APi25y7NCe8y3GnUumENnbjJr/7vKrvq7H5QPkT6LtK47qZTBkqMbNF/Ir6rIIg8A
ZvFGKjXcdZeWqLPc6vYGwwjeLjBZC9DiCTAXphE0xEEzv71IdHkkZK2hXxiuerk0Tvof63VXp6+m
s+GWBaz7T7PjpgxwegnL2M2aGFX/WDRO0oZRaZetb2/ycnimT8yy+mCftNGzNa4fTucezB8w0pH0
dcqEbwVioFK1iHJwYv7RBKSxbLLoThwiDGoz9DVgATD/4QTo3oxkYdQ96ZqmrravGYsYmWwUKBdF
aXA8J2njIL4ejHB51eDj1w7mR788nRPJCRQnjcmTFJSZqLV8ihhGeanvnIG9wi0y0YdwnxFAwS2X
eWXmlRnf5R3K7nhse9z9s8vLK7+tvYP+1Rz18n9f/h2+JWVPiUxM0L+Us7tUxl8LEzB6cq/CDOsW
b989tFhr686ipV/FQhYTesBD1EAPIY+wSm7xBzZg+VAfKKJmsUB4Ww+0TUa34ULetGc4FMoQKjpy
O3qN4qKgVxUSmuYCGzaGB7Cn/8It7sBIflHJRaGzV3BIXhKrbeYx56/U6vN11L9h7kMpw6Ga7rmG
XSVoiT5I0bbe0Cecjpeuz+lwL+Bzc/CKWkFG5CWobWSz4i6sWWw079sTcj1XQtFiKNKJ3uGjDv1k
uSEGVBMRB9vjxaGDGD2Zmc8ZJOR/2DlKErIqWxAAT1bIUIIkbViy+8rJtlpQEEQ/H+YpiH0YXkZz
v5Mrzdc4crLY1/PAr15D8IIMdZ+EH6AwruLjx+4PkYDRYijoT0OxNxMmC9kyypLOdGMHP3IsZhDi
KU63xnQclNX6yJBCTdPRWO5/wNBOpBmZqtN2Vgp5ECmI4YmPXmya+Iygafjvv0GehOwx3ddFpdFh
oYJ204Jv9+QMm72Q0hUYaL08AvuUdDrA2BSJ7j/pDb+xbEUUcX+0zFg7hQM0uh5ob1e3qB8M5dXh
D9XjHkdrVdHKoXynHTEwiXShtCuaa6xXnJsVA7LYZ5qtBiNVBl3Cl5FZMk0TCCCxl2eXHS7wuUWm
pY7dZvYAkrlXotDgblpqb5xq+n3Ra5ql5kCRNxNmYxoDaYhQ43b6SQ574zXam61O+DwIPGW3IYUd
wYocTiarsqQ99I8DRjGVL08ZWTOnkBBMHD0No4x99lGsXD0efRKz2F+yJ/PW4U4o72tLfJMH4nSG
lIoMcVX4ydgOirIsk3bDRAvYx+QHv7F6THNEb6V3u19nXRU8VNSYXDEdRO8gnVK9T1bfBXe+gBWF
GVKEwyEjUBZK0IUgC28/iPoYUNM0y7Xequ5IFUHbjGMHwPpd93cVHFdk/f3AQTI0ZacAHi1BwZEx
VtH+DXHJkmn+xDD1ynaWcMD9vxzrRz+rwuU2HQSm5j0/isajGFShapqd73HQcFpekS6MVzh6wNZ2
M95qVgapDS9WJn9hDfWW7EHKUzScmWPRP8Za2elnfMXKriq/UmgOzQ7h3fHuwaeqT5LMzQQXkvav
UTju0bcMKand+lcR4dC2wrL3Qqa1NGU5MOPBCBBnfXIfRuCRcPE+49EbFT2hCBw3YYzvfqTOBSls
UkwOPBJCtNRGbvOuXyZQJYSgarh22ys5yMz9W7XRzu3Za5iY+pPEF+q6HucgUf3YJx7Mc+yyOEJd
/ktmQ3YpzzzdprMFCKKPAEBewkza1p52BgDXloKx27wtX9pDiRuwZS7HIVz+fvx/wyla6WoX320A
zZxlBm/ovKkXKcSFjQV+bIat9REXRUiSosoDwzKcTweH+tSQ7SOkHnkZAEuaCgQQnHrzupkC76tA
BxV0oZDqYOImv2cSNAiTI1+JSM3AzrF4Jrt+EAeJrvNpQdjdFFyAeVIYf8+S9MK74AEg74KRCOcq
2lo3raNsdjhMD/BxmcCZmoS8lQftAprgSI3WY5XH9p3oYQi8kDWEtvtb/MzU3VgbG1KYZhmtiwo4
Gdt5bAt1GO6IOu9SVHXjAvZ3XZDL5aMpF9NTkeAJpY1/ifWuJXltyxnd76hoMnDBfiJjAJQnTXi0
cqsziOzXX9jFBUzkOd2CeoYS+IJRrs2USULNgLsnzesuSVyhIpjjkYkLIyguLR5z3+34wBSWwzZS
rboOM2cpW6a3J/8VJeoObavwdPIEFLIolJifEkvBzeozm06/LXau7OjpKXDqndbhnTF1olrxlVOj
KjShqxamJ2swfQajvK/D7OA5dlXWWWVTBu4Vl+ABzLI/uVZLzucnNwE6sehrnOsUllc1qx0Wvv7w
MpfSwnuNm6b3IKEQjipxchaQwLvxpKtw13DMfkTaRgbEgMfabmY2X2GL0TO47hWyHtb8CijjerI3
HvCu4V0EXGRPMHt0lFFTys3Rrru7UKQVWo9HjZDiC+0cwaf6hZOdC/F89n/bAod1V0AZfH4P51WD
HYRg5P4BPAJTtGSj8yGVZeyvg+ecNhkXHuDgvr+F7fJrNmR55KGSoFa+upCyQRPa3Ubnkn3iaDYB
5t+sHmGEFO13cQBoFdj1Dq0pjHHPvV4Bjp/R7w9linnuL6ROH2DcPpYuBhFPFumud0xoaSTbCOL3
Ao+k0mDGP9T/bz5Qwm480waMsetaax45si26RuXcsJ885VKuUvyfts3MvGRbp6VAjlw47xUV/f5K
es6ZNmmvLzlmNRu/NoqAi4WE8sLUAZ+0FT2rODaYtSVsQHgmdcXLzroSXE34oUyXLBw3qCl42nbv
O11UZVoTJpsEwxHyV9xZ46PlitB64tFSDwHpecHvFm8672QXJrfyOryVstmjPeEdWg6a6pwP2VKv
9StTxV4f+hUa/Nnz0JCLC6OKtBEwo3nRmXMwPlqnXe8RdS3bL3ccawr2CtV33ZaP2kvbTNJ2Pm9z
8liUeKOmfnHnVCTiJ7gxzAnqHYxEPUoTK1ytYm5N9Azpa1aVng8eI8mxM29/3T4Wf4ZN567AUJul
Erv2eQ6UntLK7KuHMcWR4cR/UwYsE8eoZaHfnaJAzw7NbeMfqcAHguIdqFqh92WrIAp1xQh78pA+
g+qSEPNHco7uMxeOXzG5xMuDa86C+mZeC5nFyWD3TJocRJiiKRsYLYDHUDmDTn59jrWaIVEBlG9x
PAaZf7xvfBGxSbx/GqiNkxb+TvKUIBPneHWGsMmEM3Kxc/JK9+Dy1/eVrt+bQ1g8WjNfF2GqPNkc
aLYhjsEd3WdiITt36lrdv9h+xOh9WtT56CW4ZGidBx6snrwudW3r2eFQl3hUTtj5dMBjVB3Rx7q7
cibrRrmFWP2KhO9V109LNVt8Nc5vCflCCz/1t2xjfBtzrrQ8p3/YU2jbrG2BsPDLTTGfOdzsFM77
06lgM3v4s8nwMv6yrclyAJIZ6x+jsr/QLj14U4SdY20Etb1xne/pI55EE41H+t8IQlGxjpD3UOJh
i15AZReZdfAcXryH5ncUbHbOGW6pd97SqidHWfI65PI0o0j4/p2022PmAT9ro+qcODcimdo+QTGF
ztrrmg2DLv4HZYsPIzBrhPDmJaL6R93mCejmJDtklKC4kO1UmZ+elIEbB4coGhLHxKtYHLfGSGpf
vWXlEuTspyl6nYEHs65g43Hnw7iOKr+stzeFy+ZuFFEbTQiFHbuwgjoEmPgJEUTbIOgSPoSbKlNo
fqLo1Z2qXrXEH4wqsRJLv24cUZDoudWlxbzEUPimIuKP5inTHyKBNtu0Gwv3syBZuvMbC1LCCZCI
bbEkrF5hlb7FHpgXYHiFUkZnSKASDW1oAJdk14wSLaz1kWGh63ileWn6z/V97rVPnIHRzsB+e5b9
iv/rUWuR1oc06JseIwRQ3uIpYiG7qn5znquBWqm396SkvO8eWnZi4Mo24G4whEAbChduSFW37DKr
Fm5+8hTcI0wnAFlveTyCDFKwXGxcI+MYKw5qCdO/uU+73g1V5a0GDxW4QotFGjhMy8fc4ITahJE0
k3m/EYbT0+40kyrs6hVNqmLAgK8LXWSkVk+KMH3YPqrgYT6YUK8SSnQzwmqTO9dBmfdc/orAwknt
UPw2t1ihNe7Yn5n1rLoyIQWQYXuyxEMAbWnTTPhyHSI2tknHXU6bXBxTF69RyE1GzKYf0cSFSODh
YGfwrm3aGMM4ljAxp8gSrw8PmISj5lm6VU7Zekbm4XGJPsS/V+xN17EGxjwKBSALgWgZ3Xg/dSwS
VJXR5A1jfmRWxMiyR+93QHEyiTy2zqxAPhIjleV5Qpx8JYNIOF61Z9OemfK7P0Ni3JIdEuc71lH7
7dEjLFYkZqU8jKLtG9x3dclERjNX+AhkRjuWIKSUBIfEYYnVqTYj52dT7t2y3DijOxOYVyTQtGDR
rte9mGMj6RiyxKLEUlbbqJfeS0Ws+3fA5bnqP7VahhSVEPhSS52cgo1OjuoomcGF50tUHkHIn7Q2
tTagqTxvZ/vEB0dKjbh9+YdIAXtc68qmL9i8lTUAItstYggzdOz4/lvHhrl8zT/55wijEonVfA3K
w5Qugy5Buhy02PtoFIn1aaFwTzZpw8HeQ6bNFv9fhCXPteQIHty2aOc5Wd3TpvPHF90+A2kLC+Ea
yf2j8No0EpBtXgtk6K0GeaflkXSJ2aQDY89qnwF/jr8rRJ4UnDx0Wh/vODL/hTthI9kxex6SBqDf
2HenqfIhnvZqX73v6Czozb/OHT40JzrCJXJ8kZy77Gtqk8StrENFcrgyS/iJhw9OQKa92SmiZI1I
sIij/e3iP3g6rzk/OnNn4DDK3N9EGT9Gwl40WQL+0BYueioomZLzI0mjhBF4aTBbXTeolcnqdWYF
SpKxWodBpLeA3nCzFyODZ06XFTqiEcbc3MU2aZPn38pGckOsKv/bYLMW02MCXbMb3x22mOyoEIyA
VMXYy2iLEcfgYs+5o32cUrxA96VoVuFEfOVor2gEqUOV4zS+E62jaaXcwepzeVNvggZzF3SJVdP5
x1FNVq+/WpxNxfF6NKsN3gBucllotmEtZ2IHtQzwMa3RQQfW2F3PiiO+Q8LFc02kCMLjhflaimfu
2XuBWF203rV4LFz6Yd1SRZjce3xGXcoi1UjI4XiA/LSBRvGQvCUmc52TRayXfXaJTf5384j8EmS3
Q9hEaZl1cOYmvRxKKxGR82/DmPj4Fpo7ozio7iw/BcS1nivP0C9VsR9rZHGS3hW2vYO4Wz7foqQZ
2/D4nxt9LE96EUGXcBRQFaT/l/TjvAlhcLzuTdozQJ/o017p/v4rZCdrdWouJgsovU5Gnf60odRX
AITnvg0pp1PCfq/FrVnAUqANsH1Tloaipa62uPvcj9AWm76apkeeuG2iemw+ADGOedWo1rSFdi3A
mGfWPAcztXfFUn0Q4nmsVs+xFonRgoWToNQyMiNlQ6RHzjfwfR0bscF+I8rdimQKe/LsWWkqPJoC
ussG4dI4+dkc1oapgrzDSDzm/E0TbTQukW+fxBw78cHL5MyCuilshqEIExMc2LXLuWR5P8ZFUmyk
gUG7H5faa+ZC3K+/A6cTGK1yWX0vzNCOjgRVR0sA5ojFAw//ZJU+lSJXmUA/5S0B8R/d2UUHHiY+
rUSMPrrmwLzyXblfo0oyxP3mjp4oXlhiCn0msXH1+/yf2M743PzAkf8qFPSmJj0Q9ajvH+cKehyH
BwHyFzJQ6yQY3FlUKFPcW+CxI+u1AEf3OmMocX9ts10MY1sMd7dxV8bAyvn88uj9/TiP7taYkQmM
Q5Fu/u2DUufdCZczlk5ZvcxvxuV9oJ6wotxLRu1vugaepn5b2pJfzj0PZtfEG7edKeAQlErfy9yQ
rpm/xTDp0814IIww/vBOTBKGMXhQ8lGFBDwP02LW41kaWnFZl92fF1oavXszj9dZxuShAKv3/pv5
U2rHR8uceYnoorvx0WETbfCnOT+dpf/dMl+Xt/YWy/oKrbcCqrC3FTram+H9ft5FCNb9pq6tY8NC
jgQB4r+V8UJcBG334V4got6JNbjOo8ag8WjD1Jl5jN9uf1EDhxoPhbAv6fUNNSdciX4yHm+hq0SE
aMXeNZtaz+xhKAOjEf1QYe02I4IgCOOqa2GtDQ3AYsFc5n4umJc2QjCWYSSgmxb/d26jTrwOaUB+
yszed6/uwPdXWFN1nHcEHTKs9X+dJRy+wUv8WbwIlBmyEL87dmEGJW1vLc2h1Rc7pCKpcVbrYVcn
HgWr1Pk5ZBxzecS3SovvkfBIk7ekDWua0OZvF1stVZGoa/Dh1G3MGiqmO6mvGZjIZQ1W07W5HbWt
i5aKA3RuX5cntqWawg40dd9KX1hasoA2OHs2vn3T6a/Sq51jbL8/NemS2qgLZ1WOtP0Yr4cWQnrp
Awo4T7HfKDVKINMDI95VWH/vdtfT8IrQWcLLWvgU7sBPOqS9ccLwdDX8TQ6/VnVT+JdkRnXqchf6
2u8Xx6JIuPiQbf4cugtTBwH8rgk2TtesmNirV4rB1v4MzK6QQ77rpafC1wGAkFQD5fRAJbcvBd+D
Y+vcC+Epl3NvbUXi9rrpHjZYwjzH7nKFGbYqHW2VJeP0xwPBahqwPQwJx5Fq8yuqsZPYj+7pE1QN
mU6i24M0ZWeUaWWiws8KV9oodY9oMSe8dR/Pe7te8wf2VVxrvTuIxY+jco0DHARyLbYUgrdI58IZ
1fuZXss0nuIDUO1joz6O27zrzSTSxUe+XF6P3JfhQ26lJsrCUy7zq7uPx/DPt6VDuUR4Y6yLc/US
AeZDamUWgyKuDw8goqPoud4M5yS7SucFpTdhweA8GOpYOidSkcpvYcJ7SFQaizKTui2lqL9YXO3K
IjYh33rw4tmRU3+ep44EKfK4liRM/SbnD5iGS1iIM2UdGOq2Zp4g1DPYUxuLXbAvut8T+nfnuydV
0W+WKEhTIFRB4E4HHbnECF2oaPX28qVcD9u3eUPviW+unobTJ9RSk9pazCv7GHn+eP7ryHytTQgA
Uu0+La7FCAaPCLsivKr01zxQenqRhcvEZCTCHKyLE6zOwz/vpD3sBvx5tjtKqQjQEFTTH/L4hUF0
rb/BPKZOLho74r/TutaxQjEFp0byUEVUDM8Vi0+shZEFKUwZey80j7bAkMnSrSVDhYMx6MbvJNND
95xkmX2pphwG2tb4NhtBIj8d/sC3w2dEwnZKQyQMWpAD75ahfN/hq5C4LRT7Xo7dC5MO/fvCPBAg
ee5VLvRPfGPr/Aj62XQVKSuFY4UR6hNldRqxexv/MjAM45QWjJp1NnbsXkq9euWH+VLRQMxVXRkw
INeiaSHyVNqVHXTF7LTkKgaFWNWsp+/tdGjcLKOy4d1FjAo6LxhaXyOqZc+eYcIZpYYog1cuLMX3
oqmQZN+sv+gVNAy51iy4t2Z4KCYM/s5kbnlQZFVabZV6rZu0cCKWb3XsGQlebYTlwNmddAUfmfs3
N3W1eH63PALUyGh8ZfL8HTBCFnLlRgw7ik0ca6v0+DE/WMEtmLGihz3JxgYWmO+4E4ZHVJeR7kbd
YNRM7x/9ovbglIVwos1/3OFWKUVHjoRGkBV3Gvi7MHn0Re96jQtcv7p5soKjkmsqhvJ7OQneT3jv
/ehxkc3ONr1+DKFTH7NyFUjvXveFTzmRPTl4guEA+uW8cJ1u574yw7Lse7acK1gQYj0XXY0FqFNT
VWlAsHiwKJnu5AvlQQUjptHL5CL9RzdF9/5D1BGSto9gJ7BFBQkk70LnOH3VXRqMROkj153xvojs
hqCKkVh0niKC0IQ/b7a9T3BbQfZVbn9X5kn0ezNTq1PQhrg+rpmhzG27hmyK3y1PPjueX2Zspyqr
3GkcW3nyR1EyIYZ63Qvx8aCsjmwAgJWrwL7bIE3SRk/55TGd2pCmzXmitsMCkWDGvTaxLfyKR//O
24G40VYFaq8eMj+i4KDUbeyd/d1Jw2KayEpZqTBuejqRSmPi4ziXTkmzqPDUR3pkPfJioPkYeDLP
lAC0PfysXKzet1DfQ+j2WdN6e2CuSZG3W9+n722GlgzPBwgK+GdahNFSVLzpXBxcHUNyG0CS4SNs
DM4frWI40pE/UVKtlfC74RadhLjckXo9K7usfHZnNLCiuq5d4n0uD0g3dofDemM9gN8Le+yoxwJL
Z8wTZ3KGkaJeFi9lebxeXbFsnYTy+cpCzGXJCD0pF62B1ZyZbo8cyBChpxOqdMGGySnKzMDtBD+B
0ViiUFXLAW+4WFeUnzdpvujHUaB5Afnc+oj8ROEmR98590blk2zjgdGUjH4XKleZJvgS23PsuoaM
SBU3xM2wDirP4mgskzVz0XJ7lsDsX/EiltWwRNsC5Eg2j8li9nwp5mFxMYqGI5XkthCsaWJpYd9n
5cus7geAff1roIF65uBSSyGW+zh9eGiBQ2h0ijCAHIg2l3tQdaZf+jkDUCfMBmgTefS4bATJ1Vc2
A+XYfDUGHeBv7dDLOeB4W1FTyy8VTSVln6qGlZK03CPMSoC3+++OR1brbKfjtOFaez0adjg2XYhZ
ioReAUBieYn/VqtESTwsUK3CZ58TOcbwetUds3YXN5fi6vXxWR7pbZ208epmXMKiuGfVkFYxR+Fx
kc4Mb9MeYbNR3hpibaO2JoRk5p6tzD2sBI4Tm5ax0s+jTtwR3H7RyQshfyBtLMIJpzPTDlLEJTx9
dADlvsFKO4pkSuhFedlzwITjMP4iss+VL4XujM+TQ0YHUBnIferqY4neEzqTcocZ3va3z2CqTr+3
3eSKi8UEQYNlkDeSAHk2pWv/ccKn2kz3j//gZwpFwU1YdjQVteMmq/ki0R0rEBeT/WQNHIuQr2rq
V9sRbg1eb7KwvB5rL6e/afiwTQA0VxFfPBuHNpViwkBwIOthh8iAV7yF9N1KZ9uajON8xSGH7sL6
7mLu5HDziTtbiIAfWgsKxQtyam6lbTLfGBTYoevsarc6uoVmrYqNsULxQwMlG17YC/yZwIiHki0Z
zTIctJger9iKOKmw+X8UzR3Fu9QQusP8C8OwgSSlc2jtaxH1i12VPlg+s7BLJVv3ZpuhXvYqLcej
pUatpviXwock5/y1PIkw1X5eUDkZFppLQRvYMcABI6Lfy1cK+BqTP4EZS2juw/pezMGVMs+V8h4a
GJxhjF3CB3H5gfs1Y1DObcMPBl20AI+L4pD3iGV67mAZI+CGuI9klIib+Qm9dSmsrwNWXNYV/5ls
m12kOUkH/AKxIbSBdDv5DeDc0o728088NeJ1cCGiGfKpHOEUj8gwwnFOeG3psWEYHC/O926Tqxr5
bCtsh7M4dDx3Lozu24VTFM8cgG1jt8BWdow+ww4t2IKlIHAdGtpATql7xe+clTTy6Vp4pJyCAZ+d
cgzpqps9pxGmM+puFfBPcsX2CzdQ9x5rEtilIqN0gNr+sfwG/+7BAJDhOc61MhffWJJuExn0yNV4
+o3e6QUTyBPPCMIKKyxtRMC5vGCduPE6U0DwWYb2iKbVDjg6dx1obw7GqdXAkTgNhuPb/NnEJ4Vz
Dpaa1bWcRK5FKxc2zCxDaxhMgd/ZdkI5b1gvDZR0kyIffevdOE5CJDQJjNKMwlv6nE8PWP7SOwGt
HciuFgtnZ4Cjx2Z7aYw1x9Gnd4KcLiXpPEc8Kk4BmjJrTagcD5wMH1VnkHIt5LbO03QR+uclmQxp
tS9OnFeP3kvbNRNyIbNgUhXwsVbOoOBZrNrHkkRos3bL8/19/JUMC7zQmTklK6p+x/JxhVM2c2hQ
4b6VZlC/s3BRhYOyziIAokXrl5FaGqimGxZkAeafBg/kfFy4gtucWqGFRWmlpbUfsmWYQCDVgnus
qWmdFK2vqaRmY4tXNez9e8BtjDHhNwM9DnuanzY5lYK0NJrj/neaqXktHCb5Z+ycgKdcXG0y/MDv
2OxQdyZ4MURckdcJLxEclQ1VbCcBnkHE9+Y3OrYqMqYC1PJyAWiA6jGfIFhPCYwugP2jRp7BRgFG
PZoRWw9pOYHUmEgPrEEuzYKEVmYTB0WbVw6wDJS2vLViPyY2TurIohWQnP0IpXKnBZ5qdE52WCfO
wu4A+Km4PoChzJ5+RfanW8/QriiGxjJsqQkRY+kkKbLk4An7pkp3wjYXuZ1HC2JDn3DG3WFf4XjQ
kgoNu6nMOHXSJn68+e3dKmK6MX2qobKDfNGoCAONGQUTjFdc5KS2cu0kcjCCX0nyX5yYcWXR4Yg+
yUahXdyI5m6GCdOgyJWy2GhSgPB2pzVMtcfQ0asc/CmF/tT9zCq82VvpifnbtkuZOMes5mryjCzn
NbU47fe8bjFIX8PF3FujFS1IAXPHUaRdxVprBdlMp0nwNsXTJFK+fumjChQklzt7Al/5TsQO771w
O4A0Nc8EH+Z3VHRjXBytCVHOqdi8GZANTNIXD2mBhjKtLiWkJlSqb3PC+q+o75Dqc2hnBtCjiPHM
WkkpMGp3SWC8XMk4XJm00ivHz45UxovP2uaayRB90sfxs4ufb8L/zDrjMjv52OAH8exJnf4d4MOW
SxUcEFG7kxphOTN60X7UJcIGS9OAAwFiXxBJwttSbCoU2Q0JQ4QBI4np4XJ+ecsA7SDu1QY1tFHG
O6d2h/eiMVdDlLDul/KO70hDGCc9C1NjzoZi+c6AlbJ/NcS9cNLByX/o+oNA7oDOZeelbW3GNDed
lexGHLs0StqRvrT61RPVqMm/T14QDZfeDQpFyw2nBKyeVgBp2wDejg47Rknu0FiBDMm4ORKZ64Wm
9h9k9I2VoMnOHZlRjOwBeWLEoCWoCV3+vpd0I/SMrBBNwUyIpSb/4l63eqvOw99tQXmk9mtd05wO
0ns0Ro9FT/Kxz7/popsHDGqIldfTcbut+6srRQPLn4QjA+GzoY6JBfbspFoFtbzPtqhfIYvioIx7
FHY7aK2+ajy4SUpmcIPlNOPqwRP9s49h1tYfAQaLJGxtQy6y7568/g4EOQTU1p0nLy3LGtRkb8XC
ZkrnTbMT7uhRbDNZ/WnYGZLie+dc9PCYwbrgr3C/bIIYcVE1LFQEKtgwbcPj0FYFX+ugwKUmUXuu
p5WlVKg1vYC9ogus8P1JPkKPWW7CAU2nXuDqpG5TqV07oHwsqkRmTBj3nLXdFOk/GKDitoY38e39
PCsXthST8BN3TdaLIN25bkQuiVEw7Ur1n90v+t2vPjlcSNH5pruyExRYlXDut1KWuVPEtO22SJlq
pwCVt8yqB9CQZO+gu+YQKQ2ttVFYcM0Gmy9DiciG4hOu3C6BuOCnIX0HCd0mwbnxlbpxLPRH2g6a
qTYihq6AOlk5Eboct1FdYIebRHGQUZtdMVNSg5Bq/8aMjpvl9NRidXhJod6yBmcZ6jlxZQPXP6+C
lrUitMW2/j7zP74LCOCBWw2oHzQGu/LREDjDqtse5JH8jFx7qrAhev/DYW129wJ8honYONW+aSVn
2hFhKagFutd/KDOFFGRhi5y//QLqKsBmUvxQ0uvEG0nH6pw6KC9kLKpJJTgMv5yNw7BLqkXTx0Hr
IrspfwoWCIGn+m5SgSgvBHiNz5QTkvt/t/EIc/EySWghDLegC8d9OiQTN+S3ZgiGPQpTUtf2AY+a
MiXXUMFNK66VRQC3s8dSAIThpV47bxIJRXZGiCnRLBgh0DmFrKLaAeiwkhAcpTMBYzH3Y91i/E3A
rsC2HbNjLKbprM17/VVNwkikuMT8dpKC8QPzx75zgZ3ju08qku31wKGuXslKXYFzm37520tzqob5
yFl6g/iBEfWiBXgfmql/gvz1LFcja08DT7Oj0E4hUL8NWF6saPx8vh7+mgQegT3uv4cj2zsvbZPD
hUH1e4qrQbdUGOxjcNE5RO3C6hAgqhkG8+mefeea09cICtWrj7OaE0RF1utro5mwzebHgGvGWmTI
l+ftJbT7umSL+itAxOuZ0SLoVWQXxPfTdT3XuCay7Beq3tnlJPEkCzV4p4bQjARYouwk5BcAi1UR
m6w6HvTlmmrm/Qp8WGxTWhcJ2EB5Hsxk7LcddNNHRaV7fZC4DcWnZjvq1Xx9/gVf0+/IzSaw4SGU
w5zNxHLlEB7W3MiHHk4LfUDucCv4OkY1td5QLLk4i8K9NppWpkN8MjxkXZpPrkxUWj3Nj4u7xTKM
07TxK118WLUInPf0gSDoeaJhms6tcQvdgkYcljhzOahRcD1S3PqsjIoEZ029L3AMMM0P9Gd/oMb6
Ir5k6K/7aPu0gJ1WV8Hb6C3rVpmbHsGoa9lmwNxjpSPlq3BU68bEOhS5xEx/MU9xU4SIJS28UYVJ
WGkd+O5xirx9ZnDd0v0xxy7R3+YaZav+Uo4HPZT2olOUDYXUrtPf2HLIs9kC1y1xGUEyvntOhiS4
9APZkT7u0S0+glyL7I7fjJ/H6JIwPi00z0VHm9UYkbQfQ6FA+sjQ0ioIxC67xYDiA/D5RMIL9t53
qb4qN1gNQew+ae6hSJ6k6lVGC/DwBZewZNnJx6dPHwI6rHknLWXMomK6pNaDOr2bRFj+K/9JLpMJ
PjYbaocTHKyDJSN7qUHsJEjRgjBzuv41QTT7ky/4334VN9rCZikD/e5+wDZmfoS3fH1eTrgpD4yC
w6WXhhTGeM7OFyLtwQXkLO7rUOR5TssNDCitHy4iGUuGtN73EhHIk27lN5CZFRNSSENYgYJ5cJ21
5VqMKzr2wAmU/RSaZmI8s+NJzFTSO1GlTNqSnsksztpJPNvPAoGTC8YXVNRe8CsLzIHuATYqu7Bj
B1ZWqVAgA4JaxOO6Tv2DAMCZlWSna1/d4Ye8A/e4hJTchNONdtsD/GYlXxwfXb2ed0dbKGlpMyFl
0RohXCqoX44UuWK7JIqDVNK3RSKgWEjQRBbtpIRQMOIMqE53A1c+zopi8nQD7Y4CM/AfeBARL14f
8us13b6nUelv8hsYcoU+ND+S/ERlf9whq54d6zk4LebT5K4T3qsNmhalwlrv/q+2Gy6wQVf4a1+I
FaFWWf7UOCI1zvRQWqHxT2ALt1toGeWL0vEk4ApjYTWheD6mwC8hkCGSGRRAzlY/yD8ta/Dt08ed
g7FkLs7vDctHQ5hfOvIWzgmnwm07DSwG6efHYP/LycpNmgZ6PX7W4gXenG3PuT7kFcCP4MAd9eFL
0LDaO8KmGCCIEJbwiN1gFo68GWbYk3h0SVikgtF6YNP6WrygzxkPYFsN5xlWig6BqY1yaXq19nTv
tsEkRFLdlxpILsh9xkzJhVb7xS5sEV/5OFGhGz6W0Zp1JWlrjRdJPOPe17CHWA8FKAWXw/zGRPuY
WlcWfR6ZR7TTic3WBbpOCZSJnMHGX++mKlobQfVt1eVjly1YIT/aeOyt5L9fMjazDk+vGrpPP75n
09RkYHfBXm/yrsVomN/NNWXvIb5YO561+kuIffKoyoMysZD1V204M0mh1nQKSsgPg8GD+ns8kAux
pwtx/n+SPhSaMp8Z8e6TL3LiFue+wAMCmY9REzEElhV5Zzl6B8yP1zPukVmu9/9DedomDx6hjoCk
GkoLIdSIjpJLCkRRByLH1dyaWhOxC5W/eBkjVEbQEEo196lCHaYLVxCmaGj8dgT5krsgOcXaBSnB
y62IP7odOaERaCU74bI+IjehD0PVgRac8nr7JKkjRysv7dhPTSpS7m1zz6zeesYaHIVCEgZRyTtv
xiOu+p3g7lpIFtBjSGwlQxPa2X+JojyrHtasCzhflsXrdnAdSQt8+cTbs8ocGl9OFZvAN2eVfY6D
ayLDMKhys4QH4lBiXh1Nw4ZgippryxdfMYlYvj4c9Ma25fnf8gjccmVQLOqX+O7LCj6NejvuvLly
u4sEAY5bWtaGbxxYWC9LGF0WEx+VNPzUmOg4E1BT4VhcUTRoJ7Dy7O6kjJvKpIFvjbLbhJJ9lmv8
EbqmutZ26bYOW479IbGFmAFWccYfX8zTDF5LVxJ6OubSArCkGh85B8Gn4hqNskWltM4+mP7yrgeh
0YIQb2VXGx2/1lgls8H/aYYnWT16+KjqnQGQwyWpBkVSO9/Wefk+9vrAtJXDqu/7nmwNlU14a+dL
CInYfEjpE6Dt61ndGk5IGMOymNS44iUXiRjkfz9/rDcqn5k573J6d7l4bI/0D+2QIVQ4GaZfvZi4
QaYfnxZEdPgMQd8+RrqO37siMPWZ6Al7saFogtQNMMWyxe/h1R+gSncxRY9BWhMjMrJlMhp8VFvX
orwkBlzHVhfjE+/Surf+Ih3FPL0YOpDIWAfnzRQdXNfQa5E1L5I3ffnTVnd7/9haMY/5OI6PX3zT
E2yfChmB3TiUC1EouiKkhJJIPAgHwyF7LRa4jsdi/Tb9cAp0pADklksGyn+3wWpvYTycCsJd5y63
rEZaHTKYklTx4X3XTgiB79f+fZxD5E4lztBN40ephbn/P2gtiN2pKD2pxkF+DkaTdzYn56GM6nhV
r1cLNJE2VMn0ZrDxg4OZJC6ZED1RcCjKWfWjFSp0wQ6or1gdjTqyYbeUUrd19kchTWOFgOYgsO/1
Jn+XCQ7zLLxYP6v9Hmq2gpKycBYB9oJolWFf+AiAeXNauaBEAC8nyMCAM76fscUKitJoE38kHW6A
ud9zVkg6uNNOiQoYADtRlY/oyVY8HRMMSjyvAv6Ny91yPl/5UO8dvfWdlKpC+OxT+hQOxiw6Tpx5
8iOrr8ZzXkW1MaJXJGQUG+Q9tu6lAGM9418wWqnDcQ6R1ug+0UZO9NnqB0fWFlYj77r4E6HOqp1+
Wqzcj0DOSSIBCMLFSwwNvfCmAh3dRJQGOHQiJuCa9TFKWLIu9XhAEmk29B15vrfD3ZLuWmgbC/RD
wx37j98lwOv2K7VoEg55AOq1EjUhuo8Uah7dGvgvHHTj02xT30As00FxHjZsQy0K1rULb2L9RTlx
WK7SA4QKksRq40VY3Ni5fYAMFr5ozCTSo70fdn9fFTrLTUB/TZLZaydeQLXcCO3U4kBzqrAv3L8r
pddMuCPUxj7XJfHsyzzQlv4sB99Uk//liQGXscvGWpo+kN/2DWNoiH+S6v5GMH1WfyKSfp9xQhiw
c5ZNa/XUdXXQakz1i/Ri+9pHRhqNhZYcz0N2eJbLQ0q9mirSx8bvYBSg0yfauw75drcEZv6KVBwu
b/6N3ZHj4LErnhLr30nYLabh/4iEzyJyZe+HEzf70hlnHbMobWFiZp/Jb39QKDE+LmNNTxxO15u5
I56ZUt1plbgrvscq5rYeTAhrxCtm/8EeIRTajA8HYDr0I6KwcKgBHv3qkubkF7SxgOkCYy1tpZBY
840xaSw+g1VnEl87nzmNNsrfg2hM/aI3FVptXDpLUbOSKYeA0FgMT4zReCYckQXBWkWdvAILBlnz
ypEj6U6a5D4QsE9Rx+8r/Ek3cDYWU+Qg/pwYOwEfEDMuS5NWVOjZ6WkwwonbhicxLy2GUqL30GbG
tRov7C9Xz+v+3v5iY99WSlJ0+m+qmekVYgIS4ax4HgMOEHVFEqSZjL/Mn0aANuNK8lpEYSNWGzIW
lE9qXAK3KBPKWTsyFiJpfe2Uzmrl8O9RCyK4XBifpBJhFu7eD2usrcQOwJTsKLErLL12rril8xSd
wdfJvO55DczkMXjgZnNbTexgcZmSowmYU/bslz865nvngWdiiPMbZTCWao4x1V54K/PmfLwPqJNa
SroLADjk/AZklRG5J9l1OL8GeAbT2iMyEhMEXtZVf9w6LhWtKkrMIj0M4+1pq7H6ISlARKyUbo/+
xTVU1b32qFcrBENen57Jv1lV45CYt0yXcIpUy64m7eDyIK27BEHhMqYEC83kmIC6M9WAd97ZYwJi
J+8kAoPYXTyKGItRMQFQ6swE6zWhWvpVEOsvYaC7+PHyXQplQcuki67lhiIAKmZ9XacOjsjWMfBE
FVPsZOXSjy2ypYN20DVyAkNWtsP1rK+0OcI0cXDB1xT8C0aTnJtQ58/EP9Iivcw6cGSJGJg8k5RX
IShOkriggFiHRDgC81WcPIL0lWWjnqsbVOrGD4ChYjQ0GyOb8ciWl/lDFz8QuDj+oSB+a42uzDzJ
rvkQAT9sQS2grReKGIbDtFmLWtKuF4MEypt8FXXoVonXbJTmMaGALU9wDL4yg+/dW+fK0ij3DzKl
CqS0eVMln7N1N4o0rUYjaOWDEQV2+rJIVsyoJwhTt/+aSvdsYOfifmlrJXPPEdkcRR2Ss7ABlPfB
FY+KVOWEgRGR/kHHpJ1j4iIOir0TL1IUQdNT1YYgfhDQi4gLjwf4AVW57Rr7jucfKJvXI11Zxji5
3chIt5uJ3rHe2z0LuzisvsWuxSgU3Dan13HO7NQKKXJQBWBLC5ZtrANhtBk5Bm7YWXiD7Mz4AMO2
tW7BZB2pecf9bG9K0nrn5AjFaEvlz1DqlLXm/loy9u3RqIp0kNYjxG8bMhnjm7lA67c4WB9G8Dp6
hSOHGFNnITdD4JLM4JR614CXmjFCVR7V7A4SqRRXvL3i1+Pn7Im13vrlPKBFDJY6jqwWzboSjpiq
ExQM+TNfEFtahNsmjSlkWNF0Nb2GovmWr+SpwFSAAY39qE3mQOEHDiPVXGc6rxsrcqJaetKPoQTs
fLgqI4zuTPqqOgfUdu9qr+YY5Q7eW5OqFax8tc5sZnAWofYH8/CJRP9rkoz9otaZKrkai8J7wH+u
DXs2TACt+YPVMLCCJe3KAO5J6hCmeluNb17RNyx8FpwRdfUVGfDa69npPYkFJ2qpqtGLKzv4D+ah
WW6BY1hHAj8DYloVwDRZhe/tK7Ojd35mMotgN4+0TDQRZx9pzEfGgDRaiQ5pr5SqLHwptarqvH0v
ksXdfouzHi7mi9X3qMVHe1Nt6HtFeIzhdgLenLRx0Np5wzMO1JA9rEl9UG3yT5WeRCTSAH1w/zaT
UV1cuu38Y3o8USbkIBpbEq1VvaBxoEcUJjFi3/IuVB9bYqNrbmxYrBaO8jeU8fq5vcUqcDYeyxZP
NJtiQb69DpsFa0u4Fk9j4+9LjnA0cn1ZGHLyP88iyDnPIMrFaeJ/dkFzdQc64A/rhNzgrinbl5vo
16hxX0kL5VjR0eUiNTwIGDEyZJUdBuVdkO9NGE9gr4Ze0CQk8hUjq/mv+fT0OY8il/Mpb41fj/V2
sPFWTNQAuVFoZPzcpECMq2JnYe0GLaExL5tCQEnlMb73OK2ZwCIafQSq/hXNlYW2430eX/u/kZfS
o3hc7fFHtTbGmUCytZ2GxO4MUwV2DuP2/bOrHeIXwogmIEaEhTdyuACS1nV0HzLJ0XJYLsVt3UlN
pLQAx8yUT98ZU1nJtIXJvozRiMAlEqP5C40/skA8FnV17tlOX8mQ1LzUqRxc0PsLY84CZIFETyUU
ACkr/ktuloAnRINQjLZRWTvHxD+2X67/nsHx6N0OwpmSPQVvvRkrLByIAqnpSTb93iJZEt/MHWIN
rfUXW8eQ0LnmNLt9XTKvnga5B0ijZSOrPGG1uv7scLI3CKbIRnjbcqHEM9gcLYNImJe3C8DwSKRf
3+JDzayYXcxFW/u0tnvkrxNMYPOCqGNqZPTaKY8U20U7HIgqvqS5zvrN8tItK0smY9vIMwqFKzJI
P0ZfyLUw8rlL1fmWL8EC8MiXrGLvjWYX7DJbyNDlBsU5POzp2OxFGibrvPLjuBMRe9fsijfRtgQg
l7d0ClN5/sjgIkiprSm/vhPdviUeUnDdqnfz9RGfhusrrs5qL3kQQYF5qd56Z0yNJECRSKTJJfUv
VGbElcYulFDZglOKZEOqz9MPa+a2qtIp6rAgfcBJdCmUQAlclQiWMJVQx/s8s/C/kKGdns9I50r/
H3n9B+pMESNDhVk5RVVqYNPO5hH803ITut5QXHiR3QHm39+xy97/4R3lusmy51MJZUcMaK7+mDds
VMEVMPcEK9EIcZbZpqhiMNA/ndJpfbqn2K6FGuORqfPKwoWLN+AyM4mTrBpXMo8abOxOcJDfFKLh
noCpSv91KK2qUMDkQnyGdNnfUeAXL6KDvQtoB/Q1RfC3+fM6gqZrEFgf+UYI6xWC1SsrF5kEaStM
aHO4y7mj5CTN3Z2jwoDZxBqR/rpWxR85s+4bHp7t2e1hz7z6GCuHgCfvLFSnqQFKnhoag47w81uF
Jke/iX2VOYHIdeeXMFn7geiEqPHVl+FYgDkSoilvtIyZF5mUKsiKYB4uQB4yvycBpOHbI7sDub9B
O2uUG2jICmyvUYRKbgjVcROIZFLKKs3rJ6Wrhp+Hc5w+H8D177+mJ0Yfgw2Bx8iROx3KIW1D8xnn
Z8a26RNdbVj2gJTnWbBzl0TH0mXWzmm0/X0s7h3mKDL57T5Jq2xcbynhePnUspOj0hHqg46yRuxC
XJFPzTZZ4eqznY4DOZvZjl8rIgipXslveFz/ah+6/tnVYr2Xl9/i8F6dMtGewDYujsE6jy3o3Fl0
qlJpcTK9sfkSv6XM+UQ9INmFNF/sT4pNGp+sGEpSfhZVbIxD4zDeNxQbvqfhpqKeJ8QCLLPJMU6w
qTTvZCB1hFQjbuCUCRthLQHjWnBT2dVr+n7s/6b6Ra/n9phEdNPnJEgW6YdXQc1/qAqg/ZqsbZvM
+gJnh12bGumVOL9nHzeoda4iproh2yI8vzvMu+HU3r3FZ0232J5rF7TlNOejVswM+G0AcWQmIDsV
0uh3QPMsnQlwwAnBvl+l3vbtgtd3vd/OPB0lWwMGcpfPw+LKyB2MVDgUXBq+MLhtXaq8DrFJQ2eJ
7LBWnOlflkHxfsgR18L0fTIH6fJFPdgvKLWWiHOHdtEm0Q1JkBZBBOVhjALUgRVBR3J8NxWZz/Hd
1EIDXDofoKQp28YYYoLf2hHV3gfpNgHNY1N5uPG5NBhp5SieqEX472n/1Jp+fH4XpJdVSbCMMY8P
j4uKgOVzOH1LTBMP4RcN2X+/jUAKcpP+61+paoYFNCGWtDKPe0pZZI0gQMH3iKn3fSkWot+NnXgo
OjRVR6lVTlbK0xSTpMGBi9pwsY3K07hH1jKypuxiyS/lZ3CL56EoOHZvUO5VD41D53W5mGo+JCHX
AG+raOPcioYfWlqBI0dTi0sZLUUgtyCZNGDjQrRPtwdcynqxFipdsL9XvtwRWRhAy+M5t7tgMs3I
XW22fvWfgAQUbPiduslOHrOnLkHdKF334Eorhs5rshCK3bGq7Qmnx4BbELau4ZOG/01Ft6QLnwrs
g46jMpIyG7q6awoByOQiIIHmPNNN/IscfztOYR+SPyHZn3UBCR13b1IaPR79yG8IVbckj9Sv0OLV
e380zMP326oeIB6nAWl/OnuqAUD+Nv28erMIpKbTtVcDzEt0O97s8hKXfqSke0K7JrRDBBeF77op
/NI9hAZ7YlXOKg62sMmOPhbjhXIkeoGvxhGuRMOuzarn5ihkpxJ1/RnnO6hGT8xBRINapgrLd/cw
ZM3clCzBAs+NWwLix/wgsENPA0JTwDdcNYPNHLvBNWuzNjr9ngxx2VSbgeyl3ryAa4clPYVTBuIr
A362Igz3oNF8JfNOkprmcLwUzFj7krDkTcxWVSahM3EnqwdOLS70lV6Lo21z8uVPtAwbADlAF8mc
nhXvjVP5J9RVLNwvdxBSYE8jRId5urTzz5Ut6QWoZlCa6tMq0SxurLIdiKyaSsgzAx74lG8YLznw
Lgpw46yoyE1MRkQTEXvkvmle+ZsAzcG3o8xTH1Gz4HcYwlJ0mKEb9EK/gSQ++MfZWjq9k4T/RH8m
r17kK5Z5BJL11JnTndfvWUeYwT/4yhv3LS/Pk++T+Z+H/uhzI7BJ7M0OGfTxaduooM5mYzdL4TWR
7gI1i1laoX7sLDduQ8cKN7xHldB34ZCl/kGlRJI5sX2Hg0R962hoV6nhSOYJKQDmAQ8ksoNomOPF
6C2KDWedscUBO16xhD8tA53y+Q7QJeVHsUdZuPLCZ/mU/G8y6TjOT3SLbdNuPesLFQv0m4bQ+ESv
QQ9bt8BvEFJZwD8IwhSG5Bo40fOU5ui1b5WMQn/v1ZCD12D1IAe0WEIb8zSEHVFA042zgBu0YzDt
dZtSyqcplDsllpEVA7tBmTQAJbr09ZJxbIDw0jV3tL/r/j3agnT6qgc2bJ761I2GLRz7/DMRRbSG
cPm+z/zJt4TElPxwgMeBu7KlujYom7kWqzWhpAIvkzSeIkHBh9twgrdKGFdjU14UqpVdQFIPtKP2
c8ypHjqYZhD1rDicAjTsZB2srLprSdn+Id8t38I2IFIKTgcKhiq4pWZUT/BwvDYwsPS616zQjxvj
semjYxRrX1qzdzyGFoIaecNuufB2wQRPlRyhXCQocC97tXCTHWv0JrfZIkF0PRoSiG7dnFmpQHfg
MSU3oBHHuVl4/CnUi5nskbWZ/LhNGwk7DFaAE8WkaBhykcWzdxtq8T3BU09+wDtlX5/sovjWMv5Y
tWQE0nAVrQgYywuxZgcN7mPazRzqacLwSnz7YZqyAWIg6kdo1y2GVYPciR/1QF+J0yBj2F6tdhW6
9FyAWw2B7P1iB2SDFB4DP74G2F64C4e6lmSChgHRkbtO5wtmbKawIjOs9QvlGRhh4bx5+xmGnlX8
kHA2n1+NVr/03jxDDXEuhosytB7n+zZgiGppnSHonBqkqRSTzNxebHFyj3fR1lEFXjvbwcYAAu4I
JrOJyC91PP0DbXBx4IRy4tuo5LMghHp0XcUCd2n9muQ+rjB9C9l5HpynEke31/FNHh5sFFkviwgr
11q3eICy17SFB8nDNRrUqqY6UaKQUtHF36CKjvQdIndglkDPiVKvXJwA5Ca+k8K88ah5MCNjGmM/
aNImT/utiDiSUCl86jmwrDoOb7KZUoJC9XTEluB/u4IbvY687iFyU0fPnTAmkaAji/j/qEjXZxG7
6kO+B3C7oTpcMWK0zgCiWeeDCCUTRecCw7YQzBnuyEbK2bXnYHZZ8R7pn1CWuER1DwrFIwBtYSzN
dd0UDn3yIoEishEzqiq1MNWti9lR7cSZdV2nhsz3/nC8iRD5+ih0+AuH2ZDNkAs0VAgszbvaqAM7
tooQqbsgYy/Z9yLH2r+/S0oho+xlFFWdSofu1CgH5z4LkNNKe+0zhEJJkz/RcPDAIX8OTMJGA3iX
8as/FL1VZW0Jrmleky0ab5sW1FMN88LLQMyeUcO58xisT0AC1M3+z/HvNM5mddAIik//umjrkoRm
QFWaqjz5CwYZ/aWXg0NJeDwcin1kLyffDjJKGQdkMmFjdlEetbRfOqPfgBmoSWT0rmMTSU042rAj
As8xX2hf4XSqBpYaf2GZ2AaHmIhUpDVGlI+6TzKZolRfkLViqE/cz9oRVG2nzBWp5vVgDHSGKVZF
c2txlkqyOsqu4U8XiveltbMOvAqRiFOqKne/jELnDU1WjJXBeGHnK0858haAZvb4z6kY+Ir9Piye
JRPK2g9YIj8E1oZT/ISsAKdclm8db9YW2i4upeH3jiePOJbVAGrkkbXUhFhCexjJ2RvTj3v+FflD
AV3ixny5kS/qbRuRm/z7pZKp5YZXkEHTJIGD1ydjhS+h0kf7o/P9sDZ4dHvf7ikOhJiwmwh/c1AY
mym1r92Drd5ytWyaIWlYbixm6NrSY1dxPhLLwyVfpdbaZaz546oXeIY53u+5NBh2D6s016dWIq3z
OS804k5l/xEcoGBnziBqFK1WnOgL8B+ntTcdN++H0YGo5cfT2QDh29Ru7xA7O1U4JHl+2HTXVhs3
x53b7yL1XQR/XG/IU9gckj3Asw91Egb4sDPszwxi6oJNH6HgQO/AQEZzFQvpm9/W3/48rx0N+uGF
l4ZYkIxdoTEMc3C9oSmz3so71z31jDTCqDeeguUUWX0eOu7vLh380KBx7nv1v8mtI34N0w/WbPCp
gLJZFE411BozVIGNcXXYOLl+nBO680iUAkHi2UeS5rxNkJ38p4t+dm3wa/gYO+aE6iO9J4pnx9Qg
JpFkOhd8Yu1V1o3MoFrbgfg2Cwyj1bLKRusAzywVS+zdf4749ufZrlYqtU8s392dMOus7L4tJA+z
Uppy9iCi7w9nykzZh6rw2DibPnHQjkuv1FLP7Z6HjSeJVhfThIKr9TWVZ9f1CMHOweajY7ygETqJ
C5HgJrk3iEARH1QGAjhk0cEy9JYdq6x/64yf3KTeWjE+c3Aamj3r21YMDweL258gWNPSjJGcDaOD
xK9oWEdHVazOwBFILvrWnvu3IkrbzrOHh5RhLCpdnB3WYRl9xM2wIpOGI+VO6/p2DKe25qOV4pQ4
UwE44mrl27cukq0vN+Duoj2owNnBbhIefNuc4m/xErcPoeTyMsuESQzuTeXDhiWl234SOLUmqo33
WNkX/0j/3f5Xgc50T9tBhfiwPA1ZqSa5jD9ZD7uGQsZwVCpb+tL4hPIxwHQ4aB6dztxD2ROpXhzh
Y+kEpV7ikeZNs7RZseml2/jHydB+mJ211q2Q0YbcYqCX9fUYK4NkKZE8n5WaqrmWqTrQBLRVEAyF
o/gDt1TYOB9zeGvVFTBCuiGOV3Z5mrOWFHCXF4lMJ8GGgQTHvoKszfyZI9wyaOVRlUZ8gyVMbE2G
WI3T5DIV6MS4o2djIONA3zkYKQVhhjWe3k5kJY0FUDpHVzjhlHmT/imtXupkildosudVJ/hq/mom
YHSCDNAc1grL40+ewcWfquTX4wtzdwnOad8SHR+yYdNODmnqonjR0sBEkzMtUen36LbsXWBVPbQ2
VrTtp1yAbd3JWAFZRkaJyt1ryTpjjYY95GAMKp+WjL5GYgkEdp6Aah07i6GnJ6t/RA14xRV3KykV
KIDDZgzTLhWtvgAZYQdyKWHe5U1vGAJx32FVDVoGYhe2VRaieKqzJWW7eehU1ALKluAGsPAmArmW
3kQ9VoenH5V2d4hcfUVnlGpMwTiBvFi7ouLJiFAHgLJAwARI9eNZ82SBlvtPf2FMgbbV6kejYLsb
BHNOg0Mf0fwxnUN4YZ82sIqB+KPQhkgx+avAEYBsdcu+KaBaL3tMCh5fZBsD1DkxkHBBu1kNw4MV
TZVCX6IQR8FrIbw6oxZm3xTMbNxKcZTzAvz8AjpcXaw9BqAPYE3cZ9JXflDvlLN+JV4ygGmlwtoF
1TF9gfTCjCOmRIbED2QaMjCyNi4CKhUKoPZhufZ9VVoA2VsbEt4aajQcGrjS/orI1Ka/bKET1W7t
5FQ3SsVnhcDSnEO2QEsgviftLlWUj0xhJi/gnr0aTS+qUvO0uB9bU1IAJhPTxHECB6wZGE5m8HBR
nSlTj6ClsV64L3bUqrvaK2UmNXaKDrCTX2vkaTAtrg0vJjKdNN2VN+Xl7vWIssVDTsVm/JxXW0kn
8/Za1GZoRcVUQNw3Gl2RQ5/8JMmjI9RPfqZGGRV3bbKrNZSI3p7j0W4eDkPbG+sGs0hcI55OHczx
hLh3XOlyJgW+Eznotjh9DXxmTzR/M9DQ/236XgEDeTVA4Sn+ivVEV9TV5kuwCGGtyZO9V6LAmbOW
+BPytyfQGDuB2M97HnGNoDIOxZqOLVqd6HMDjGsQELm08OOz24thVZSuFCiDOpxk3EmiOWEiLxyC
mvkYPCE6IAE1GvrOL8ZI1zy1OQg0LQ9F120CrRVz9vzEcSDbp1mlbVHp9tyCtNUain0DDNB+XGS4
ErB72SwePWJfEkM4IW7qxBBNPd94Xl+4u9j7WA+hFOtgaNjTsW/m/zmpofvCLDDUFxswBa+f+esL
IF24Nk9o2it14sQ2wJeOox4+U5RLy2SiliW1XNFsbf3/SrwCl4BbJBOVMsIoKK3p69gyYz7dFzun
/pCxBMRszTK2Oa3/uGVEPemNNp/1momw+ubyoaLpaujX7EAXzSqxjEM+kS5OpHpVt5i8RsM9P4mu
/N8Hhv/tb/FDHuasqRFs901YXnnm79mxftvE/xgH4fjMocyyYqvHN4uO6UI/49KlmczaRybi9+ww
0obdluPzLyubYR21o14VVnc6Se4QS26rWKEW1EEh8hAt0y5WX093ZXO44LF4cOtHH6EwxWfSxFvt
4WO4E/YA9/UY1oB8Fh3HkTbi9SvRiHC4dwCQJsyFYJc9wu4K0Ur+OltpHlOjdaKZuxXSybtgmK6D
I1nq721uNMtYnfha/8jZOTQSTvpQ9Sg9vgqYsy/lTEJgM5gdqC3RxfR9E3Pw0nH505xdTyNG3GIa
2Vdw0jdwoqg0REj0xAPhrENhCmkrTP1XRzRh9isLtlQfvVTm3wvA/dVMlEpOJTOVRQQa0Ms9phY3
W3kcyfjfsCv5HfUEpkcf+EgBF1v6ZQbK+/E7P5LdUtJ3M0h1K7k1Em3nAZ/+AAMa5LY+HHM/Ia9Y
oHMkKl8FNO+Kekr6JTT9zWZe6Kykc+Uwnjh5J0Ci6gZx1JdjFhb5Bg51LT5Di/fStjKwYy9Uvzk6
KxuwSs1j334KiQnoafhiiRWQ1PHBE2j9ECklrJDuIwnXCt/kN6rhvhH6S4YZBlYq6BSj8erghKJw
HPSRbmEJ6TEI2hAnCPmCjfsEl92HXHrl+BiZEcNOtPnWDOFaqaX1fnamlpvg42sVkwAFx1Etuicr
pX+pqK184ohzYvjjAJcWnDUwucxeMTiBt7Vf49puHH5x/Xgvz70XjK0hje2VmhEfqjwFwdin+NB9
y5nf2+cwx9wpUnjjSGR/zD84uEaVYz35U213EaMPrxdR/HIJeiRgUfIkeHFebuvRi8+LS3RD1zSw
6KxbDNopjNGPOrLtdGhRUMrpgnOAOCqUhNFophUUQVQLZvGvKzMU+MuCc4UDamgJguYb1zJwNXDW
DVlTSzmW47fEAk0SQxoLkqP9plX4Q1IfugOkoMFuGxGV5Jny5tOQEzMji5/GU//1A0KxX5WeVLjL
y8uGxal2NFwg8PPvRoWIPZtArLbJCpiKtrXyZ2/kIJU5HdGXy4WmmbODwyZHs7N2JvJhj0/lXdHS
PSk0YNkTP0cyf+s3XyL/nmGQ3gTsQ+bpQzld0L3yYxZS8fFwfMTFwaAE+YyiJi/F0hCLLI/Tshb7
Ww2p4qdDl7/Mwlb5Td6XmW3pyQmttvXbdzdvFy5V2QeBGmiwbcfPTiXQsOJa84f+9T2XT2vi0RIO
qdLE9vssFHKVdfMqKAPXNwRwYyjguBmfsfWY5GeOgz4IPE2WmXKcaRg60YJH1ScDM/fmcpukUli6
g5CW5wiJWDTZnQAtFr853Nt0O9Z0NII/YLqRlx9jE2Hb9OZNUwxjKnVr9u28Cb7+/wu3uXEl6wcC
9+Ca6gA0ChEA+ELam9AEwR9nX60/AOKYQkBFx5PbZxxnrS9tXfKUXns8j3wqnm6HKNLKzXtT0Lpg
8TJDSSoq5icOXd0j/xYUbVFS8r/s7VvbpW/06U27rwdrklD2QxG5dkKsLXJFAtWoDi6WgsL82b56
eMlxxv/8mO+XLua2+rUPn00xVAF7VjredLJTQeYrUb1A2x9gxs2CaTYf/pydb3Sr/wneuHLEoltQ
zfFFZ2oxBQc4kVt2ATf6Scnq5/IwmCiaEvm07sq1mklB7sJ0iSrY6gRFw+d01jZ3Iyg5eL7+lEkM
JhI5ER4lGeWbjgMMqbqbqK8yQwpplJPqxWRovlMfqWPcQkMktUUaxfVagm2nZ69ZiUXtO5WHIN1p
sJLPDFC3F+HJBexnYcC7EoMwNadzpHQa65vxHWGMVKWgD5E0YtfjJvn8A37ZKZILabn7cpHfbTyR
sCw74+OG66sBY98TTz/v6LiN4ac4RgnO390zJYxNjTWyFi2VIzUSq4PR0qd1Ytt9B1Kp2k+9hEHC
iJRXsCoIQ0qcJBBqnNfaD9ToG6TmiwZXj38/i7K2IJTmUvrpjdxL2JavxlnEwKMkW4tyuf0N8Hv9
MUfrlItDRJNbectrfC0AWlcdsxD4CWAOUw0HuEe7ldvxGgUdXSLTUW8rFZCTa3vdCSajAKBGTHwF
5BCtmYQ5tWj8jB6hCLhvHAWRM6pG0nDWf2wMXH215P1NsdV7V6X1CHYpNqZxGj8cnVENvCdOIiLd
+BgjsFZLsa6NHYq5qeJW+z3uGouzsNNw4GMZbhQqlMHEDgRD5Rr9OkSmAQKUdSmy/Y2nmjC4LV5a
p0aPp+5IsTd7akJ9udAzkWjC9VBmFwnQb91+tovzXcu4YnI+AAowyaxvHS6ncuCWqpPaZMM0vkMJ
JkcecvpkbKCeUo7e9O1uFyJ6oVzS3X3ULyFJOC3n2DEeRnzOfFpK8BEo2zJEMnSNpEz1MQQjIiKK
MHwvwwS3c9G1zpc0gLOZab8JWSlMUM5jK5426NvhAqQimrsxvCp17jx70+AWFAAdfgsVcIc/37B6
9ZlBWd7oF30SANT6m8vnDZgNNDS4NaJ+Geqc49/1PU0vwVbdXExwlxCxa/Z3sIAqUTc0Hy0958g8
iFqFaeE20uYFw1PWwc7Qwo0Vn4OGwQcsPhsUA0XZxuQR8cAURn4Zctjy0U2Gg6RfoIs4i8cGnfCg
nE1fJhw/vfSe08qHHLTJW+KOR/DYAqJUdVDFr0wnu4/VXwZukUHixaedJNIO1tLhsNaKMnRLJxwk
0VdgVfTappX3pUo+B17Jj/tH7Dk0GKtvczwmsnrQzmEMuEje9aXCkKepRPzk4jmnUPvqsTETfwzO
eD71+ITkEfmuqY0SnYNCZgfGLTa5WWzmOBQtm6FMse2p86j0UbSy8Qy1TKc0HPwoCaBntMmAcYUr
Lxx0w5wgNVXEkOvoybpuuApIgeax+bHeplj4t4KD/OQ/js0P4m3/p+EsWCOp9H7B/99+s861nnuB
O+JG4nsxgEPy+OPoZHTOckbUvYdUfbNtWcQ1eSjytOqqYfhV2deOKzpOARCaG1flSFeH7g+YdVHj
aEEBHOExOfiANOeDxgwIg3jl/eVo69peYdNhwJZuUAE1QIq8EbTXJow9wt26f9xLi+7bdN47Eo2B
34uLTQbwpV+npLliq/0dwNoHC1oGprX96s4XddfteToKdv7o5iLxeEExQDku46pWW23CcO3qkQ4j
H7Uc3z44UxNAjE044jWWSjqz0+BYl1eVkiwd2fsopcmvp1RPG4nobCsKOsKjim0LTS9N91CEPDxn
DTWOj/0M//y0Asjfxglw8zVmJ3ZfoAqYJysjja7dR3IQbjr39HjsTx4XydRFgaEoQls9qrR8ovLO
7kJ0kHmZTjbJv2J4CzFUhUjaRfIBfLsliM1fKTxpMxw+MaiTFbENNhI4jh6aNcimoEYHEN64t8ny
5bpQsMrw7+V/2al+EDOe33Rs5k12ywEcGrF9a+k1amFK8oFMt/QBGpyb7LrbETBqQt2zk1m/Q/+z
BEfgPv4eSQaF5uLpheaKazF24YCpB/ebSKhsejXMX6ZFEOFtKOpkEGS5LigxIA/4W+DaP48if7/2
csYqr6wez3SWOnVV11bvPdNYl36gZ9erI+w1iC5mp6NM9h4xWECOe2zdz5MyJH1cJdTGy0T1PrWg
Z+SnJp+bLnRL2n0Bi3C681KlqmS3a0i4VcyR8853XylEPfakUSZv4KvRhff0Ctk2ezpYOWw8clTx
bALmwH8djohuFX5kHwHpGjfSNOUQnWIdm3c3WlTTIar6ssIxIVQ1raYAMHwFYusDFAtfB/faH6ju
xWaOJnWBZM/lHoOSDWQHBBFivixlqqqHeE8hp8L42Cjwu0UYtF+0pfwSeY53vZk4HXOSVlVk1Cbc
OpL6KDhpN/0h7qPH1l3sosvvV0ouDvcWvOnrrDCrPy4nnJ/MaBkDenlLZFj+A34gEd21rBKRtPrx
/9+LJR5K+zXrnOZb7jRjePwKOPRiuULSM6ErnhwWzyGOkPynQQqLc5cf9Qd2vJCl2rEsywG/TzYc
BDryDIVux7HiCp1XWjWkTrafi9FPQNmicsbRISouRfzSmIk6/MXjsZm9LZdTHHMqIRSgimglo3WM
FkrEQvCbeRpULyFOeOBoSBIynTNYZACD2abptVHF+6IiYjSj4vCNOFIIb25QZKY0CpMHRy66XKtM
jma+QWbZi3OLoEgNBBZXAViBtOJQGx7zBgUnWJvM2134VSS6fj3Fu/ga7DD/7x4p1omNuZFv38yU
cp4FN9v676sg4lBFsK9wWx/PzJS+DLFON02uDWOOLFYb46sbo1wm7X9iGEM43Vq59z7qjrxMUMrt
xKgoClcAzyOVCiXLzwwmYrrt6XuvyvcKnRYoEwenPLytr6HTO40okWpQXK2f9Mr3bAqe92f+w2kZ
Sz0CBrglEzlk5kvFXlZ+KcrL7WSiZlSIYgXO0+BowkCtVU1qV/VPIkwyEgmluhF+j01fKWY3gUME
x7Q7FLCAYnAAuIzxGmUzGQtXZESJRrJS8gB+d8IXEDeWFi7Y+6+Flnu8YiW4aMOgH3D9PAEAUe0N
nlGjvF7GwNq04MWwfsvGetVfj3EC6oVGS4DanupIdIc+BVsvObF0eArAllPNDCZmirjTQqGOIvzR
cPl8nT5kmFBMZtdKDZHATksBhZA210qKMc+iHQ3n8WJ85sobtrab5D8dij8piv46iXXkESor9czo
+2PeyUp9FdtJGZRgCJGYMrwpQ0EXZASjNd3QmJRW4+vGoBdqi2WPuCsImV43F1ljsuM7vKZgxmU1
KQ7n8W6R0u5JzbCdtDXcmkr9wlhPbTlVsIuPr1csuLk7Aqb034Ye0+OiJ/6UGevu80NRQN2r4PgA
5lQM1shSDnzMKICIX5QP9tM/DD9QoRj+5feEclSbXR9abIXjV4zp3aPfq7hD/pMhHYJsNi77FUgl
lrl6koP90sDohfFF80aGiH/ea3nYfq2LHn1jNcz15EAlhhnx6QiyKEw5A6Bs92hC19dlSaIauaEA
61Iqoeeyb3ygYjcdl0iZXnnFPJ0LuuGCGEQnD1kJAfmOlkHR1u/WnrjWZDEt5r0P836nNvgTU8yp
7KkDBt2Stil78hMaxcgX3YQ5jGrIvU9WVwwlzVDYW0cDFr/HOC8JUgZsOgGkjcmPshTiSiSzlYin
wlIAoSpW7rBQhzFvqCxpFS/SCtJEySXwGUvhEfrR8W71QTpvMdOlfiiD1pTtHWAAHabLoPAlwCQa
M0ypWLcV/Do3ORzk1I3hxMVPkIDIqX81+718LL5TW0ipTB8ThJwGoZp0xG4AN1qqG4QuQjfRHG+k
7iQvpMBhbiuf0/I1Ulch2HAyQAIRAudoXPnmKVFXZ67XGT3bwSOwkAimH3/67FQyogsPORJ13Ab6
gTdPPtZZ25loLSAhJONqUNLxj/PZXYreQ/AwKR4EFu67a94iurzOSCNkRFlpyY7Ia6X2bt9DE2+y
+p7VYQdb6JXUzmUsSFq/dcCw0fAly0FwONiNB9PoXWOiQ4JrMxWgBtNkeoB3y8CybGNktBSl5ASg
M0G5DVDfnb3sp6P9khjNp9ezccW5uLYWo0SGwn7HVD0wsFrRlBzqXErV5J1QFvB4EQLBn4Yl+EpQ
5Fzl6YXG69Tv0Zrk5bxPxCURWiZzqDdnChVsnwqo0vqxf7di3RDL2pPH4gnTdxG6mvvNy+DmnCXP
UlOqJgbfd9EpqELXGJlrOf2TbUUMlzMHDmL9b7bC6215etE3QQpDrekivTO9FX1ilDp/yTHnto3M
+aoYswciAHlopI1cVlav7iRr1GxXewfB9M/wVQcqcb8xEfmASjTmcKNG3Rr51eBUnRH0TStkF2Ib
5114TpxC5guAIzwgWWeDs1DRx4Ie+ducrAeGZq4zP6el0aIEf8TKIsBoxa/heDCSGx0+zDfVR7/w
/mnmEjLqgg403fl+JY+RGJI2hU3pyGpNf/zuSejfY3cx2qaVOrx3Z4lm/XHZkTsiwm4WzgqebSnt
rwiFokf1iLu/UGtEc2F/SgwS1NIV1ckrelcf7gCUNm0lnXJFYzse0axHEYICHj86jdtXuMzAV/SQ
elnjY0nKgyy8hspOWAKl/w1trClaaC52PswqUGsOk4CFjjjqwlfkRURNqunWpdcEq/qQBhqdOk0X
+pcvGQ4Ntib7X3y9+3a7ED6Z6yihRbpIq4sMZoa8eh7bN/MAINlk16K0pnXc7fbBT54Vg8r+7u6u
iLNII6c0cwQL8YPoS6yUOZqqnLwVuASC+EmmMVTM6tbI0iF+oKaIFIbIWcDTHzEzK9MqbarZl7w/
AChhSolLXLkAIPOOlH72wIRWTllG+djj0sKM7FYXJ2qH8/VJye68UnFyNGEDt/NR77w2vVDbkeVG
clax/h6Ym9lXywDmKeB1mXrgH0IgzDAPeWo7if+Pt+ITxDpiiot1z7bC11ffKqp0qCphOUw/1wqP
CJFkbnxzXczz4vNHYPTXTPXX0p17xR63dQaXZycG6hRvdBDKCTn7h8kowzZI533aPuzlK5egsJU1
G/1aVdf99rT7qTy4CtCTAfuzp4+c1urspejfLSV6FEVdRUEWhWfYIU+K9msrw/Cfz+WqYTevowIp
i2oSU5mxM6ebBYiMnAQM1iVLWywmqlNZ3mIdXl8UC9TkLqjNkIWd6+JbrjB1FdI1R8k/EL+rQ6bG
0oMFpKH5pbeVw3H6wYHgud8r7fpXIzbPlg18q7GSkqR0XgnYnzf3RCPED9QD9uYUlergjzAUI5nC
dXcBnIw3VAsd6oQ73Jy3MzAwOU1VtegD4td9uF2piu6rnoJaEvP/tEu2pZ0KFb0g8+mn5o6AGZ2P
08dv5UOF8clcAiXTKrStZLn8tY0E25c8upMhD4+50rOlh1st9tmfa9eieeaPOFv5mSuwNlmW3Jw7
09OuTQ2xlgTZvAsr/pUEyTgPKvpeBuTRMCjRi+kBihoVABFnAm/yvzE3uwvEgcZM1m9K5MoqSqjd
GMKjKhqghOKEwU4fU+fWMwO09/c4hp67e8i9iHoqugG+T9iBL4rXCsd/kqoR+dYrp5f0/658UTpZ
d+682stuMuH+Izgr9nsw/XlfMLStOopGEwlLfJpCFCFcPlCr7xCdlUiltyEP8G2Z73uiqo2uzFxy
dx9JeyYWafrS3ik8Zwt146o3CJznMYPMuBTxV+TA1Y7Qzitdo5D/VaOJ/4sNBGqJb5pYINOBNUEi
YO2QPUoxRvSzJcfMV0sHLpH15d/VhSpTHEW9ovKAYKAi4An927yMeqpdKbpVmR35Ygm9byXev419
CCLFjEGFAROE+vPyAk4iKSd7keAwg8xuxmAggdSTBMGPS6Lp4czba2xRgTs0FPPabc6D86JfYes1
TniAH17+myH75ZnEz3/KX3QiJGWPjUm2TgcI9GsvqLI/NlZ1gyOaIuQpr6++YjnJagAk5hR6Q1DC
VKteIo63lu/AmaCiEI7pn3zDa5kHQ5qqz3SN57MhKnUZFlcR5QB/eHcLmSmLmDZ9NUr5Mfwobyoe
Lm3oLGNOusCaLdEA2SDqdv9bSdEwKSgBmYwIw9cJpJqJS1/yDNOhYZ9ztaxeNCKPcLLzzKgKxeUP
1zwA48jppwZyF04WR5lEUqpRNUl6i/9d8EwN5FD1pHcMdFH7CdPzx1n5JIGr0BJ2Pf8l+weexipP
yPAWWB0aCJEAlUUJghzcgEKOPeZVQW4VT8zGAyiLK36s+a68uu+nS/EtVkd9op6H943hGcF05ZbT
NifvVG95X3fP43128UlHZh9wV3WV8jXxw9FjcYzBE6lk9e2E2y6KN1BOGSY7HEbUuEvPl5ZHi4ns
aGZ17OLzYfUFPZdMwrGduFRZB4AsxQavBzDHBe2u/jbXUWurwN+pvBpqUCR9pNGLYvUrUL5bFTuS
bl/aSldHeffNwyvtdve0oaPgTuyZz07whhIoWpxnivMmmpDUUUu+S9R4diVnlT08BdMi7t+yM5Ox
ilxOZSJYilImKSZ4Sxol5j/ScqFMvukiBcBChWeIXuza5urFfCF0lXw67RfyRkHyazlduaShzXlZ
YsELpgdezMugO5wThYMvnO35n/1VVDYHNdDGQ4dOLBLCDhcXvz5/7UraNsjEUarIIEOdABDnwFcP
eAMcrqV4kJWRN+LF9JE+GxB4FAMNLdhprk34KvVifoBOdMOh/H82e4t7tQmHiREV6Whfs+OGV6YK
kfxWAu4miiNIx3SouIzIyFHfeMIkXwkzfls3ZJ1Oe/nNS7pHmmgSLPfos5hXBx9bIk4wshQeceVL
Ty4gBWOTcYfuXBhKqMidX1Orq6LaY9QRxQKJudef4G667Py5nQjWVojzoTNvtpc7BLD219L4PITk
Gi0XUDEfae6B66iAIMsQNj/KqY9sBSQEmyeGGJscqZobt4r2oY1TDiUccr50r+UzZ5aoXudXHZic
mk8WZA5IZqJvR75e1irftOW6Gqkh8ixPZ8tmM5Cz/ZsWxrACbfxjmUO3egHMg0aoDvoTG9hRx1bt
dX8E7No509feAz0xWRSjM5fARldT/5Il8DPZ2V4eoTovgw8YAOwZQsTQfCPo7nFoDsgSxDlafHuC
lRmPvLOedblHGVRjjf9hvCTFar9gUhhnNu3YyGd4yuzZCkMI33uQiqv2AdcSYSYO7RqN4p7YQb/L
uKYgRCVkkd8zUfhkRNVdiIB9yBGBqmjuzdSSJU79ogmCgh907eNFXrseThwo6ExEb3Pm/2KtRwIb
MjZgM32hHffLQsmPtkLJXbJhbjEuKRMTcT11koDkxCiIs0DJc/HFUQTfW0OazjU6joCQNZtcbFG/
r1nR/1kN945N24KWnrpAxDbc9cltqY0bldeLXbzDjRhfEwEz2F3M+A2mwFl1Hr9MjbQ+mzxS2umk
ZR4Wb+BD8BgZ/NHjv/LQulcGVFMce5GO8FAHnui5l96lDfXDnE5L/A7BYkIN/8Uh4cOcGxuaBHgp
y1GqTa4CAABdtQBd8PX08Tw6eX+Z7XRof9xYw6nQ8ZOfr2Ra7n3miHlpd+UGGIMlHTT3Y7ZyFsR3
CIQBedBNLbAXbRwx6/cPCB930GszRaSjoZ5aQfelAmRv/SNtVsi0pYCxQpzILDxT6cSZEG+KG4iV
ityC3ZOoRkCadCBN457ihUGcfW5mCP6cvs6Po4y/V2oFVPSzi+U9s+hhE52jCIuPk4kDLm1DANl6
WrsTM3dta+FP4jHZMivCyhq9rH8/orH6lPFFibR+XCJ0HDqDBxYi/lkIi5Sh1itchS96lufcY8WO
YJoxWoGEUGksJnVAqQbhcDH5iBlnI2UOrkh5aubaJNcaMkABcPjdtY2GhiUBq1rOl0PtxKBuHO+Y
jotSd8BTpSYAqG4cLp58JmJcFPjuOH9oXIav0npRmcEdo53u2fh036b/sOTwINEx+K/Hg4Soo4n5
Zk/Zh1N77gfhk2ZZJGrZDmnyd6QDN6C89NZS2AL/34h0TDPVpLQsj75EQ5fWMSCGmYOnNBLzOAfV
5ecbUGl6TjWgeUJ/fLTmCYE4/zaqLnXNqGotcO1PldIMil/gOalJSqoo935kLoZjX6UIzbu1WrE1
sNgOsxgLguFJf4Wk22t6tvijonWnJ9R1ilDiwbVJiRnnHqMWm7NlAgs69RsMFvGeCwsQbHDN2N/u
sUvJYm4/ruf0Ys2Ki4fapC13DQ8vbcxFSaeZS+NkBU9ATlTVNAlxS2Gy3eqvTPirF8VBgtAcJj/X
0zT/zNGxvenacOWt1D8/Nr4mKlkADzZOG6+wtJsJwOl1FA1BwaSDfuot5HwpzvCnsXpFfAlpRP7c
qoCBCijzkjnzEsxJw/bSKj/fdxrIV3OJ3/gah8Gb9g+ZDNdHy1QaJRp0Id4pKHwAVAF+7VmwXkhM
20PA9mka8ix7QONhHrpGGTVTtAvfkttlu+b/tqb4dYGGNxb2cCJajFI6WLGbXov5z22k0sn2AYho
EPkh9hU1DtzKYc6ODu6REs/JJK53QtaWWv8gvcgJ7EQFVx8hofq2munU2vu/26+qd4RFv5yyXTtZ
KtHxnGHf1H7Nb6qPLfOajGxB9d+G+/8glZiz8wr3ff5kB7N3JjlcQh/9smY7bzEktc+6KpesMnm6
luMe8pENYjx3TccQeeu94aiN0H0Qk418mZlV/ZHTDeirmkHPIVCN84SNFsbUsubzNz4+vPDZl4Dv
VpShRbRYmOUkr2Tdtm/Dj9tCn0S2+ADFzmSPRUxdH8adw9bsobuHGo34QLlqwPtzmYQvNKoTcz4O
k5C7UMp+dqn9EHrUw9XuNQF3CJzegqrK9LSj9f4spx8LNsYc3v6iM1rPFLRmLF5HRWeqWljRGt/G
vxmj/A4SDlRidVjMiQbRsGr19ZRCMD9Olu3cWsF5vtaR/+lz8vEqRjaN7SfV9kEaREQKX49p6+ZF
LJhkkPTucunLpgeY0PdFBRPmEe32nF7rprrgibwucpEjfLTubkQmSzuQcb/IE4TDHgsWenhlr4NB
EY8BRKk7bq/CMWAJPWAAbzOmuKr+bVOsP/SObH6uS1RtTeEdzTXbA651ae7RZ6NXllUDQd9RwCJL
i7zS/L1GuRUPkMToa+kSWRx8cAXppeyRZ2iKv0FJhGTu9JqHubkAiG2NjHdIWPb781Y55ViFhK8a
LfAbhNmDkPpQKk5767P8cVZuw3d4uRlDr+dIqq3zyLViFqexsxTiyVl3umrKzNOrLLf6uyVJcQD1
QoNZC3XJoxQLc/fJG+BzRWee2STFfh5k0D2D0ZgwHsizn6BvDSUmHtS9RqFWm4ZT+/voWQ8I6UHn
H4okE+hx6Eb+xdm7LCaWlz842fbD6Sp7uwcyNNhw6Nqv09puec30Nqxzr93vB0nzbFQ7PixpgcqE
fLPazNyTofUEZqyPVR2gFRNmaJjmQ+sxd6h30UoErVvL72dUddRT7SLf0rfxFk0y861smvtRXt+0
R/NL4EDV8Ze6w9jZ4k3wIV/y3r8zObRFIov5yIpVOErr4lWYAe23OpsTNyeBVrH3wZ2AvjpR+J7W
ROfiHdOPg4zcqoZTVN7KD+wB4VlqR7vygBQ8L168RGSCpmz2wEH8+ZSFyJD6TFE3ryIcNRLGnPSv
7ghMl3cKzji8xl3rLoqHfy3l0Q2+A0zm0P2pUmBq8+L3PfaIPaCX690MCF+vZw0Y1lNMqt6kMz/f
60m+wbdHJKGX/tWSDNKawBCScizh+KaER7ySN3GNYedJg4TuxaTsxG4EHZrpuNWZ4ThU3jX7TSKg
K6kuCPURAIB6WHn1VXpVDdEWtMLOzxmYd/AobQYdV/R6p4mUKF9VwzN+mSimcrsgr6g+BMuQHc6x
AFGwz9GpMMQbhWw6blUeZND4anfJ2ThsOjwP0AsnSqDbNpa9ZAQletvAcHK+3t+TXOjv6Whcwujz
TVWs3vPw6CCnZf5e/3PEhS5gc1z2IJ+hddlx/pPjo1/LHPDJP2mznmEiWmWB/G0yAGKDwzSdyLpU
RaYLecVoJ5oMlmumQGzXEAgwc9bkhGz9B6lh4FZHE4tfR9gw87HwF79Hpnc7gYyHaes8VoVZtVUi
1Jpq28EfnKogjqODty7no0oPuWfnpORWen/0Et4IlcTd+QGAH+fkYhAeTgQqqCrKPCMlf/leHIYz
ASEwY2FuuKyrVzfHP4PBB5aOaQg59I6++UruHYSO+rnNUONWH07aQe76NRBwDxUDjfU98toGDQ35
6E6ju0Q4drcS0FAbFnpZsRLG/L1kw1FMqg7yU0rmQwLkimh8AOLrzVIFKq1xIyqeaLkUrQA0r4CH
XOywYQEfVsDlkDuyyTR96/sA45qR6ctbT9hNL4h8zCbOjE6Av9bTLEUdjmVfPaZlH5DHtPdlDeMs
RSWm454vnPNPSNVsl/++GT56+jjQjpm/GBokQVIosSBxkRVAAEn/f87o3z79In/l08GLOz5Q2AF0
u/92hnK4MtsG3kbNc5EjxGVhd4TeWqgaeY+cL1vBlRqVXiVOBR/00LunruUs5yp5T8c9KLcBbpc2
/ISWZRRDSmzbZ8mwFcBbNgE62tvBtmld7ovf44JNTNxroO8esIhfybZYX56XQ6zeXXSmiOr7VAUr
F2lw+d0vCz+nZYbduFzjKIk0na3qFaSzVDF+BnMKr4W5ADlPtm72lPAMDGNB1m6Ot7Irmour48u1
TUlmpXrpA5xrDps69Ij3Qy96Wn4ZjkWr4Wp+UX/XljD3N/TXgq8urFn/zPSycMFNkd58dOw+tYQd
Er1HMg3vErHlvccDdbYTzweLuJXYQDiN3Ld7t5E47QUNfvKen246nxs8qEnKyVn77UvoK88BuAeL
86yu/IKyqMt2y1PCfES50uqp/ADLR/NQ4PczAvVOKZyTJV2zfiJFKWdNXN57ykho+vQJazFdXEM5
koRSgdSjuz6m63LIkF2fBdQgRSB+oE8zmY65Jt3JDjAWdvjbqYsLno3RwSCrCl80pKFBgh4xKRGg
v/Xn7uzegw1fpWhNTr57T1dUH+NXp9RfjNH8mSalAbEcs6WjzmR8XgW9kytde2id3JVVqjqpIitU
mTV1kfT9JSjEo6MM0amgJmUbt3H6OiGb0k/AxB5tTO61P2IBYjSr9ihsRM1ZGCzE/wLZe1RbA06M
y4MEPe9SmJdmD9MSaKEOI1oBfGfggDDakokhr5zZzvAxZT2GYUJoCto0BdP7rDk+3NZsfSp5btXm
GA2LcFS94uv3iQGuBUSKVX0uimik87iTXS/9hH/IzqaXs9LVyhH71fGswuwluFMlU7L1CSvZcm29
GfezPgOEWRaZan2oHJx1AdVWL+g+B7+j73sDmRUlPJQPIBMriWG5WoIhZTCvblC4NyjTYeTH3cFm
lT/gPqQRQhydpSjZuM8naYKJEK4yCuEpmC7wXavaDW7JcVwuaL1R3Kqz5kgmKjDBtrtleAxQRpiZ
IigaVJ4+0rHMvsKSxZ8COw9OQ55xHogSAdwCCTk/En1qHU+Xj9BsUEAmzHPtzpwPy521GqRvhmDl
QcmrHpY7QeM50HP56K8mUapPyU9UELels6b5+eVl2p64MXq15KawoDx2qt3k1BQ0DpIRucBkGjCL
r2yq4+oFZ4AfMi+XR0ZBC99BIouFuuhnL4cfOulWEI6B6jofvzeucHTSweW3iVF/SiEF/srQESm2
xM3RF0PTtzGeb+hVALuXUbxCwPXNw520Xhq88IVH04y1VYNCspJSmSOGxY2njOpMIgQJ3wTFuUVK
e7tUg4ULPVxicCH1dX4+85MP6aLnE2kv7xgU4D0SZ14vzh6YnD69wyIO5T4rIAbrTCX61mWi3dtA
suXKSF51eFCFJMCKHD+4RVI7wP8WCDAeNUYlIlqI6Qm0SVH4FlJFpuoeP6t/iQgjRHY66BlXdKJq
/OtLOfessLSLu/E1zauj3J8aOurB4QLaA1tEQn6mu2cuGfVPtXoT0+g0/mS9PjXXIK12aAwucsgi
QjAT5u9rb3+9lTThHDG4mxtp6pRyE0KeEa44aVsvfy7j4ZBzIWrxOwKP762HsgVerLHNb7jEZgcO
1RE1fg0MdQ37G6N9zuHK0QO9KkOhWK3wFHHE22Xz4MGANgLDRrCtwNt/4lXkxCGiuBPxf9/D3jLQ
Lrs/30tZTB7jPi9YKR52VbcXqe7BP8tbYSif9WS1nYzh3mBtXJF8wpZCxzkYgBUWlfhmZ92AvEyb
yuqOmWt2ysi6vr4pPdEpAEagtgBli4JpSvNBQLZgkUUsRS6jxQoaXAF0wTQmxHHbbuW6+U8GfJXJ
th1PcJAi40hdjyT/xn+lx4ZVBwJ+k5iLVa+B4azuTGQy3qXN+/lWXKGCdOcKIPk76481Ah1Fo5jy
A6xuyK2LQbWTW3zSX9qZ9FEt4/xJC2LdpxCcY5/Ffzwk0lalDNtG3TRrW9aB3eryH8sTQQ2JBIVb
SXSXIy5VSVAUpKhbYaiNHAH0/J5UkKbS8yqgHP4EjvBPG3JJk7p9WVQfqZ974M4vMYIDc/RlKV+W
3t0ZH5AdQ3g7rEkLPfOirLpIqgfGveolD8cxNZGFyj+ZQIApbgyqETCTdbCKj8UOZLxMUFLwsOaU
W1Vp0nIHNOJQnf1w+PAg9ZZrC9+q0ZkokW8edGchHvukRqwLgF+YEV0pwCftoGmcQTmacRZ0MuGg
9VxsNZuIqa9OODxggnygTKsfr3v2+HbdmL/rR9/C6BzS1tD8vquJtl8Bkmast7TBKqGWufRGxoFZ
F8w8n1/dbXxx9I2JhP/l0G9oTIoioKrFmwDMAsVc+tbvQAix6a4zbJTLRwsvVRNAUezYvnxcrdgR
GvqPrcoaGO79hFQdYAdHpd0b1SMXkkwTWNDIwfIe8pDjhJ0ZBDFgvf++VFBzl2XZ4XjHN2spEwQR
KssOst0tL4x5/lR4qhb4CUhLQ3SyMSS7iSUMkjCA5RtKmI/RrScQ5QIRCRbKvosbAl1wKHyx+El1
aRQlb4OO1eXY0UhgrFkNzXDovb9BDI8RY8rs5EzUQNgHI1QIAbjWXT1adzzJo6+gsuVD+AuiXe5t
Y4tyEHuEBTcMrUeNodNEPiJ0osmbm5+0DjrtOtYvt9x9JMRYZyIYFQD+2ZdUQxwntmu0w7+A+L4B
gE6keyIX6KqX+zNeXkBx38j2m0NR/57tntNPEMrhpWfXz4Pqx7fG9WRz5urRDa9JXHlpZCDJfX2Y
pGyR60AVm4SO+XAvBpaVejABHuFhZ4Q2KfJBgJLu54sidcrXdXarZgMojzE2hdr+YS0uysEtKVcS
pJsfeMdfTa4w4xQmPwFSRKcVafjcO5xQFon0RNzLjCHnZ5d4nH5muDVS3/XFHBE8HKYi2gm6sWjg
SIOD1/KQLKe42RcpwcugUmC5bwwXLwyPRRdRqr+LrOvJagjYSkZct8cb5gBv0t50VVwpibRL8c7o
llRrS3mjOo/jon+h6tqxPTpDhbmHVTymKs7y7A7drWDMajhDthSgBWkJSta7PyeJ6X4L5gcDCm3z
qwLMaGqwlY76ZLrA/s5t9fzIyeIXllhjZd90oSntpkqIoMZY6uIMDZLLRrrAjYljKO/GuvQFprX9
0et1rCFFJ9LLTBKjwtLYECCN1S/8Cp54BLNISjIqqA0rTEeYw7NWOXVNmcJbST8RYeZWDq21lvcj
xm5MFA69hZ0ksPNqX+pXmtVnnqwrZllJ2KROSmXeFQ9wpvDDGhPmZcpnHH0HBtmVveP3y/jGVwJf
exRMbrGOKAhw/lOxtUhGTHiBNeR7q5P8ucC06NM8ZqYciIN4TxLQCNnaNbmurOyT+ewvCR59ecS5
LLSDhtNh5xuNrtNdVewribwbrmLeTGY8bA1TTpU6iiCyi/0/BUxJj3woQVxXm+RPEI1HNWXC8SZD
xblPDQFHj+AsoCP+iZx57IBA4i20ltvMb2DudppTraFoaHsAu4c2z5SaepkeQ3Un3IuUf22CT+HJ
Bd/jjLaDiv5OaV6PdgX7lqWS2BbynNOb2elQ8V2d7jHGDJwYrGOTgak/biEOVIlyJUr5sXk4oka4
4olqD7sgrozjOx090iVx0kgzvHELoiaMsCe+DWnTljDPjkGPdxZv+KgdeNxEvOBdD/Twss0O8LWT
ddLA/7jBGWJSHYEfuVqiYHNDjOkqdp85h9z9g8dyvEuaLKILbh0T8gRGZQB+vChk4LBmNLIQ80ej
XXg1bJngEWWVMJGDtkn7VEhavHltnsxVxskqS+y2fc22yhx9c+4v4vSqZDCMT08sQZhvYnzu31zD
Vnm2Qu/nuLytxRTkNHjWsNqJum6weOMD0zAKAVjlVC5Q355C3qCPERcbOZDil4rYHRjc4Q7+vTjt
lgJ07DljFr/5VZlg6uxlUqL2l0x5PcKKolLUwTj9U5Zo+Y1E0SVcsuSYGGzsepARQuYKf/zgETev
R/niR8azg11YnDng4kt6BbbWBQsAGc2qXHWYo++DkKviFhJozETZLt9jC2kdcvP3tHTVDxmOgy/t
C+tz6unDAAHmoPbnGtETgH8tw8KNuxMmOGeJ6QxDRE0UHJKr9WSoyvhyapQuksdTbuRBHv5IMpjd
LuT2Hab7ihk6vWC2thEqEmh0ZbFRqth6Wvg7qwxd+BvG0eSTZxukNkndsAYYfmebgPcblshJTV2f
3qlQyMY2HqKrkq0+yXVme4MURnbRuY7MWq5baprLNIsT7gZCm3gS1W2mlMjjcWdklgjKGIYzmzec
N7/qlqhCdjpEqbRkbOiMCd5QbLgTriOk2yC7Ir1tGViqEA45WhcBMiMn+mgZ1n88ezb0IFOoKQEj
7dUv2Wr8/Cf4T2l7aTJNDgDLxbxqwmQDR8ePB/dehqk7vzTAPsFJxp2eMW275FeGDTiZGjTTOJAc
FTLM9BweCvn+V1kQyf0sF9VMTgmxsfkwzccYNJcsIRYm/FuAu0JDBgKucsEW7+DiXEtK64aATZeZ
ncCd6Pbb81XZV2NFOECeISpfADApqQgohP0Bn1hrxMR2+IZzjNjLznu7HugIscOQSqkqyhzn6WbY
jY4r8YU3EKLmPqsnBn5nvl8cunoQDZ/94Mgtpmuaho5f+gsN/vU6OhA0Yj5foVFsd1o+Ptp4q3qU
K18jF+UPe65LNAM91ipdeUrKXTF70VwFqfd7J5xGZQ2fqzXxRqbMpWPzXeQFdPTO6SuQNcKVQzX1
BGrVt0ttHDonTwZ+0v0NsbcxZJ9bU7R02xnv1Q4Ecf5dptgPWO8O5dKDjxHkE7cHhbS5z9w62hu7
shQcCJ+yF42QKMPA2vT5uiN/1Y5mo2HSbbUUodmYXaCukf0G9blhJie4ejbUSB4dU5VseQesOZ2Q
mRd9R2+P9wATbLl4bYdLGIvWyz2hDDjznahp5WgfunQ9Z1mP2H4oItL752TrLaNWclgWNkyr/ds9
bvKG+9x8ec0SPOw3oau6fd/uUCn0txhxsnp97OE08crAYQRk8Jf11CltrGY6a5ar3kBe7wxTwStu
1Py5C7thNaayuBBJ5I0ggZZ+vDkhcal+VSZwLCz/jsYaRPPn5UoWUEw9jWTYzU1WGv8V+m1pfYq3
EVcoS9ZFmwzicUx4DqtgtvBbQmkbNCrHK53vY1eZt7Bu7BO8+yIQnE3RFBbXM2sAgZEscxf4deix
y702D4NrfRD1l2zIKFhi4Se2TIb20QhGQgH+empAvckxj4/kq0S8eO4dsx8XZeoZLZgLSUW7Z0Kr
Fgd80KaAonPa/mRcowiL1k4Ly196ucboXNwMDLk89VULbjUqeLM1t11Do9C9QYtV4f9Dq8di2xnk
l9deqvH8xlhtQplzUvV44tYDmlJn6lDYdoL0dYjOGHUaC0bfHdXdX5YZh6dUHGwGl8PKRXuMhj/F
Saa99FYfg3oaD5DfsmFk6U/CxIOLzKkMssDOt1ef8GhnEo718+3jkqJtFZtLsZEQMoqEhvUX0xPI
xgKRqyVBxOSs9Be9yVcHbViv87vCOUN2EOGIL7xlJUhHqGl/YyI9qTSPXeqxjdor7sbup3Xt6ASo
NcaB6S1lqVCCZ7QGY3StCNcMpjCE6INVTlWhUhpV10Y7x3lp74uJYeLKYaBDOzmTwfRJ3XeSSRxi
OK7ymDlEnF15dlgd5XKeq886ypOvptzkMY+0SRGvISoI+UD/F8g5hv9cjES8oBScwNR3pUOw/qsE
BxNwmy0s///qA0SPxoSLxHmvovR1vVkkUC+yzOlQqftDl+/ZoxQ0qqrvrv1NFFop/34EgTal5BRv
53t/XHDrOzFWZPRWIZBQDQgTBF7tuMu1Rlu7opIOtqgiKW74XFnhXCWKS17tjXwNjPZClqqBLFSi
YlPlR2p2w0mYPS69zWmlGEx652E6cUt5ldh8JqpC+MKABwlahsEfNox4sOrVLKBvv5lyBdMOxQdp
fyhpPJ3k2ehHqknQ4vBeFgvYyeUdliSe7yPpbUGOcp97yB4EUNBxdoZXbYpPPW+RvKX2AZk4ONfM
Y0OyikkMX/PyOfbGfiaUEh8GCCPjyp9GDj+JV6SOeCn1WJkXdupn5RdtL1fIjPEwpmWEXgnsP6/C
XMI5n5MYggSOL78C8Yp+3AfgWbFkEnSsy6hDu28TExYSl7lUxo3FQccI3FvhFvKLaToTEfkp3+iD
8grpuFJR3XTvQU2IbE+/SZ6BrnLKSx2zGnVdlnEZ2tL5ge/p2n3UamXZ3ZuOwS6gOlhvdz0Hxr01
PaPPNF2JVsOXmvFvLN0FW/KjPz+paBoy6mnboq5xxONpuCIgl3ppxiTqbua4Yr9HR8nPB3Y5s971
mI9AvPWH53HdZ2tUMc4KP+pTQCtJfeoDSY8BDJeOXbSQonSfDyswnBSD2H3t0zRuKINELTpivvTt
zJ+iNpllaDTFKZhhYYKOdGXmv7MjURqq1BifHJ5HdHFVuR9NTBARmblY73TbYQBwnICAxNJShKCf
vcvpauL3zV0bcqAwoOPuGYRL8f4hLSc/ay+jvJ7UF38oUw+vQWjUjMAManydexPkNzkq+GqycZJv
hyDLOlJTGLV9ZT2fQ+prhX7vHriA1qQekNIUVnysjGW9kxehUAbsLfBYG9pSlzT5nid67VBUje+s
l3M5nmxS8d9hpvaOC60SE0Zpfs7UJRWyqYJuIEnSyR0jzKF03xeklBXctGG1Uow2Bf0UFPIYmcWN
GS87OGgtFPJx7vbP0woJuK37dm2NrgRS5XPfRphkrIrKt33tOcTMSAeQHzmtGAVGvCoch1VEx5Kv
ubEv5O5doX9nbgELiiZotzIsKmTsioCK5YmRu3v5amKCy7k9Wu09Q2OIuShCKWWtc5d6KPMf7uTg
b6GNgs2bdtlAZnQebEyY84AC+JA5LmM3Bf3wfZLbw6SKDsbY8LR/siMqb6i56DWeajTXwDvwaY4S
herb/8qvyCbP9HPap2y8eoGDc/SlUaLPtBmYlG81PspAWUC4IO1ParWhiGcFXMG9+6FpypzkY1i2
ibgU82D0izafTyaXwaiK26uZU+AbXt7y42iYpzkYRqIcn7s6djAuS7Y452GwEkuAtC0pmkI0/43R
CeZWGhsFtYVnHFR8/zIMN7R8U/uZg13y8/5V89LrM8wELH9EIWpRPiR5z8Ld82DUSQjX35uY/+rI
2hmeXat+1IdybsKmuTHRM8rw2wjaDr6y6GEDIwVroSZgNuCCYVRLLDW62SGv3l87CjXVN/YDf7jv
RcHxvFRTGjZOn0yx5ratU5K68Tiz/DWieHl5H6uBQRzqqBcP+F89K4x8ExHwpoyRgRZUURqH9VX7
zueUBSaQ0CGwOfJ2X2Hcr/ckEeDe89+ON+gabMTZnROjdzsA10bUjiYX/yQEL3X3RroBdr+fvbXQ
ySDyHFRWAaipN38QkSOeLiK5cVPkgWkcYm4TOFjQZJHVsoLKK7TSyUriY74QYPwfdT5uwSF9FSc8
qlXPQB/Yc+67KwegmuEUlJndGHmvCa7QpwD3JXEMZ4TfOsDvuem0h8gOl0ztID6ZaXaBiU0lhcKg
Jum2IxOdyoOQN8MXpMhRmYcO3RtOOb9yr+ssqdPrETCU+TtjS1yJHB6ShpS3H7N8iw2EnXhkpyP2
Cvfd4wtwcuL0o0Ub79+Ri4yIhjQRVqxYj6Yo00YiCNOCpX1Kk26GiGzXkojWR+28imiPPMkXFU+p
g0dYosJsPZfilNaJyI6EqMPUs72jwFhMqghKcX4rN1ANyavFymu8DZZdwj745jayCD2OCLBFIfpe
jYiDm6pDG80cTVltLFd870hoIvQt4Q6xAgtTOUzmWpcHUoIKUY6Ymiyj1iN/QrBzl58AL5pHFPXj
o5cV8Yr+c90zrm7iXeP+vSiQx83y4PFDnJasLQyUaKEj8eHC9yo3aFdhLIaeJqeMeITzBrphqweU
ZR7EXBIVnI/a4pz+PHNpH6lJwOUYlmvA+pHmFT81HfD7YZBbM7YcKwPX7EqsgH8VjxVuVov047H+
rTZ24qQDYvuyPgFKmQevX/M7FFV9ocauNZ/aZM/FZgWjVemUxN7We6puSykH4B9Dahor3pJSfFlC
V/f20HvwBB20mrVHTwbzOsH2k34M85kDC8gPymRwgOmHAcghVF382rDCk9auSleyYepw/6T17voM
5Aa4J2fN4F9Tx7zjTHZEFt/VzJfAq6aYWwXbpqWALZWCqWnJry0NmaKmlG6mNMy2/Jcx44fdQW7w
8n2qXjsLttb3Ni/IU9PzBSxrMbO/c9OT+zSCjIoy/qsCCBUE7xZwje2MXxI3Zfr9Z4risEsYbJ0O
GyNPZI2AJjjH3aDJI0qSTfj0QDK6x1+65HoqW3AaBYYguleVSN7A/tyTRd6pGHcQ9xY85qtKx0ug
8i5PurcS3/n1zjyMn1V6OIfcRse/wwCxScBMpQnQ7/1bQHJKGsaQOgaMuNWXrROO3Z8PyQ8JB2vm
RX+hydsZ3CnaTDb3nVl1lcWc3rvb7W4JzvGeg5cVrKKYqrP2+0bsoU9pmRja05rDSij9OlLlFFUe
ka1OV/bN2pquBWYeY0sbX2a6KZopsaicu9IjrLTaBnsMmhsAxvgm+fy54Wq5HXSApmA5hsiHNbbm
IcBMbv9vzbGvSCHPN/y/HJ0DkxKwsBfwULw7NRkFmVk8UJrzM2zTytcGpJnDtyQdRMhDDeQTYiUC
pWRd1AyzHucjFcGUo6X47XjWhA/lKa5j+Q4p6wrxTIEJC5VH/NwXuRFnJysvh2A3oDdrNE4kROQV
VqCi1MXKT7d17bgSV7Y+bWGLSzxL5cuGO0GbZCjYR9PJCDhsuwqYtvOna2HSSEb34Sy+IKXDP6E+
jf5FyzS6C/qq8zI+LpxBN07NQC69geOmaEPXdc6D2gVZm2pvgvbgR6nyWJE83EXxe2vvLfvAFgTi
vfFQrJF2CETc1Vm755R9W1t4vkz0udCK+t6rpz5XYFQSDFLB7b+BEcUiJmVZmFw+Z4I/Fa/L4o8r
bp6MDHK+uOGOmli7ZvtpQVE4Uu8Lqf3Qm2fDiqD3KtSy+UQzvFE22EUKq9xctHZNR2X0Go7+ej35
8Yi1ia+lbT3ge3Q+XiZ7/mAkU/xGgyXTtPUl3Tf6IDDDHnn/79iWDP8Bn/2y/jIw4hZRaFaBws8O
2NLPhBjrrGBieXwoJReoleamrsvOorKZomKrkHEdy059yN+HLXonYPWCHmGVmhLq/koIG1TrzqDJ
MEnXqQZkhc2mmBTyUREZ8tfgE4NgPbVYNWWjJjI9Jv1j5N8E9p1AP+tWyigzSelUut2XoyNf/oQo
2e8QX9r1fWW6OUGNQjmYDqikR0F8g/UtGKsmEcDm4OIMUuazO3Hv1At9zTfYJGO1io/AhkqIngDI
30nX9VHZJgZtOEXr5iVk5YsC319zR3/RsXQzs8SYoK6ioJh61fFgvOM6Y/+XyQtJg6km2TI2qk45
MHlk59Ly2tx68m0Jd3g1CakWsODGTvbVGEPFHfeE2D4QHe2OP4kOuSpQwbt8EUgvK6V86O7N4yTJ
YXZe1hWB7Ar4KmrYfZSoHWRjOMEo3EM7qxM6X5fL1k2n5B7Pd3eHTZ4ukYUcaO9Btc7s1Fqhr9D9
EmiLbJftRRy8n24/Epe7i5qEDW9y5mhd6ZC53V1Df9Zj4Ays7gfHqrQaft+w5MhlJVP7JmSdR5Go
zej9cW6+l0b8OgZQwU2mAZZLGEfCZ/g5/q7qX3sNaphMyHqvFEAEMtOLdnXPaadGoMXabdllrxlO
jslk0uqY1piS5bpt2EysL6++L1O5JUwtukyymzC6Zdio/66ychbYzRwyOXoQ3xiQaL2t6zaJBuPs
vmFNHyBxVZaWeJEMjiO6DIoUlsM4S/yysCNbjBDmmFmqjvUf1OIiKvWSbbnqShe83CkriHeLAtUk
xKMPudcSOB8AalP9QACWxZZiN24SnBOU4FI3uE+lC9WxkRI8TtK6qY3QvX9O/YiGGGiiJk1dV0iN
8o24ufeoAJ9mew3W38Y9PWNAur+0KSr8h/o//NpS2O3aNV+zHMBDWPoDdIXjpmX0uL+gtpYTRCuA
Lrm2NVeBF9WpJr1bqW1Ujdb+c4xiaNOkT0gP7t+ZbPYDswggUyDBQx6Xsa8x5FzLUdLiq+cie3hF
HQn/mKYL4JfHKNeHXMxGj0u2Ao9wX8/zbRbFsWyZooZATrU4HFcjPK0DlQmxFDd4Lm7qgkRecC6O
XLp2u2BpcueW8Hg9zDj2NRKOSm91ttkTvt5lW/NfP4Und3aX5DBghw51G/CPJEfZJ4R482te4fet
J6DVGiuMgGUtzRuCKYQsA/oI2mrY2BWu4++TvIPNFo30DygyIIfEliJPv/806/EWUuF3vj2tTuYI
f8lWuQyZ15hJCfs06qSXJPc+fjUNUjusZsoLkzhHda8iUaA28R4vvI2jckcofFU4j/rt+83O3gCo
LAfMabRgHrrULeEqpDue/9SCCNPuS6VAu8444jXceOSCsXyXVGxbuynzF6dW1DIgbiQeJ5gaIQhr
jLtCVm0CfFAhdMBY6ERawRaoQexyiaxnIzEPGYWshqRKVzJ9sa97k4CnCAUq3K8N7C7OvCM7qHR8
JM9gjCLrGTsp7CTQI8NffZKtjoVGJEg5Q5DHqA9gsz4GqDPK/uKSH5B+jjAN4cIf/UWnrLsP7Msb
EALPOoocy8P0gQrgs+0dV+7VyyACtjhLbC58rcLMm57ik5k0yylayxdyUaY7nQ/fJhWcB6m9n1sc
u/1y1tOr/+4HroZuCkQv/VHD/9WtQgNEcOk3xCsaMudV/CYxjp7sUJKWAbtf29zv2jUnU8gXjfnR
KeBspTAPdgWLrMyQnLsQ79PrHzVXzm+6Kkx1S0edcg2b4JnosxjJfU1POq8XD5k0c+Gmi4W9lWJ3
YqzeGnSMv2feQ+34as3kePlme+hr3hAk7kOd+MjLflV0Ljc3UXzYde4lete9OUpjPxgLiM1GTqhP
xmCGOTWcjlc3FCJBkh6GTttxeBtsOHxz0984TNeA9UV8vO886c6LbU53/0+1mOHx6Ja1nLUbRmUQ
0d+IHdTK9b5lhO/PfTf50H9hBnZUphs5u6VDE2chUuPNYNVmOr9+QZNF5Fsd47O+lmMv7VXsenu8
L05GR+5q8B8mXn76OjjYS7rPCY/ZvLO8dknu2oSI3QS7z/LTeqnYw4VQ6r8lleEv/kn7ljNOE6KL
3gp7fW0WnHJZueFgZwI2au2fX2dKL1CMSRcsPNtaA8D7AJyuATrPT4i/fXjK/uQgP/I3gImxiD5E
RFTxMEfb/lJoWL71gnRrI/B3/NaYaG+suxT4xK+LcL7ZKxEqjdNJFqKYRLwK5tuP0afmX537cMUV
ZXvzwhV0Ib9RhGHhr0DH0C+/R0vhsMoy8ndafSNKnDBTQYsTiUnLnCXApZ9tYJHDHsDAxgC3lGnz
s3koQbivjimCDRYOf1p1o37OANkkF8+5+F71OwKoS823zZcUpG5JiqoraXZQugsn7bXJ3UWf7EHc
tJJ8KPsltpX3XTF8216UQrabbI1YjPtO9kSN5TmqTDzbA8vvQ9Ai5EQ4g6nIOW7yrT/wC+/s4/H7
ldXKvrGLgk4tt4xk4MqxeY6NSdJlxXkp6D13YbbeFrszeg0PYRSOpyEnyXlFfISdJjn2P1hNA9xt
RjlPC8Ze/SXHIqtFB+0F3ivxMTabwwLYQT201n3lFfv89la0YTaDD14N0HUUM31fnS8vTYf8xbQM
uVZCqTwn7YWlfnlBK0UjFORNcK5UhfcU/5y+UrZx1RE9EoAQVF/eI9G3A9h6sEAQF0aItZpjihvs
ukLFDTLIUjtgmVEsNHUaKNKYRRnJoMkwZeUshv9D8aHvFUmE32m5c5XLhTAM4BX32wdQV24dS9wR
fvE+kaQOqCwRfMU0UFVQjbZJlU/k/pKlPVxZHYV6DTl5ugeXR6SqF7qBSru6DuJGbbAV9U4zLmK2
vAc25+VIqV9mwNZZBSbImI4fU5DKnuN/f5A11qaohv8GR+/zeECPkln0prida5HzRWsw7amstjax
MgQfsFTxeYn2LS7Thbv0tWWTZxnr1uezChkKF3ZsAZdVfsVNexRfLK1KS+ClNlM4NHcxPUJUDLep
EkxxjIopEocbc9Vr+JmIcjNToX6Z7t84jFk2ccKQ7VGagmeGAI6W9K+BEjaLMok4uHDej6e1qlPh
moUBCPrg2XtgnBiwyrPrHExzAkNj+jhBgBABm41fyiXGyajXE78wQUVbTqOqQsICI23502oZlB4k
B10WfRu4susvKFHr9YlFG3j1LzqEbNxbWvBpCusOA6WjJ3RFar5fie5KlAXQcrOJnAe5jbOYDKcy
l3gf6PWcXsawZIF7YBDe6exniP9RcwCb1kFUemnZnc5aGZusNvi5g0skxKlmz7vdP3PpwEIwPolJ
1uMB+37dDx4R1pPBHrqWRNf33S6QqXOCj76SUjTal9H5DdNFOuAG0Vq3Dj/kEm5dTl5ziafVqiIX
cmkmcHZso1poIf3qvQyB2KhgaqhfOczDamRHAIRdbXMkxVa8YUJZGiPA65IVVzTU+KZuCTL11U50
rkpbmpKO8P9RNl9xOWsTVsocYk7g3gd5rCCtWOvo8A2SQZCkTLMhQF6Nn6woOLvIScIuotO1+wth
KTq1tBNZCUOZ3NYMuO5qQmQdNuAOpIZQOOf2UI1E8j0MO0l4yiYy6i6qDABieo0U77ONUlkZzdg2
b0HkWn19of15NrEGQ7gQJpVrhRseDUZ9qDgRI30/1p3KKeuG2tiTilJnsd7em7F+lnLo3A9exXXt
PZ0yiJPTAFsmuuiNgpqEsRduzMj/ahzh1oDuO9wEsZHXrSAuBxmSJUQXQLDbCrDCPbypt9aQJaU1
NUc59yr4Xm6/T176E3sjLHgVe15z29pvFdfmqhgJS3DNoptnBE7D/9GvkmHDkNPOBLq1n13EoajA
IKb/6QflHxJ3dKf16VW2sthgkQCi4KJZlzQidp2+7i+TxNI4JX9Nr3PJ1NJAyDwNcmgiJnvgN9Qq
DaSE3wYWsnc+ToGvu0NphWF8X+Ty8LbcH5VkCMnnqM/8KENTaifiF2Lb/gJ9OnhnHi6BjH7X0ipe
1KLhgrKHByX35HEKYR9ArUp6hm9RMEGbcPV7RZdeBNcK4jxDnBblZN2AbPrN6YvVSxXbN1jiWa81
E/D0jPOU4oG9gM/ObhuwzxDoOKla3NXCUoz4So/kiUXOzznKwAoPOU73fsEJtcHAgDOLhUUGDcdL
CiuZxqXSdfo1EpIr6tsMskItDZI5zLyZaiSt+7cXYVew7mTC7s0SWg/mXan7Ni3DwdTN5XEvqhpd
wpECQw/x8OKmFvsbtYWByeJYztpNhK0gxRWXXlBQQWxEZoUuLfyM+eKWzM5sjmjoWxKuRKkO3Rga
pPoqjM2dPgbiOxbgCi/GRTSTNE60MBYQ6X6iNrrZQq9k6tgqnpy4pAUM6F+UKjjYm2csxloeQXgg
LDNcvU483AvKsDIkp4Dbpyf0Q1xBzUG7iOTy54mSIzf1Onjty+45abDTwA5nDVIMJqnbRELHYvv9
Ub2l4H1PD8yv0Z1eAYmnLTXjyAYetwtBexUj23Q1YVNSrXjQNkiUS3vzoHjWtwnDEMeo18a5mG9Q
FylZ8u5phz4CjhsXPPAiOkWbaIf9Bk7eLwR5DP84xpsrsExnMjGSocvvpJ6v5Qg7uA8MBKbFdJhJ
zE/GbnnTBZ7ebCYuF9dDink5U+QFRgmI9NsnWpShl/26QSbFEVcixWfsPJ2t16GledM9Ke/Tsqnz
SYhuzhgj4yQ/ojhtWVzx9bmAU7f14S/8zBK5Pg3+3anl2Cr7/R8ePznnOHpXjg2q49+Jh/wxsNMC
qaxWIb7d2lvjzujXsbhP4+HqjU0f4eGqT+4Is1/n3AzjZ+HOltH4gHVkrNmYOh0QHf+L0GyKlu6y
QgvI4bjIMJlXwTAgZYcEiN4vRC0mArJeoNlA49hiKiRBtgXZb7/OMbsKNWACs6ga99Qpw8C5yx5q
4B5BOlGDtX8uoMTZ8oM5OoWJiQq1l6bTP8foEF87u7UaJmpvKlJfbkqAJt075MBfkoLRCR34kG2P
D0rvMvoBPxpTTG54mHawh5fC0d7bST/oUOSrbNxXd6NUAVdFGRytoL2wUKipb6pCfzcHEd3beJqw
u0kstFJ6tAMaQmbRZ3pwVbk1kEY9O9WYf6vdz/+l/kGM4HsiJKeFli/Ai/TajEiyghO92uX/H3Sf
hAFyveGg3wp7EP6OIrqEXgu6MgaCWpU0HSwvE+i/DlPqv1/zx2cOOfnS4Fx3JLjp5W6744f1BXfj
1EU5vQyqdQW0F0e8hEIfLSGFcLrZkN95vAunzFqDuU6Z2o27E+fIGGOBhXtIyyLCdpJC+og+PNeh
KEV6R5t52UcJ1H3Ydmbk4eDhTfW54N390G12ucB+HO8j8sU99Gw8knb1Qtl/H/+P9SYkL50/n6BN
zaRk7+b9ppdZFNZRY4FBXX+TCW7kW1MmKz3818mVQ8+FZn4AsKdPHzlWy108h881MgSaasa8oxQd
iTM+LiQpc2tVQW8WtN2k+q+iO5omL3p2P3AZfROZszP/s+VhPQE/4HW0OHBjnu9DRAfRgkGVa5JW
PpUVnyT2mVRYeW79ku7tkXhzHP+gXbkarzj8HYRTTNs9fwOuxPiiUqBa1zg5igJAL+8Wkimddgv1
KcK/9kFlwwsx797mAodMgxnliZVI23Z1LCHoACcOL0+gl+4BomsKIc94ogQ0Qphq+JSxOif36zIz
MrvUosf++yJLO2Sj0BAbvY/Sb1re9kP7LH6bN7TNIARY8eydhzQJ3ZgjZdJQ0MaUDgegaoQX/NOU
5ST1aMTiiJGcsAbP/3jjhzH3CFOZzIGTR7Eyis4QLPQv7jDHS75vnCsi3LWPZo2WxT7DFomiLAm1
FHzeuOpLhqCiCrCcTmA9WfMUvXRbaCGkyFTj8nVV1+FByAVrQn73SpS3lCwHeIEAqL71b132OG96
xS0jNipX0S3FjMQH2ERRJkDpw7XLLLzElEzzbPYfR/USkps3F8a8X0+u9y1RUn+Cn25JZt5vQ2l7
N/nu3TPvSmBvKuFnn4SNq0HpGUrASvVFwcjyjWkxuGipaO4mVpDV9opLQJwVLn5FQOhHvG394Weg
m0u6J15APg310V/HJKbCb4jgxf0xZgfZdB0Ci+8f55gyhQcX9nrPs+CD0FzTYlG7JM17IWx/nYy2
EDktrfSuvRdunlxngyedKh4ZV1XCSKo+G91W49u39R3qqewbv7sWwzn24Dv4F2A/CE55b+2hV2bF
HAhDNqq+5iVtjRGqd6Cw/Yk489tumGB+kr0lZoZZPOPwNkNEuN7EqUBoBPsZMXwtDy3yVxS7y5vg
r9VR41do0RJqj4GcxwrEzl8z2IVIa9oCrYHmnvTJdiQFOx26eiOSaI1vprKClfO1x5MkY8qb0Osp
bPnt2w2qbF+ygEyS9koKJtHPgYni9Hc5BRMI0pGi30w7HoMhHz6MiX55xUYGXmXPlo2kGe2S7Yhy
0zibBtNtyQhb4g2lPHxT/6WAwgZscRh9Tg485GslvRcPLythOz28w20Mu0xnb2X1zfKOmbvXRo3n
u9kUJrpvUTEJIL2Nug6+dIPj9ilmi4a+3nmd3jX/UGQ0zEJz12DVYtwoRrTPpxkD/LIbfHKOvPsM
CY2ZM4LgCOmIsx3AQDTV34vR2yCiJolu2lys0G1LC9pQ+snveLohQsDCK7ofWo6VoXb8wAvVE9NW
AjKmrbN0zPHTElrh9e1kw6vwK1wSR9YK8HD9a5WgI/w/MUYd4mp1/WwYBpKHV2tRwT7P4BeXrdwX
7IXkcddWXiHzvjJDZba3RuP1nu2LXKPkKJsu6Q85RfbXfnJtkw9n1yyl50QtXTf04mcbkHuuC4s7
F9ckx1VYiHw9NOlopKhxdmUpwVdqi0efhfd+HQNiYfq8ex9WysCtlM4Irl1K0rrZSobeBqRg8CLd
ofPaLZFd7ona5m8DkR+nK56hgqW5YXEBrz66jW4o9IYOYHFL/84OLPWWVVGTxK2zuYlJjG1Lvatr
ImzzJf/zPZiMnOQ/UeuaAL/VDRR4DWlfuwA/AezwcWnYMWggnq8UAvrJpzOJLFfn7luIJf6eZA57
LmU+QjcH6ZM1DywO6YgR4K0w+O1ZnkOSbdaCphnklaipTifDdIK1k/gh+C4X6Pfze/bN/ehWFSct
kT6STte8zx5OeJ8JZXTfybxh3ClAUGUx8GsOlomouEmDIR1prfLKHcNBcg3Z6JjsSY5kisEFKOJz
TKaix9thFkorGa7tG05F0zGR3ANsKlkigLXoJIYpzCbRLv5XVM1cwUD1NQur99cMyqVBg9+JPrjb
Ei+WLH+Wv6bUqU7re7wEf51IWr/WnZzoC3YKdoSmzbMSKUFVltpFutdvkJ9B7G9C3ElZtmVMjTDi
CP8ZiAWgIYmcpSoHHkJhZ1UtYTBVW0Tk/K+9v2yxxm4hzmVop+2Kcx/0RK8xnIzF2mG1n7dh8Y/P
7yjpMD8DGVkO0ZF0Nxw/ap0znM0ZOIPYUxJYGeah2y6kNExqZCGy3c4qDe+lPx5S6kGLDU/QWOWU
70hmaDaU0L5YTtUCxv5M3cQBkXZQj90YRYMZpQerHhhczKjtBV01EmPHw8Ywqe0yrC06BpD7Bkqg
sMPV0ZefuFRF5aR+Edd3CoJCVoiki5+vWhkPmEJUk23V9/34K4J+cXE6XdeaN0AAQMdmn2uGailQ
l1mXmLxBoyJRTNtPpS1yK6KZZGr/CeWE+AiOGU4Omm7MzKN4uP9w9cq0nO4wq8dRORIcpkt6Kdxs
aFWzNLZUicqEKPhTR87DpXCj06YjbSfPYIPC3f6winPAJgXdTJKIBgoYJNErTAgE6Z57frLQbTib
q9G7evViJeFa9Nilg+dHv6zI6AuRrdr9u13Qm5TccAvt+Uio8uDlxLQU2K9dhgELZpY49mptklK1
fdfJAD+7Gm7YyTpm8z45nd9RbW1ggd3DUyyCCLYk4DueLkOJU2+apQOUKLMZutGkPIMru6eY4bK6
6USPhTSD/5yKTS0/51QXssiW6aoKu5kcGuJGuHiCDEzOQpHNqzl4YktACHv0Wiew8mp1x/ypyT9Z
4S/zN1ZNvVe+9houByyma9cq3O95q97C9lg9ne+hNWZy9JWutzkABsHOJFYqOgurXLl/ittBL47Z
9KwUwtkLgGUSn1sR+E2PVkqfJLf6/dQdE5YD6SeYmpkIUNEUxe5jJcG7INw4gSkLqwZaoJulFv3q
aXcLdvYmxdWL6RIs7Fdb4im5/tYABZEkgeDcGSdOL1SrYy+Jk1sjvOstb3ed0Vcjff1CsJreDwSs
XUk+7u0MCUe6/aS1VMBDMQzPFyv1YpZSsc/q6ou8sAPbhbogRNPtx/XfdAP6Di2HPI6vzJKf2U+T
dy8NiExWdTFceoz21NzMRZFJizLoJk6IBssWmfR6AmuYiNWVuj4MXm1IWI5YEp6fd8T4TNcvhG/+
xVmEO0PUIeBGO1N5dK4s1YnZeAVIGE26VOQMjAtW/noetGCF3NANaaezVkSXu1mBN695RXXEGc50
s89Ebi2oX+reVacIJNApFt6uzO05enJdCZlERf+GWPyCiKDeOXPM0qxv7XAWaHpuCY8eHx2Rb2bM
Y9HQEEDQnKZtp/6exLPt+VUcFfFmMMPbw1iqnYzZyrlLlALCmVFdHQCAkEWxxkqlax5E56y76G4c
vIJHXgzLV3l/bhbx+IdtFTYwxAlp9+xo/hfRJ7ZJkfN3NDHe/Q8qFr/itkM3klt10dKeiEc7DudB
SM1A20cgkRgzsPrL0JsnuVDbHZrLNEHS3nq9l/vNPsMCvYpdDoF8wcuotYwccUiCYM5cjmDwF4pD
7afYIIQ+yBzDwMamqQbiHl9gPbPX0LHlSfWkqTzIrzAGCn9QkDYucW7tj6Rtxc7WchVdGFQq5yH2
k91XtJULyzIvy8q/0ym5EtLJxzWn2YZPERUINQClti1OwO2dinCwXzbcqWcvvjlxRJP+5ei5Akt6
ZVKZURniO5ojhZ4TS01iBfR49YBI4zcdOLdZP8JAkZVTUN38RE+jDpErfvipcViLGKBIwfWX6S7Y
dAEkvs6gC8ERoOp9DbYTqlL6megibF6wC1rNC8HcIpCgepzLgm1kBgZsxfu2UNFsfaHSoTN2yeZF
Elb+bhj7PiOe3NBnBhR/6VA2uWVWRd9deqsNKisRQNWKevu6n88IJ7fakqMhMRfALBqHNpjymKVu
ZIyZKhrvPef2HXS4dw+90tzzOIzH3Yxx4KnCcK/+KVNNDRESTe8bSf6+vKHu5aWYLYownk5gFBpc
RsuOC8b8bdlxxzXddgNPjPa5CsYtInNoiUvtbH9IvlYUtJvl1fPD8ki4vW2BF4txtmJtI5qZZ2Hu
BPON37+QMxBVf6wUdQwVoiMhJb8TIy3bQV57SyVnPMxrzHHHsRMBOgbBbd1imJ48+D5zS+kTsmAm
Jq87gdIgRqQ5sMDj4QblApfq0SgEMUJ4/G6r3hnw8ZwOwYkYT8As/6YNVrPvN+vvXw/GD3Ukeqio
oa0RxyVe8APFgDwjSoZpHMsH8sSBR8l11W9RdwPIqnPKhdwL0yHOT/u9ar1noBMbD9nXPjgRerMp
0hDtQGx6A7KeNUjiEUz2ckf3zcFuY/cfXMi1v6z5Bn/yQhOTrpxiuOjy49dcOtisOdhRXcaivZJQ
bw1KsIeV5ra7wJZC/ftqlpcnPYTttjnH/VXHAi78KcjeX6TBrvlGYHMown+5anEAdA43dhD1OMKJ
x2Uh1cxCRk/OgVaa2K9eE5m8UH08cX/u9IxVJXMgzlmEGIvG1UxL14gVIt0Dalv287ccZ5LzcQb7
OtI7aAHmsOj+zW/K63mlImhsogXJgD4kdWnSXsJ0jt5QBXo3jUAYi3ilXceKH9odm+DwFdqioKs4
W5Z6oktvVAdS6uW4Qniddh3NRL80ZFl0oeEr01FMlQXuZoxi0iCYCaEyZVIkqFiT5xDOSyQUHhhX
n5IRVRtYGm+858SlF2AOHeMj+JZUCMwz0MWLmwgWYVtKelXxIWIKhhrkkm3l2iqQkU81WOxyxiwe
RJPqfm7Ii/eh2jbjs1pec6nP2FY+KK3y1Emw3vzMugA4M1jYuuG4rOF0jPzeMX68EY52R5ZEeDwa
FH3/Js5hDh07p+QwMKAng0qVSOr9BH0nBGnaNen+d9+O6587XPw/lmlnLDBvrdZORRsd3stmrUJ3
yL7wCkabH7VisGj8Fjr6ggiMe+F95cgtTQw9DZZkoU5eGhSkKULkeIvFT5I5Iysg/oCvA1fP3sNg
neDAdza02RLaQZjgg7HUV2uObkYdvN7G8hRjAfDXQqSx61hHwnxl2xJeyueW2A+x8VsNSPefvq65
sh3LaT5r6d0T+yA4Byu/UKtzvKvkb7TY8c+J1PvQnlgFtYuCOM1+6IEiCoxuOEuP+lL/ORuBQHcf
OL+kA/5gZiMFWN5R2CnYtv3iMwPboacZa+N6/Z4yv1h/0A9GQYQiKthhmu+8Kj1aO0AWgiIRFnp9
/vzjqFyG3QulUiFLroMSlpW0jTNR5wiwv5CbkPKDKU7TraFkCIyPHKjK7DmrNZsNgrRzB+pgi3H+
xE2CaecHABqacAtBSqIlpJShTAsP8qULL7dcy3qT63RjZ985KYRWRxViwp5ylo6eeav5lZyeLxUC
R2HnBKRj5zsecE/8bAQQshuyzGhhXQDtQV9i5nFJz63JM8cBEkDYVKS8FFyw69zQJ84SjkzIiCtL
p6PSq1lGRHxxZb4yaB34c/TDurqEbmmQLSi2JasSY16s0mdSafAbW8c4hyGYZnsmJjlx28fO+8iw
Gyu6jSILgqI30Mfp42qjeGnzty578aW91Ui+4bfE4pN4qxMQFOz3d0Xbllf8PoUvPejBQL120E0u
cIFf7a0Loy8JlxarGJCtoelfONRCGsq46qTQ08fabwfhBu4xSH+O6fPB0tBcXGmognxbS1HDqQLd
o0dmCT17qr6fTH+l/L245NPbuBzsqllEOxZsBcKesI4YPwt8I5dZap/RJHbNALvhy3e9KOM+1S72
/QO50c33GJSqNcOLmeqzrvSildRukue04TXyqtr+Dwrz+3vB+Txzgn+mwqZkKUqHe8lrOXF4uvQh
kCloY2gPpONgPfANhqO5Y8dzFdWGRXzGVg8C7Y/+yaVKcQWUaODdA6n8JmpYjX6v9dUZKq+wAVD3
ormvESfWw1EWQCbgb2RlzLwPWYVEm0t3F+5OB3b+gLzw0Y++F7a4UppkVPn88C/6jzy2t/N4FvdG
n0ElQlFbTmHBur8jZG94cfmj5CrQ88MyqmjiIMN3xG0tJOSTF17Rn09zenbv60USi3g21O+Y0Opz
5PE1tcavxCHlEAMGZwc5Vkv3U0TcdjKpkuFY0l2XfIVof9NKa+20btfQWqg+O0R/w2pbeN0pB+rt
CHoUpyHuP+QzUQ49HnzDNixY5vtDcHkZ1Q214s5PykRQBzL3F3XlrPyLtgYNdiXME+EQkzIVlYub
6DV4RuaDYJu+hsvZ2xJ0S2UYafGXxS8faRTxnjoo81R0ppnbepIJMkI2egDV/RucwCWStLbfbEzK
JRtCusSbZHp8NrRUq9XSUnwM85M0HayBqhHd4YHdzvwEdIeA4wEQYSnvk5N3P3NgdGzmtll727q4
yBbo360wbVru2JJmvgQ+oUk2RWC+M9wFhmqEKOcTbvp9qWdOwYZLXpKONpRRu7LRjFHceUMVSzHO
iNViL8KJjdmSZ7agRVfHtTmi39rTSsc/UP+IbOshT9d4CoaUV+C054kQJFgOfcfsg3dakPS5+Qco
A4sAl/oR+XxzY8KYPdDLnScbdyEiOYj/803cf+dW1Kth7PD6BTyWOe0lV2/ujtjwNBmrcv4A6wi7
nINAhYrLgxwCYM8kTFeM5T5H0XusevIvBJFOhJDOvK8pdcVsv3ywPye3vd5fD4pCo7MUftxmHQ/1
+lJoUi7j9O5B86KJTUvDgI5e2gf3KR5QJAjUsfGtGvpYEphtTvnJE7Sj37+jnLDKyQuwn70J7b2x
zIg8ujgpPFRaUI/8mwXirxfEtzvRpl++9H7P1TSTXGxGrbCmZTN2q93Yx9wGvdTmJe5NZYw2uJz3
V04lc2w6eiuz0NRJF1zfQFPnl+4tXHWRRh67X9HZ+Uk5E9NLSuDuMOUhjHQ1mgiVpDqegUUHwPx4
0raMaNg5XfFFQHn/gwa+sQKGyJiVR3emxgiUvQNNgUuzkS1qa4W4+BqVfbsP+YrN9uiQ7eEpYMI7
8C7o0cClXYIuamqJKjDqqzldJt4eQpU+rObe5W4wfHb3hTd3/4gcNTINECa5xB+9eMLTyyOJ+s/8
loQO5xMP3l9heEIdWbFDVCkaRT/HrRj5Jyki8atwXuDOYUtvX18yrP3BjKjhcchlUW1QakZ8yZuj
9+HIPMu7cajumbaJtyPyYwYygVepOQpISXyuIifOXnpnAplDx12PP/ItM4l2Tj8nsxgLnwjLeR5/
4zQbAbndhI5JuFdA3yPpZ75EflnyNe+sKivyTL20P8OpU8Q4dVmeJ/V0UFmtFIIGZL2jI1Qa79TO
fDltgv7tmYppYSKTlicaFELL+w1+Z7gQmTJ+vkVjmuXyi0ghrlbvDdrzPkkLTJyZeCcNI058RcgZ
t+aiNIDiU7Pq4TDwdMaYo5mwfboC14K0sn3kfcCxsvxMTyd7RwfZSwhqwS5NgOUb4v1gX9Zbf1xv
fRLA6REkvdDyRxNzEkxbQsL8UdYxM6iWR43QvQ4+XPFR6eDz2RIYk7Li906gp8hJ3YY2BZ27lOm6
jGsCMop4FAl9suyty3FP2w+4dTrck6THqcKY4kaxJYXiI2bZfFhN3jsa8+0mjGvY97xTWW87ZvON
fMztTj9bXu1FlI6BuE3Jvi2fV0OGn7PoSJNxgooNoO2J4gD+gL100qaEF0J0RGMTi1I5xRI6Q+HC
9j1Lnze1vGNy35XhmdwLNlGnEEU8HzLtU8QNKz2SuTP8e1hBUc+XgJA14/mWMU2Us2y0n0Bc1tFW
cqmPq/T4eQAThHrGWK5WN6TKYIQOhj6h2gugxJMJBceNqy9tsA7m7PUzaYV9m2FUWR/o1MIk5rgV
g74ZKH0obfcK8/HpiUILBk1ZdIk3kpTVPglbs/7z6xRREq2TnfqACphaU0SROOTVsVRov/q677BZ
cL6jC9+gGcXcq/coMpk87XPKIgUOPvDf/tJowNbFsgGLquEFQWQQ0Jj4uoaDCCKa2bL8+a0X8Mcs
sTEmWIeqLj3PxshZZDwISIev9iPdS/6mMBQjAoH6cjCFQXaLxMaKKW0t/5Ek7X/yYJYBOxennTQY
sJ2xZG54qIhRhIIltsuFKilbmX/cXuWkue/m1JrYWhtWWjFhKNOaW/O69TMLUtg5kWZI+b1+ONsn
jB1ZP4/ltNgpjvPu/Auwc7vK20HP8bVaahtQhzD8m4IRr47cRFpfIkcDe1z1d8TmcGcIdJgSxLUL
/+3H4RzBvRZgKp+C2PXnnr5NSp/zVSlzqPxFiD7E+Jd0qtzmK6cmRtNZa7h8C1XKUlnUgVRpoZfb
BEZzbB1KdCj04EWxTJax+g72shDC+beT/+pP41P91VBrBTAGV5adowTCjKWb2FgzApaJqr4l7Co3
OskQxyWPLfR2fw+Opqfyjvwg8lbiCTwcikGgHIqnJP99AvWlF5q9vuBp74or9YFM/wFhHtTj4Bsd
PtT0tNUtrlCFpFMI2M7U0Zac+Kwmr4YeIeDj2lJAQj3c1MU8qZTON6ytcqFb+WX/gFosuNvt1rvV
QRZtFIznbaz2OhSN8Twl0q+lHw3bGxdmijzANe049VtCy879rY4WtuDkvLDigjNaSyrPo8NRz/uy
qG9ccke9k0kk0EgOm1NgKAQInTTxAOIKCoKzeeyizVvp22/a41GsmcT5lD2bNJWQZVBE4FMINyr0
g8jXBOJclmZ6Ki/FW6IXZPNJ1AafQac1rW0kErUG1bD+ihU2m2wZsyKyrmomhqbbw2G0+1Rw1JS9
s5xQPXjBaqC0EaluaHnnEdS4n3ZNqig1veGs/Ulpm1gTcdxOW49dtiAsCs/CjZLTyIKwWHetLVHl
e0dELi3tLBtjeEtEC+ZDoJbDBdj1d5lRcqTAy1vDf10BphxUPM3akEgy14RrGmAtHfKxk4mhRznx
QON8bnAAlICJFyZbscfjJD7zep/bta3u9HZA4k3kL26LK6xjkqTo4CLNRQuZGfLmi7keT4MiNoQP
eRRNyLKAxM2SfCAB75JSiX0/lLV3FXoFBoWK6tAlFwQ3LCr06zMEkB4/VzvVZqTHy2BLwzO6v6CE
C3gN0ySdtICdMj83wp2xEa1c8DDODQ3qGthVNZQnq2L25bKkIBJNQ1w7H26MXJSm6ge9G+x7S1It
30f5x8WCl3TGjou6SbqLCnD9U/QPln+uUuCfSeQFLZjKFIvd84Uw9ClAk45yRDyE3gqKcUqJESn9
1r6VziMAc7bBCBp/12oav7J0xQoCPykIUA5dAQ6tvq8dmJzrty/Gh8ALFVVuyUc5ptLIDrFZOIhW
emYIYf9Mr01tMuGKbwVVFOWpDRcs/oVMK3AURwR5hgqXnjNaCJUGftQUzXA2yweyN35nEfqiW6w6
+UCc1WSo4EIe6Nql2Grc8/LjOBrJ0KbHhfqx5bybmc9gSx/ns7SGQ+rJgfm3SBisPc6OEB1F3vAi
xaikN4hq8/AOpk9l32ZdHVM3oie6C75lYw+ZedDDDG+qxsDi0l/8igtvMS1M3sr/f7U5kMJUtEL3
9CvYm7mYuqoGWFCYSEm62BkQ7vwDm9rZxGWZvdUMGrdXV1ui3lnbr09CHiU/383Tpbet4lLcIzUG
Ql8HTSC3St0cA7mdLxGr1OVtvIgBTKqOlc9jWforYZDON2MITIiHX6z8O06cONG83X8HBKNkU1WB
Liza0zvdoUtzjfFV4O+mCDRXWn/5gTLs2YYUz4VEkBLkzkWUY/sUP555/eRrGAztLNQgIg9PxiKy
h9umtxbB0nLlOkpO4oeMUr6+9PYCXDt/8KmV4ALfzQ1e+Nw3H9rnC38ALe8suTuWzoaBBxXiFwY9
cY1Mv6L5qjgE90f2PCqwSEWUIn53mNhqThk8up7g/OLEVKD1PTTTk7i464Vhqc6zd9VE5kZ4n9Ev
3WDo9IbggWqpyfD/Hb1UBKImy4UGAO8ah5NDu7+msmdYIr5OEU3mbAFU6vmHIj7blN7eFjBy37+e
DV/dUXuIdrPAs+cjujQE+MNZwSBTFcvbuahRuYhnAaQC5pBkETnAU12xEd2kyv3+0CbL2Vzb3wsl
8wpeXL2GIu7FadNd9Yl1lZcwUy/OPXBdaWGt1nc67EwYcFWTyxqZkC0ytPT8Sx+42gwEIP2db1/5
AWXySCcCRhUeyrqh3V4ddq8Gwlc10Oz0w4NdVskpO3bJ5C9ChCnVbHpbEn/if1KjWxuh0OMJ4UT8
UMkfVMUFjoXIaF733Q8wRqlCY1x+qM0yZlQJTPGBVBp1ojBXkV13hL3BclnSAGn8jXciXgvGukgU
LQJdpvSKxh7ntvl0n+2pY0SMZVacOqwRI/SwrugUB1JspdLbnGbZTBpCSJ0t5AKAiZcXM7XWP+yW
w4W7ZirZ7CE5HseuIMQ7adC9r4yEf1LYQ2bWyXnbKHFObDQaOFiUCeCvJo/bbeBB7Imq6UXEK4yr
AVZtYMN/3Mm36EQM/b/ST7YNoOtUoOiKxwyrSvoUexulYAosUeM5prUKlVLId3X91FM5ehVpUKWh
rUsr2e6FC6RhQBuNawViSO3IazjgYYupSMDjsLX4x+LaZ3/nhCTQrCznzpsb3P93dNT5cyZUCXNZ
IvrlOU/fM14e1pzmleX8tHaNBC3/Hz9uQHJUa1M0mXSnj9psR+AsrGmYBRcLJk8TT/Lfzgdl0N0A
GdSudt5vUJpcdGTEADhzI0R05dJwVXA1EWAP9lTE81unn+/7Q/a3tLVjXN20nc+GdguNdChqc5y+
TZbnG9irBSJ9wjPOfBdKdOTP88Kjjhk6Dw7wuIMrenBZYF2nTup1+ZV8o+W3v6M2FQvc3F2NtNv1
Q0+z0Vh1aJGKxUIkqDFaEvTlAL6hGm0VvPYQgO7mycjgR571FKQ6/BE+wfFJsoQDym7IEedXOlmw
B8J4NwpFu3hXbcZO06YjuWP0oz1URsTEANzeNVPr0iKuy3bJTMqAboHtUDPKPxMHf8XzDxLc32Vo
SJGYr4ahdiF7XFvIPo291Pomz7v2UylJBW0wNy10zodJD38grs5hj5wL4HxXmADL/Gkd5cAM/zPD
shW3EzaueUFZOVGk1rpPpamA1iXTkVavhiesdxPfKz1xl3IAQvlW8rHdYGxQSFZEyuf3xBnWjHLf
9ackdUb1V3mWd9JkB8s+rxr8ryOhtAQHtS2QTFoR2N4PkXhDWlVLST9V7xEarlHoD0aBhivjO3hq
eGYNUpO+Eh2dw4HHuMEnvAw+2YwBEpmknXdYl014rAOv3a7OlNQx0Flipv73seagdkZE7syzzZWz
GsDGhPv6Nk5QmBWlKUQrTx2peVyoGc2pu++o6Fak5e+X54vahXacazFGAWEsxvci0VSv82zJ/9HF
/rUgD+tf4rNwbFZ/jXtFB/Lyyzr1QUTbAWafKE/cOy3gP6YITg7ruE8XpyRggFOO1XkTu2EYgd6K
6c2aSbD/gYkquX7IXQ+7m/QMqxxTZkOW+gcFj0pv44QkPw3HrCUcxVMDAIW/PSjK9Ev11Ws+5eFz
Maj4fYd1y+jK8HeyC6p8yJ65HjMMwsU4N/4fExnRhHEOanGRJbkLGcEk7sJUQ3fsfcWuN54m4TI/
nd38r3glm7uGsjCegxQAhl7OocrQcHkZfvb52k0iQrUFAPetxpRzO+x6eby/7thxt+1f8GVZLPzp
Rsej24nlygralDOrzDiBqlSNz5xRcPosD720Reab0K5d6NFf/fN6gQ9hEVUVMRXRkiAe5OTXuBhu
DpvhjqHqqN5StqylpNIs14AcbxEqSx2Hl0kGaXvakzR3SbK68ynp3WGE5qjLecyx0Q1mlj2CJ5V0
eBYPqv6yNKJCV+v5pSBKWP/Yv3U/fAeM/XnOWlyj88QDFsDb1klRBazyEKnOCQdXzq19MnsJYvad
F0H+twuWDtbgdD7RtOk/BwjwRU/8wO2fXpWT74cXKdBA/gUfEoqOR7tk3Xq6ARbM3frX+b7x8i6K
uYlrLh2uojWqAXZR+8PQ9wY/rleIw6v5ZBd5kvfZPg36xxS4Gv2mL47HmqP/5ZnfwfmanyYBWwhT
LTlqT377ay/DQIWVlvuoHDDJkQVVJJhDN1Hfrw3zUnYrl/9m/lQyqgkmjwIiVBSoNTS70/bTfgU9
pGp7SJOti+6HfXDQ4bRxXNmt79Ul9+RpPR4UX+AX43zVbo1hQXM4eMRyv7UVP9MoQ7ReesTEvrPE
fhyeoLjlxSexzjA7U3jQK+DSCPDjr0uhynkOP9bWsGB3TId1QDlsRqVlFP3DrpwOvfh9I1z54CBJ
7mte9DJ3+uCmg97Px1E+FAynkBSc6K6xT8Ngax89EYauzRrEUYc5uS18mFyKfSPR2NmMx/AwBg6r
1fmJxC/eCNsTyhG8u1uWK5vtGr+W9siRYK0LX1zkwbmOyg5JZlpPV6IlfbTRvxf3Qd54sZw9RyNP
pArfPM9nCR8gfxlzzCsg74C4Zsox4z+5u4HsYePl6+7PWmOZ1qrqyGdJj6JVRAn+WVlYGajYOTsm
zuaFkRwvp1NsBpmj0LsJQBKMOHQlCe+mm806bspxYI2eNLx3e612/TBexPnluzJI3kPP3XnYGUpi
t4Pv/QqqobHz7hbK8+Tss8w7EoDq74Q801/j5Dyu0qKIFxqKT8FDQJp3OXiY48Psx4tA+g/05wrs
yWtRvkoZ2OFFBu6AXfpSzacq71HT9Ucinm8py9a/YQfJMWFDfLrF8esVVP/o8UHHStHFRJwiGUpE
zfKa1a1GeJpL00SldfsKf+ueMKd5xe0mNfbdnVsG7mKfM8OTKIEt7vPqtYs8mi6PWvQInx5LR959
4bQ1VvAWdGEKwYywUledc+y+803CGdsGJugH3bm8/l1+ahsjZYJ8QBx76t06zttffM60bGf4nxEh
D2XoC6o4b1gLJYUfJKV+4ZDHfWKz/qQ4fpuh5gX5PJII7B4n8+HOqFYhpHi0sGZGpy1S5GHtDyrr
fUJrwknjtm+7KHUKLhOWprLiImBQs91Lo5YEfOfxo9GSthFm0huREM75i5DchMjaCDVvAgtVZ+rP
V1LnOf2bIBzKW4P04ECvCAVW61jHAkudkH2BjwGI5Cw6UuCAZiesSKSz9ZoC3RVqiiN1TwZlyySi
lW3uLUXc7djTWIrDSeYfmMlIRNBh/pqQovXHYrecp6bR2EeYAgABzXWFd8AigUhZgt3UEr8Ts88Y
HKaWj0fCRdaqkpqEL3F9R0Rop4IRJPIsYFeIGmBBYs6slKr5w1UVMhzU8NgdJi8W63w326deuagc
0IjfOiLnF3iX/fifMKt3VJFsQ4DQrfcUCEhGhlEXfm+MrjdC9g5SPnd1BddnTlRzJsaA5RCKU/iG
XZfSTIE+ibNY3+zN5exUN/6OS7J80BqXmMuBLmHz7sTujRW/M4ttS97kEGb2/vCnChCbdJy1HZl8
9UILqGuEJDEFdTVvQta/HWAKIgxQiwP82rOniHATqYNa2x7bEPWP9NxYNt59DxM/pHm/akxO0+y4
C4Un3bO3/jQ5AqfZOdJkEfaA6GoQOgkRopBfhMgBiXqh1iO0DorTSCkVqt4tSTHvzpw44+5jSCET
KLqwIQ/dIUTPjTkAK+LNbHS8xJkTqHQe5ZZTOKEaR4ReaGGl/DXZ48J2sI9xTMT5bcivVTyBq4bW
KSxUHfmKOLr8i1PNPFzwXvck2aJcCoziwHKPVSopwRsGyPs4aDV4S3USgALML2iZGmEpeH7vOaYq
n1kNvF2JhaffnFT+PILT8y0b2rl5vtgCR3DT1TTnZT2CUNYKFKjlQnIsEBJqQYb1fK7aPq++YFoR
mru0/WjX896gN/hYsIPR+KV7B0LiN4dNwp4+3qfum9QudALfUDnrIVOS4NvCfLhApeg0+XHsjmUA
FO+YWLUoBBbZAD5zCdQhY6LIA/BWKF2onU/cE0PDsq7C25Ih1lYHbdbGze2L/HAgYvCezi0GCsRy
LtIU6wP1ZsMPccCXwiiQPeTY5ElHgm12u7SCoSFy9Tnkwd/Ae1z/ZzSI+214zdhzaNpMS03xIHMW
u0rbYHwNyZH1pz+nPpNjf8xNx2Ayt+jmDcb4lLSQ8OSH60+UyzxlxYr+GibZBrASWgurpPmqzDBs
mRrj5ErjSe923TiFb2ar02/5llTjrXVLLRnB2646rZNOPHh6Aa7AfauGKcVL7mbxKFRBw4eIWyRy
XgJqN2GntCTZgc0XvJLdGLIuCfJzRdDboZUVljd8u+m/ZwzsTyX0g+JiLAhfy6XRR1QN4B8KH4E/
ARdmR1e4g5kkHqr+13fnAttM+NGXTpzqLBhcVSeb5JMrY6bh3Lm5orhgRhhabSgV97v6wZDM33WP
pSsCbpHxuT1PFQ5GcnX6t4rpVyEeHx4S/OWj9dWZpI1A/fTFVGflmZDwJ6zE4ItADeCFtC8/+AKo
7buWi5gdirkLIDWQrYFuEuCmrT8XMDhFV0/dP06b+R4jnL6CDna0+CGbJmPtf2sxg9zvCTgPgj+4
Xwka5x/b6N9pmL7aBCezgJmJo231VXkWda7DXjY1NHDk8OouFzsnOKjpN4zlQBX18oAqe0weJ1pa
obUUPCkxE7rL3wCicOtv3/1//rmuKpRHmn3pBSV5WexFr+b//1YOkg/KNZMiyGOM/z5kwbCgo6ge
Ul/swKKWkQhGQM9QEcgMZTpc/H4NSjSW9MMr1G+YqHwLldq6ukboxQOtl3fSFwo2AzDAT29nBwmR
1eNLOV8qVswBVBghVKHCIYtebzgWcootEQ8W/xqsGP0aYVHMKOrPRZCu1rRAvP3ESLdBXV7on1UT
PwtZgstsE5TOKwb2DZSN6v8rPqmjx97MA9tp77eFAgKtC7TJr1o9EmcKISv2pQstQ2MhEzKxcfhd
DVM/d07MKtrnW/A03yVy0RcrRmNq2rHe1W5qf1S+7mxR3sv+o5kJUrja8FrxXg0Xc9RZajVu70FI
PcBvz/V6hubBagzYp1aAGzjEj7u0QsDBy6T7suuw30ku7W7u5kBoukXUofi3kp8zI4AeZaJzJ8i8
QalC4kq5KmPuwAAQ+lXhF++u5EydId2KG5c0jYCvIaXgOxo6PAubjNgrbBBlcvxr1V1cbJwbLwtm
2H65Gv3umfI5ZfB4huZ3vm4fXwFCJ8VeILbnwaz/b4gENr3zg5ggrlAAksk61XGi9bkpicZ4G3G1
PsDV90QQfq2N/c2hxvM7SjPZfHq0UHWTsuRgJqblLTWqCBxBPvUgMTUIv4/QBeLksdwdOluQdEtT
GoT35VjySqRFcJyJrvERo+MUiI2gQ6OQSo/3RIy/AJEVBAlg2NVBeSJTuEfEhG4kcRTnWCaTyxly
wC6CcgLAOkCfMOGnSTpFed9TTPlvFegP3ZSclF+19z9JRxlk/eiS5WzYPEanVaZuYXx7AmqeskOd
p9khotdz99d36IWC+FFCxP4oVXXQNYEzMefTlgcnlgoAsn9VO8kiIt9HNmxCk3wJnQ54SMREkCsE
oWlTR0sI2UI877RdbYNbiso/R0R9vTEVcVOQl0NrzzlGQkwsRpKu8eiXKSMxE0Bp1fI8lKtqYwAe
jT9Le6U03YHZcIn4R0tDtcAlAr942q43+szW0XfBWMRou0X5vb9dJkiw3XhpfgDsQN8NkH6OzybX
4G5hPsd/KfKQXbpdpjqqqfA6TSp+eC66FaQxCOUoRMyui2FHNGNaJNv4jYDW4m/Haw34M6+QGrYi
SqqgFIF5o6VFQxLXfs4DQJG+NkCZHxZIcURu60Q7t4g3O4mVzGJhv0fUML9IhQbNcQGjHE6LQjeE
X2d4qNzsxcgzSdpM6p8sM497dGBn70hPlxgzjOuE9ip7GEb5SJyQzxKI5CdBi5iSzBOW2fpuyOae
TWUcW1HM3C+oerMBuE1im4rt8hozvYzkbXtNAEYrD7Z+B3R8S/qO0TrM7U+7p26lLMuqgl9wvH/o
nIirtNIeejpSQKTAIWR7niQhSHbtHS9fgGn2S6o5PkfET0v6w91JjokLG9co7gJxdqKKSu/kR953
8+DHuc0xowfpDPO+bRSfF2TqmPhYG1pVbaH26pLCBTQXhqyjFSdsMeuTEFpiMbs7m3ylIFjrFcmp
sWNfbYUjQbaYfx/O91g0Ozfh9+uiv7Xjpau+1Oc8IGzIMKLdvtlysmD/2ofdas7nHlZQ2d33Nuqw
RlaE0AH4MVvdeO345zy564j34eQJkNJWgKtEjngk9xzuRSPpPzvItTd6PsII1zzppRkuwcVpCova
HCSNdsrivoNqhwHQamaUqnBuZACiW2EdiEhr6fV60oY71D7Xl+Jse+fFFAwW9hnhrzKRDVVgQVx7
agE7Ku57m3lhoP7VO+zETlxaTASVh+0sVkS4j0epj1AokEL/+zU86a+uh+wdvn8vsBLi+8EiEvlO
uGWKsa5idvexEY/Wlq2X+2LMJE+/9OjK96c55c46tuidHAoclqprFcwIpZF40bv0V6AFjlk8WW9M
wR/wSBwFbQ7xGjZET/Xwt/FiKJwB1AD6p8Tqnkt1HuoLqJ8Q8OY4oGQ8Q3g6KoF//rZrFu9sgQvb
lDq1JUKbFLxHW5wUvHf5Yxa3Xj8+3a76kh/Q39SX+6e6AjSLTTYxqygfidwxvUuzbglxkUh3nrCR
89CRQQYewgDop1KjAC7QiaXRQenI87W8cWP5gonkgp4ebD+DYPc1BXUDj4JlxA4/HN9UhGsRx+TP
45+Ntz/sJYdaG5i3m9maEOii+cBfvJf9MI/Tszp1A70eSyAXx6o3lOBtt2+dvHf2xtaVFFUZW05u
DWsuWBaIoJMdLvnYQ0U+ivNLm+ItWOhkUsTI07CAQEGWV3+u7algZEmtALc6HvKaSQCvWUyo1ckA
NZKEfUfulaRWFoLWsqy9uJoq29oRUcuP0vdX4GpPWgpySVnxjwDHWC1sAxFgg8RvP2CUZDDl6ewQ
ui/eNHuNGnt1k28MpbangbIcUn5UUxl4A7XSxLtsvDYR8crm1Yxo2eF8VUkxFJScctyTVJZFw1Ji
TmLYFSqUnOe1H9LSMv+vcW+1+WkegD7OiVb5RZ5buk2XHC9bXzC5t2Z45j9n96ZlSJ3G1CBg9Kje
23U97OxXGlSmRHv265jFhCdXn+9K/LFyMZBGi77IoTn8tcN9vlMGIpoZ8K/7IMgaw3ABQ1jBTh8p
IA0UWlwHbTJeKQjmdFxapI27Jz0gjdu+6CujIY0Y/RV+kyaaYNSwWsyr/17GkaX7dU3V0JPn7qg0
9PWo8XHy5jDRrojIMFtLdq/esTgUAaWZUYwNDQWnoJbsdN+LpEwSfrE6KO841chEklkRIzu4PUea
5RNgTnLp6/2Fshd+WzFw4+OEFXnxXUrTbfSWYPAKEjSMeWko+CtOEk6fdVpYLokw6zlQsUtOW8oa
TetAE8Dr7VMncKcOyrxwITwEcFnGxfPwGpuaObAeFfC2jHXW8CR6TansEDdySWjLvPpWyYeW9KLO
KCe4yYsjH3z9y2feUdsGlame3VuAmiapsp6juCXtaXt2/HyDRXS4MBJK3vpZimj4ThkHk9yp315W
oN0C2rj0paQUoRRoTW2QlCSvr+0CyoWQS8RQd0/Pq5hNIhNlIQcScrd3/8AlSLx9lva8CgBUg0Ef
in6mY7NRyXE0ZXYgw4Hu9KPtYWCvtL+x8V8oNzDCoctEsmgKma9xORxrqb4tyvemyZzkM4m5mzDT
FO7tRX7AChKry9lBOdqLlRxe0caaiv0GIIrIRsYu7tz+XxzLFugTyLoqrPhzjsa4w9u+Ako5c9HI
Lnqk3y3ytNGvaep7vmzcnvOWMNk3rAhJbP9Faa717Xdz+vhzNm0WjkenAkdPk5Me3/bu/soKX0iO
3xa7VEWdvBOhQwL9WNhE33Z62HqtFf1H9RKCG6UkCCOxdGHDtRa8EezVbhtCowcs8zZXCyBxN7dJ
crX03f6FvyecdlL5zg41/zXDzNH4qkoageMdbaK1V/Oc0sAtxSpQWnlArFjvdhquT2dix5qy/lO9
ewkXgwl/KE9JfGxodRz1V3bkwui3ENaXMVdZw6nwLS9DmYaPaL1+RC3ncNz9yFpNTOvrZwDp+Jxu
Qz5MTYbtMhMuVA371qCYb/eDfxRMzlBKVnAILYHkUrNEvbnlep4AIMfcKA9si+9eL8PqcPk4SKlj
5sgcEGDkjdFyZxf/4SyCj8yzSkLdQ+sLOnN6vGmZ0fAcnIccNmWzwFJhcf0X/MJusyu56OVpiyUL
Zgo3lBAl4Fb6IzdaHzA46ma4N7rN/UhYFlyNiOZzwNuH/WalO5jUy2y2WsleGSSl182RrYzVtO/C
peQZ3aKTUs3Tjz5emPPb+WO+nMsxgzyxkojGvqremxmBwhstD6kyxYi7qVGTo6VtsxGcSbM9Y/XB
qllLlRwVypFz2XHKEo034QIy+SAzvTVRUqDaaXOuCKPSF38n/hJ/go8Rz/a38xSSTs756d6LY7dJ
Ij4KELOdEmtzaTzqx3OB8Hfn+JsA5Sv8WylXKmnMC2xt8QuYzity3Ru7fCtwgz0KZO5aj33Puu6x
h/frV6pdslTGYK5MgMzr3xXnJDcrxDxrhHsc2IgA1RUPq9A2pgfqfsFGx4H9kxv+LI1H6LKkdN0X
YLtMKWnOa6KxSUuB+se6xJkWg0MW3c49SOTpJNJjSQ1K5YQkLf2f4R44EZooign1yxHvj5efdeGs
sn6irWcWg8IGzaKszsBPiBguKP94/r57QQpwTa/C0u1c0mCFJCL0CEIjugnL5Ix3kd6oqsXCCLyr
FyFs1SgGnF9vlnFXOkuRVAznRyQckxNivNHM3k4yBTwZdPfb1n/kDUAT5x7f73vTc1XC9P93B633
olLZQl01YnTWNqho/rRq1vDMjN1YYIMJNsANB8LbTAsAwJ5flJ89yMduKw89qAgoGu040UdevEsG
3YBe8lgshBKqOGfTfwXA0fKmTnmlhY6F8xz5StBvg1WHceo8Xb3QDzME2+B27vq6vX4WmHf7VoB4
NuR0AS/VIazu2IGUeRKpvi83oi1vQPRDKP2YL0IIEWtZH+b4nFtt9CU7Gb8pLnsxR8HXrENxE2ZR
p4zbtBCZH2z4gUWBSEcRDR6U09nZp9YPk70ps95UhLSFdWujMiuXMR/bUfN40w26cvUrWoe3oOaH
PgeFAJHgxmJ1GRhPlIiuB11W3pPlbzkoQX9cmoDqAVdfACQEZKhWtb/gU5JxbV8O/I6HGnb26cwC
l+4aU0Kjgd4zCouIwNrTKAjrLAncczIVwwdwrZAGznXxZf8u15kq6mHXJcvHYToDX4nvWfj90sA/
TtUhh5v+wL+QMIG7j+5obR1eBl3XBQ40I3a9Z3BtdqPOPKJfb7GxwkkYnXHKN8+N8LugHZlQ9QV9
D5t9w/wp9xQ0/UcuxCHAUcvrbivR8BssnhaGXaOOV5gR+mToadgPjWQIgUeJbJRGRIeRmk793Oi6
w6sq2q5AeLr7bB9jUG6hilBvAmlmQ0ixLtW6rDAJLeSB1mDJ2b1CUSYd+KXIXEfs97u8KsT2iT8Y
g74BZyE86EviPmZV4e9jBZYfZJMp+2vTbYsS2S3k6vuiAgvoN8OasJyoWtlmxpfJDBHeMqfFvAt0
l3i3MzHc56YJ780FP0Gi4lIrTY07RYA9EPF5GntVOrMwR7RM3wszDxJ7k5ommYAvLTEFC11aqePU
PxXtzrKHkU7Qmqh4iCxnMS/b0UiRatl8n3dfxgXENLNkkgg6716zRy1EHClkRR0UFRAuxDh3/Wud
HjNLXjspkb0tP8b/K6bZTzp7h1frNFQeOq+7Yhie3gFWKvdtk3ssuK8leeqLaes98BIL9TMnhcaU
Y/m1Mpi/UrHSHksloTUvF90PUdqNoazd4Jg6uXregyjAEOkpxQEndihe6Z+ziFBUQtC6xkfu5Fwp
IfIt7Br4IGhU2rFAJ1wchVaziw4phVahfTlQfr5Gag3xVtNr3vrD8MEZ0zDJ1W0tgU9h2P4xqwI3
yLDEo4eROycNPQTntviCG5h3k1tAw7NZRhsHoFiNA5Qm6oPoDG090sRfiHPJNKB5lR+P3AV9EAI+
w+2McIwCzzLeYdauif38AJlPqz9/4IhVNPSu4g2JgIDeABpPzJznmQ1hAt2pXHmP54jruANLCmI/
rDNRjGmKnDC6mQkU7T4vGZpNXa/Vh3sI3AY4rYLcryXDgkhdfRnPE0BAUY5EOsMPaw8un4/3nMiV
xI/gfksoxMh1PvFtZqgH+4eZr04YLXXLHhEryOtl6sLyCq0XsCdOQ26mlfBDneBe1c5bIG7nqGk+
+U0SXsWK1aR9h6NhVN2FOpeZgki6CbtrEGWGUta/bzcHPxH/xekmwn9cZc5jyVQUvZ8KAytzuaZ/
ist6yY0f+94l5qHNpJd/z3bvljttpH5Z8a+hImkSoA3zPNZwgKuFz34+kirdeDKj4WxJZsO/GpQI
L84YekXg3XG6KyffzTZgZBTbMEiIxyfXQ1YfpqgAbwJTPu20l8X8kUh56DN/mc94kkdbvlgW9vFo
wctzL3b6ERhkhtkRiRAzre2kA+UVpPLoDv+eiYiVoB7Cle82QYI+1/iktAvf0lKl6yZF48ZZQ3Jr
i2Rtz9ARfx2UolVL4Wq8h2hlUQ34V0N21YlPc1+hEj11H7Ye/jf79sNzi3KaF61ARQ2clV1Pt9em
gjTRUPv81bYPoi7bjlHQa2Pd8FjB2hoDlZKuqxbLZLh1M8MUD0NQu/P7ZTemS1JQ9saM60UQaBhq
iXGn6aQhr/s4DDwyW7azuf+opcAaMvkYN3yeqdDUl7FPoHTnHZImdihJC9Jn8ZGygkY1TqPlzuhD
igmBoCaz7aqOGRkQGRCX/Jpi59mZT99O3c/5tl2Sd5y02Y6tzweLRU1PxO4etSUfNiwAG9CIYYSo
AkTN/1q91FmeAv/eIHYcrhrHzXV8BzMDafmOPGJL+Rcq9jEy5tSqDkhQwkbIFGlikyLjDxTlgJnV
C0k9ThPUUGjVC+e/KH8ymvuFup9Gz4kw7JYFzUvcNLUcLcvqFgyHgGe7Gt87eadF+EVJ+iGbgNWu
JC6cZoQblZqP+sm7Jfb6G58Njs6Zw+Lh25alTSa4CkPmWpnnniwQFgVaJddtBIHr9/b4UGcMT2OO
MH0tHAMtF4Pn64z3spr7DpRBhnuYPzDCSFK3GzEI4yDj2HGXzjnqQEL+G1aA6QQoIeqPgQXwvkMz
dz2PJ4wkO5kL06raArOWkVyvCHLiRw+4CaJqHR5FCofPy6K4nX022g+qHNnlIjZvuBuKybmrlnJZ
2U8RupWnRFza3ZRsQVEF7iQJ5aDhBlIcV5VEkKyZp1FveqT1uJnPpECHFR2YeOPgLDYLD37o/jhS
3ZYtaerdhF7UP+TVLOf1pDdgne1JuppuxnPK1jkjIeWo65D1OqCTot7eiDobUgzHtrWnPxjT0OK6
Xl6QDSq7gCZP87CRdRS6GT7LKjKtJrKKvVgQ0IP7QacdFemX1oklfdcA3qzeB4dYN5i1r16AcRO0
GpQBcF5RLnOIIInqYaiU889y8TW7gvYG4xkPypL8TR9EZIcXV5WuDdSMGMEPWA+jdntDon1iq4Zv
57obZ4HRf6eHc45npneavoID4TxwJ7KDlVh+s8vQCZqC89zQCyZIvS4uINvbACMw5N7Le9cjHWes
oYw76luJSYc4Semz+3P28S2sCqXaNqTkNy5Gxfk2JjVtQTLJLw1UMtRVLJqHv4apHb0B/yJPbEC+
+7nTXwLj/+YIQ0v2goAcOw0YqBotPw5cASaKMnjosNkckvUKNf+yOQh3h9vkQ3+j2u2L4lVAg3+a
zk5Wfe8T6/QpiFIT8KeAMGPGEgtU1uZzNV9pmLT4OO8iqF/LUviZ5EV8L2taFYHYM8GxrXnsQlul
zKQjXIXhAqJlFJkLjlb5sOrzzfHjyfKYPHo9fFzbv7xUngl7FLxo9ImjCu4k+1undHr6fp0Von5i
1DoxfH9739XqHmI/lHRjzUe50K38MKDymrfCBpBmSHG5w7kZVLQ4QaetefCNWybyb84QSlY4Zy4k
1GQ8aS9tsch2edkKW9mGk1DG8rW0vH6F+80WrhvbKBA8FWMAyGRUQ/jnFCvPqVBY0f9Ok8IsX19x
f+RcpDMlk8lfp3SiWiyxYAOyIRcN+HmuwpzTN+NyOr0004MMQA3q7JWmYnwn066pwSVr8oMIhIfk
unTNk1jrRyygTJhzYoZpPtia226wFy74TzXpnlPmaCmh/ib6KEBxzzSwlWrYO/zrk0atn8N8g+lP
Pm1FSsMDZbboZmxeVTTnt2LIeOMI9dH0diEnW8iMrnCUF9M1mmfwBytbeRVbcEWPoBBbUIbRaURK
rIzFuphdlNSRxRjTJT23XVFxgnQrMZDagGnVGbivTRAs4qk+vCOuOLNfhYEv/UgvwCYUU0o9HPbu
meggfqMbBezIY3wPlob4sQ+jLB584grFstLg7FC5byv2RwoiggQzZlxvSm2v8yre+oNiD+io+oW1
H7o+O4j2YrVdYezsu55gkr0TdDvOoxyIZsfaRoNRNL6qYpc/88HhGNXmHEdWomMtRe+TkJYNb/0k
sqpjupCd2/sXG7tU3Nj+4eMS7tyChbrIVcypFfXr0m0dkD8SPQu2Mk9yC2tcfOWc1pGqNxLgKxHs
Pb+Tn82Aw1uZKQMuDVXzdAXVji247/l4dNNlsQhdc8u7pNXZGFQ1v6G1LSj1HKcuk+1xfW9EX9dL
DY/K+yrXdYtvC4dEW/iiOvKFsttJEmEM7eywEPbZBBxkYbpjZq/3/VJqWE5GYPI++XAQnYZJDUJk
mJwuMdj2NM+xAolCzFQf518OwXEWbBGZhAYDkNKlw5hprG+5U0TcLO1Vc6LdKl8vO7OB3azmWYJm
HjX7mcYGo6LrOOn2Ve3EX9kyPoV2e+1hovQmefroVrBdFRIMeQKnk+9jfowopID3D3BLzpeFI4SN
nDIe7BHJfdQqN0ztzYq8jqO4+uLb95coXiHHNIur91IZrlbL0CpeYK0saxtOE5F9Yb3vjlzdHxKc
2wqS4qMovGpH3L7q8R2sUX2VFYQQG7A4Wz5C9qhUhmfQLNC3zfzTJAFP3hjxdFtlCpLRytyCgIlt
BVlIUEbVWeQUtKdJVEEEVW/3CV1B0wFEsy8CdURms02GhJvtBatUYDFzHsRXlh0UirZ3dX9Wiz6M
gGPs01ZrdXeNEOcezKbRkNW5M56gzXuFyhLVDDZozXp7jjoQAtVNuCbIN12n2oZpgTn9aydqIa32
Knq4z+A7mcITNdCR6ePbMJrAKD+zTqEr+6B4LgNV8fuUBZdauAn3PTwahDfJARL+6bVaO7nkld86
AqQwg6JC5GzI4v/9SsT+rQc5zlse2lqFzR5/NN9nEpsMti9097Uklyue+Yt4aY4Gd/o/ZNtLFIun
C2PEnnKHg73UX11knaOEt47KHflbSL+Pd9CgJrTeNqH8IhHDHtf6MtA1JlglL8mXHFfXqhnB2I0Q
BhxiV7fB+I7IsqYV70g1jPrN+FlSoKElZEQeW7Cp8nZDnWYVMUE7DSw2VbOdRB4K92BFQdDnRRIb
sF09hPNOkk86DsHkH3xciEyc0pwd5apHTANHTuMZ+CXEMiG1rB2oWRMdcBm+SkegRb3DCQjKYAr0
qupg7zNHDHZvVYgiEsvRA275JtAZK1YA7We0NWO0EZIcmPuHBAnHi8h2vMHkdCydK5r4TBCJJQCD
hBBPn+OqJZopT30VXkIGEPShTIbRloAJtbTNfk/Ffo+EWjKPkzRVdmQKzLBoC0Rn4rMcCkJqvz4E
eKiDlBVO+NpsS056sk6T/AkIh2mfgICiZXhMRI8uGHREMxR0kxXF3gfRHmpY0lT9vw7jSd6k0Lzj
X0aSqCLp0pCqKxWnvNETrvxa/LdE59t5+YvbS6ubmkWHDizVm1OOjhsCGQPl86DDF6VpbcCTGcxx
TAqYRnTCD2IiaW+DZ9reDx2KeGM3xiiJOMNQEXPjGLY7Ybmi52FW0lBDismug0S3PLHwiL16Q42B
3/+KCfKPBoRN4fZ0nmLr2J2ANlMZr83DJrRfS9s9ydvy53ELHHTPuW62ulptDiZUsYx9UAnQgoLQ
LY6flkieFY4KlH5CRrFrelMgTrAw9UViak0yQUSCcSGyA+CfAxAAx0lQP+F/23zGFBVZuvfeScWi
S64nCg1mWF8NA6PuZw9/UrTfbah5uyKHureIJsvZpxI5hlKKB4Y2JjF9pvZi5rOrDBSI75HWzwBd
55ioBCHd4Zz6i2Y5em+EJgdRYaM6k96QB7JOZo2F+qo1LRR6B/0QpvZrV3WNjWiDxiUnzJA98u4S
aEw1yDn0YFG7s+jlkWt6ija/8Nm6+tEVVj6F4J0OsEurcMndhgRMhUrm0LUx0+e3hO7R/NN+iZtE
qNBhEPmgUxIHQ5qWzjsMiLKvot89TIbWiZ377egqtSlMgGqkks9Zygn4ESDoHlfknj/2YT/phCr2
89BU6bdTOrGUVx+suLGpbrcBfapzUDk6AmW8V70WsaZKypUJepW70qdb9TCYLGt7JTaV5NXmYOLo
/4/2lwPsFTGlJodEdNIyk/NI5dv3h19xKTq/GthhREHWS2HqCSzVkVcR2Dtbej0cqh1odzhVuh+U
QMbX5r6RRCtHwGydwwNI5E/C9zUGg7Y7w+XmubNM90HM7jgapphZYz+BEFeC5E1M0HXy1yIMDn+O
xV4HNxQ7UHDMobaF16UCH616reDU2i2InruubMjuMQuXcZMALOpbZgTMMWDkO7W3qEsiokujM/Cq
2KfJLSX9/j2Q+zv/IG6CYy7uIhgZmaonzjkdBBCnfaa0dX+S5gsmPtLcWPJMjCrkTfIzwjmbXO8G
IcrvtQsFXD1ClFNP676Df44DhyWDu3+XUCM+oLKYWpyMzsJK/YTpNMy7ojuzFVNtB1frAmk5o7IP
/mzixYvJZdJ8KcgZgiqzP3Dh4krJz7vxULmV8ZY7PfdqItUEwyls+mrqMCkiKXYCUv9BCZOcbxC+
lLYojEjAFN1OTIJCk/zfkILSsj2VbzfAXBferWAPB36ANW9lqJC4KGYvw+Dt4uSXgDkC/7MBV7YN
usCmKldhI874Si+QP+0J6G2ojuvvRr1BlHY4H62Wgum+zoKJ9XxEz0xM2l0uTV3d6zMQxR8wVRA/
FECvcmhr/LY5vRV26PWl11r0DEAcneYKEXeoNfiSqICbPe0usI7UKbeylkIyjjgzUikRamRfLoeb
ZNHkl7jrjRPhSpfBFNP80E7VftTXzuo4UX/C5Hdb/mtnl250A/C6ycuMZ26pEPZFA3fCcu8Lawg0
CDHld7OFsYs2XBOzgq40A3R6ojnloRz6zdVzuwr1jy+BKbwvkRUcUa5q2CoUYQko/uvKp86Okp6Z
BtwhAwBPTO6Q4p+9qyLFOWUNpP5WV7wQ+dWgmI4qL3JDNiwi+hfo2DCiFbxQQbWI06Kmnl14OT3/
O1hUVJ7hyuxAC52rctSmr8BdkMiwRXjZMr5JtN3dANQ1ofAKZEcU9m5kXekGYirFX1ZJ+9exgDnf
AnrHz8KQdttOsQEYSgIkBgnLDrnDpFoOX3IKzOMF46dCr0yusylJJSepf/iSEmG0ZFMRnTq0HBjx
JMdNT9QISgUGpPsW178OhIi3NxlaG/XzK6O2F0dD6QfjTec+MxoJ8CAfgAwHRj3qBEBpmyZL4ZRy
1ZB0IMjUdfk2J3CpzmPxOEWycvVqSPCmaDSgBSM+sB9NLgIAd5MXIzN0V+Pp9R07WNKO7UCKCHsl
KIhd7CLXK7rmbV6kVOl6O6KjsfVmqrt2I8cdpYST2odEQh9BBPi/F9FAxzdFnUl5ZSca874Q5HOx
Co1FA2jMfXL+Qwx7wt9OjNwv0Fa3UFqkgf8RoZjnsxI2Z/mMsNNjxgOvx2B7P2rnnoDlgwCWE+ek
SCrUspvUU6+UMP0X/ecr0dyCsiVTu0gKt0q8cBx9IffgnXNGXY1fhFH4t2ZPbjJQUYsRVQfXLp5p
XLTAIfKF9UH+QM2eCGZYBEp+KzWhKywtRUazTgtTzBYb6bYAagPdKP8tj7dH3BtoY0TpzMy8Wubm
X9vtGMaNBG+JFWQu7+6urSUK9bTpt3ZkWviCI+oJ01cv4g7RxhAKI4RF14GoPtaHKwXeBYP//lxD
QZ5VfX1DmT62QNQ7qdJW+zxHu5t10e8dKdnOd/cgFEMwULzWjZ6EaIlg+lA+GcIgEQffjqrK8v9a
mCnRb4fx8pNj20MbPpDn6sTMQyNv1+3yDfiYckD0j68G91vIe+QS/c4w9T/2UG1wqjSdiXxUIV6c
Rybs+GDVdiqQoGHp/nuJ8Ci7Os7FDsReCqoT0olCTTrYhi2WSq7xnidcZQuNWnNSxFbJjSfHj/7F
nrkoDf6yu8mavdjLbsVqBgwoqlD/k/qJSaliEqG0I6ig0TTKBz8BuCD4qlmDCobVHeYdOfsg1vhj
pKDt1svRXj4/ARJU24eHR81pD9HwKm6ct+wz3IYY9kJzgSgJ1bKKoCNFc91+UDhfRXnn+Xl/Raf6
6iv8Xdn6QHBsrLumkYHgeQ+bF2DvT+8qD7FqOHE0zZZ2gJkBBUfIZy+cAM92xVkWjRRi78or8Bmq
LP6e1HDK/idhMdf4/ZupjkLKE7yo4w6ObllfCjLgOKlbnTBYywlw+PUsW+5mABJrUTAP3ncajUnQ
rsG0luhYQjWkhs4RrW/AlWvtENFgZ141024a0XJYKE8SeRiRDfiTLI92taRggbi8qDQ2o8ahCOcM
BXfe6pdvx/S3kBozRQw9t5DCTfqI5Ge1wwHr2EKdZ1vPrq1gSwYDN/+cgMCUZfaK2qSqmWnMxhpN
R0CO/Zeh4Mcb1e4ykNgggqyv3qbSPRm3N7Mnyvx9ISp5BG81Xj6YuZmG7B3R+k4v9NV3pKkVK0yQ
BMlvn9AxUHH7aZvOWImhZPmr4NAUScStfFIYp885qpv28p19XkhVXgpBeK7Ugw+7NYqwoStgFAXQ
iM2B0pfNDRbOVBUQiV0N+xh+egqKNx3Y0mOU4/XPYM85IwbRYhJMtVZut4c5FRsgCMm4656GtFs6
rE5i6pSEx8beKlWVjMGO2/F0JeNJvg6G4zK+21WScOPNoFirBHmzbwhIy8c/rxWCLNJ8dNVCdxcl
lLkTnil+OP8CmtUhvAsndg9ioODf/kgeyefXkbKyIbD1jbtAaezmHLmsOK7BEikVx8r2IRsAiD0K
iWEhy1UttwFqAT+5TRMDg2Ot1iSGuyNOPMlSuAKm44jPWDRg4YGbT6V3IVzUrJkBrxWFTl76Tcks
+an1N2hWl6mI1jhtc6wIKt6dmtyKvxkMGx7VuFKEiNjmnXPRHfk3ygYlTMW+xKe54nkL6GrBsT5x
1PlRBfDlcoG0De+xs3Eodk6pjkd5fbcFGq/LwdxLy+cmdpVP/vJJMwhtd7oj59OsQDmcPm0YQ9FR
lG7h1ANBfnPxzxq8sqM7/HQ5MZxpvaVsLXCP1QiIyau64SNMrD2vouhxmgQtZTprwpHcVlR2pZOI
S9dt+uot3K/iW5dCS5gEUERCykNm50mCJli4Yw1mW4crQqW9en77m/9C7guy7LF5ZcckWclZxNP+
bejlDD0jyI7KRQB3Y6AA/weJVzLxmg5jZZwOJUWSA5EMN2YSxe7ywpGDr0//TuFlknJht24Cn5TY
FeJociKdmIJMi8EvBZvwQghi2XQviuHo0HAoEHRnkW7b6qJpU6ZurJrA4866hzqXla2YFZ3L92Xe
tlTF1y2D+S+Fy+iR0qv5VRynOwKvG04tIX95ecdXweCg62PEAqaIlWnP8+W1rLrJhKzEYLLfXwfH
96cJY3jFMeAkHzB6nJ2EXHeBbpP7OKbY3dvpdAdgdTgp9hA+eRPstOXA1vLQX1HZ3k7wi5ZfbwZl
WPvDzpcaQ6ag7VWS85HbyPmcP6oUWzvUaFDcqaWpo09+NTfwK1QYZLrR7vZcl9v5s+amfXAJV3B3
oj5cB2yBFPW9H4yxdMuw4Wk3fNcT44rGaJfmkpSsBzlaqLgEN9izfGIUkXL8EL/unDmNtKgWpF4s
HzCwreRKffCULvmzeF4r6Au/y4T9PC7XG/+l/iL8TGYL2KzHS/Gsdt7k0G+c5ply93PIPtuPA0Xv
EH7BDdPurAalk5JQfvIIZu5oAKkVwS98oSBgmIVRHwiUzZlF5Y50Cjyir0ql/+VakC1XAOemZ9jB
PQ1u4YPGTwIYf5ZdTQgXxysyZPjXJdQrvx/g2OViYq3FIf8ZUEx8sThO4nXGYtlOQ6ERkjkc7Yn4
Gfe4RBVkGFOTGfxgPHLaGGNKfb0lmC0GMNE3rk2+mV1k+2PR5shLd9F8iE09jkWNoRGxWGUe1tPE
OSAeQhMff7p/EOXUAkhRXOtgFp+W2g3A+wsx56i8SNLTLraaY3sMdqpSjxyaTAywJCts60usgcY8
NhZmWV8tkNLkJy0xNyMDcp7u0mlcRoJ34qIZ714bDnPLea7GZkM/CK+GhELFwfi3dpEqVknGTzNd
7Odaw5jUNgLAMDWUKm2EAVzO3rM0vWbFW5BkplDYEjFXUfj1XMe6ggglwZv5oymS34ZXyg9vJcbM
PaBTg+cZ40e7BAtVkW3oHT24yHnkfbFAb4NBUXTRGBBLDsd70REuPTHr7GrYqptCXwtDtPdaGhkK
cpLxIVHl11RD2u6USsY8Iwa82lgm0gRVmnop+XhCUxo64DcgYL1SuCOoZKARWVkx+T7W2aqGCEIj
dkNfV1cu+0rpCosltqDLMaiDmVbp5SX3qKd/OOFQJrfHhjAFk8Ytr5wMekubwD3J63SczbUWMX13
G4azzHRbYoKHT3B+xVJeAcrR560SRvN2bJWnu4A3J2v5/dEk/rshCJ4nJe1Wbak6AYnTKEOCGQ73
N/faSN2k+6w9W7sQW69mUCzEJrXwOawACq5Tf3hVUEDctqbcWQXedczw4wMrmyU3cqYLSUu8Nn7c
0zx9REoPV33nZGHe/LK5TtDrCtQq9ulDxH/dkYXKolOIpb2CmSUOgtuuQNSH1/WGFZAFaP5SGfW8
u4FFQuP+XTAgAgCRUCp7VtZzqwBh8Uy8stsNsxsYp2t+6mHBzf2XgIkG/ybzNMUu2u2TsJ63gNp8
vv3LoKDgB5IxDOu3X7QqpwDF1/F8t2eGaYO17D6DzaZ1zgJqgg/jbfLtldNE6J6hs7YbAMVMoHq5
9BQa8kowQfCk5pQq8bt6ENcOCbD8A9sQLuQaPUlWVdLXMuQAPPw727fS5VQkzAW/J3oPZRKe6rl8
eRxurzxWuS0AuOKo82/i1SQFN3cY6dFy/x0S2DTLJwBanjG72kDxDmCHt5LyNcGnCtXTi90fZ6p3
bxpMKUCSwHT7d5DKsMl+oSveONckDdYv3FDVKeFIygCPZrj9rpE/7EJ3KAkrd29V8Qet0BgnncR8
5W8zbVhQZKYubXmEjqhld4/XWP3RsMPIECRBMr+96qgylxCSrdOCzWC5bJgM92L/+MEw1aG+pqzd
uGHdk9tfYK8jEW3kGN1GD4LUw5vNQxT0kwbpwPosdfJpl5JDOjm4FsMiIcUFnk4NP4exi7Cgr2DP
NZgaw3T8HaDYc1G+lo0U/8Ej1GMCHIopSo2fsNb5/XLovsgdBtxskco6urrcqwg/Amu5+f/uuPpZ
Hc0NvfvnPphj0CEAWVV1HsQmgn1O4gHJjD3SGBevbzU+eGvik5CKj2Y3RechNf7EysRPPGYkMvjT
Ft7hfSCqnGyyyFGM+oxd0UYY9idUvk92cchPSJRIgD+LWGcYL5G3N4bb9yt29gdMN7TJO9HB8YDi
3WAxjrS1/QkXT46pZyk+oAe6vL0RPzyCLZNg0N+LUUQI8fPJx00ardBnQ3BDrAOgLbq0HIzzxtYh
KDDr4l2LdMQ3fCzY6E2z8LA9ZzrpMeLmya4xiW2C+eyF5rFY1fk29Ff4PYr6f3fJoUc/BXRXQ5A8
kGUmHT6edPxhpQ0slaP9yqg0uDbZCYt9N4J8GACyOd2bL6g46SVhDKAJwYAx9N7ynPmiefxNwDlP
+oDNrSDoQiCKuxZQYYcskvVZmz6Wng6L4S0ve0jvKNc/plyTLl85xqGfyOI9QpcYkYSBzPJJxFHt
819Gz/rqyXpZML/eYKLev4vQCG1+6Y4cp+0MS4kSbyUNOq2KbAjwFTJ+WOy5uZWjGZ2w4stJTsGX
xJjnOUe0S2lh8sWDDagHYY608KER0pARkEwob8ZdJlIdp2+ppMGjP1VrWlXxdWNOcnU0+ARsXE6F
WcdrRx67z1OdNK449zx5FJzGOzgIVwMQZwPoA+wNIKTzS5J8yM5EQVyE3w48rmZrju1UoKlTT7wW
BOzgfy6ihlp96ELqkvpp3IKKhjllFWcLNnVVVjRX1ZpDN3HR4n50kZDW0sr0PyefY4oBKEYeGEGU
WCuYCDqVSRQ2TvErjveWeL6hwOWmxUyfy2IRhAu4xJswCHCezCGmUAmJ2Weohr8A2t6lbnXuquSf
K/0dEzZEX/1iMnjabAogIXQ7AzTKNun+9dslaps5Yo54LPBnmo5c1UY8ADXx+IQcS8w4q1yqfiOJ
Z/3nPg/HRiPoVppC96W9X298QAhUReH2SAlGTLuIl226TFnALn1C+ftta/Z3GUNz16Osa022APmb
kk9Gq7M0DtmyxxUn72RJzzXRN32hkVL0COp5UUi7R6fsDUcua1Ia3qgvilgChf4C6Se8SRvKj7DJ
/NL/yvrV+RF6GCXSNI7I9dBIJOJJR/6C/CJe0c13bvd4Ut3pbACgpCj2wP7F0mUbPtb1yEJaN5kr
pUtr/0uwwag2QaHoQFW3b4eRkXHSS8E4lAfdRTwOTWGAkRSTYPQTGK2TPPGXRwJfUamkQOkMiY7R
p3fL57quvL8u+8809V256VDXepB2Muyh4hkwwAphWYpKf4DL0LCnz2j11pmbes6nDIO7kfp/irHM
95ygZ182sC1tFjetq38E/ff/FMiTqWnSMjSgOiJ713I9p9fcXxWRpSHj1yLje/SUHTzOeZnsvnrq
m7m3vR6JVoY4QDdmuBC0BOPca92dod3Uqr9H3OsQaxevJXpIsdLtko8+UPj0a0VZPI8oXIrNTLOI
CtlUskZR48XIjkIrTzXXm+vpuE5XIkeZJkz6BwZx37BuC+5+6Ck1FpzySl1PdcxG8pqZOwJmvIfZ
EgyZ/FMDjwE4S4qAN8lFCOSU65LOiKz8zIiH7iLmLT/1RXDPr794LB2SSCh6Dx7N2VYFNFHNgL84
qrkt8V4mxOjd5wuXKA53L/LfjDPKo8tdK3WYX25wcvWbMdgoUB/zzVj6POKfgmyozedwcBkN7I8g
94YY7HH7LJViX/Bgyunk1NUJf3hAe+HUTDwBoZLX0txc7WoBZUcfmYMvwSkAWKng2oDoCDIQgVL/
hNasSaMfdEdwNHaBDEXh3mAZRAbwKuKR4dM5ydtCnKrxr8pnks1d5mvTN8pt0wMftvNl2/lzDnFb
TRnEtI6ABtSkmzeQI3PKZj8q7sThDZmgYOxUzCtk7X6CKjrOv6GiLyOFAFd63ATCdjg0na7j21G9
QNkRX3TytNPqN8HHNjfQDny9cmlmLyX6bWF4cLVnzAXKiusDHORtJB2NlQ+u4OTIHxLzSr8fgOSw
pgzzVuKuxRFsQulXWqAFdgdw8tqs+5iJLWPvkZnM4EbpuRH9it+z6GvV589s0P1PYqbWuZrQlC7l
BRQvUO0E2Ykj7J7haeIrJG56z0HntMUX8VpCkM5RL2dNqfP2S5YTWo2kxE2zaQCxqOi1ocVMw0Eh
rBff8H88MN9wyTaYa7hCLawGNFG6kxM+aFGEVac2m0CkBHLYnuCK2XWmEyEDZ+/ty80Ho34HcDAJ
qqNzlgIP3Lpwqjo8Yq+l8mj0VbwTmWgjr0JKq+7VLsZnyI3AvjGf0wZLqXjxix6zI4ZY9bG70zsw
G+AYbs/Euv7Lz8k5MAddiRYLgKV8eD+e7I6n3V1WIeKiRC0XqfxxsmB+QSeJfnnUasi7e50juE/I
wMlWk5JDYPZazs+hV3oN+oSadGfqMwEZtnmpxtswOqTKrBLKJ8kRaqYimWvKt/CXl2FMhvnmhS02
CMl6mAQSEaUEXQImwIeWF3HqcirYWdnulBcRUA4mt+tTYi4NzRf5v/XhQZ54fvLe2rEyGS3P+Q9g
S3I4yZ7lUNztJWq3fgoGdsm7msduEHnTT+QzRxt9vImutYXmIUAVJ9gv7rfO438/RTR8ymPoWYcF
wRdcZriITeWyhJ+L2i6TCPlxmEv6nG/t6307sGVTElzrODXZQ1dOIiFAWln8Vt72JQV1VTbTmRnx
O62oNYaAnj7K5n7OIDAmDssRTdZo9OgwIS7KFCGowJiHZP55kZMN+rZc3mn7mtyVM3rv2cjjLT2Y
ku8wuFmJt+MxdnQsq297gxaqSoaX2WUh9A4mu4sbDfG1q7+G4Modr48/s7YW1J59389SsdKhv0xp
wPjhJR+Kmcg5jYFlPhE09NqGk/uWEz3m5h1hm/pb1vePpXfLKMnOaf2bUYQylQtVojWWfKPllotO
vlM5HMJuvuOj4yAlTE5gy8M39xUxHKnNet7zvowQLpLG2c+u/8CuFCfIOhXrQQfUNcl3DVFoZdrK
t0r02c+b+l7mG85vb5lnkc9DwbCkYC5UJiViBJhJKOFeEoZItQdoOp2188trp0RAQrEB/DPZ4/jE
tHugTAN7Xy61K8Xnna4rY2M5BVHQgzj4VHf7jxnQV13B/QoJWobhynmvW4+N61SO0CRMijm8toJo
gnvx9kOdZRCwc6LB/zzZlcoRDpQ1ZpfALjrILKcqvNxOjBNMomcumhO7xo25IBdGU+WIOYnU4Bv+
NM1Ncu9ndbsNTwHNdv9ukGkAP9pI5yilEB4SSqAiam7W7WIm3Ast9PUN4dn9Ybo4eyCh+m3iEPd/
OIWdSuql2t0JxPjXX6xd4oN/+2tdnAPLEmi2ejtKhURyVAQ+cgvWbgDnOsmLwUj7Qj4lMDj/rb/j
/p9S25QsPgCpLLZnKeoJOE4a/xdjdGwtKimfhbvgqtdapoW8zyxbMUBmO1qIAjKuRlQyYqyA9Cn9
ChYfF1TiqFF59N74S/u5+Hi51X/28EWGayD/NbSj9SRs/h2iWTQhkN9zEN7pJ48O2vYF65v6tH1m
ZJs+I5y+7TEaMb3qJLqKGu80k5txDX8rJr8gP+6aE7UIUzyjxP63CHK2kqBYiwc4fJVEd8n4asmu
m8Awl5E/uuHi9hng/f2dtWja92f3ZI9WA3NS+7ddvRavo0EovtXfsa0W9EGhUy9ugMlhg9B/gw8+
xXiihAm56l5+eVp3WSACJflHb6hgPvPg7tqiSbSOk58oN5XBJIxODIVwoml/W7vPS1SP73QHDNwJ
onUtKgTXRb9J3ipiapZqPOT8TDc2YIpZp8Tc/95JfqlVt+hCws8Sdn3m/yNGgddprbyAGzHryeoB
WkEByKG3wePFxajxLsKjHEciOqTMfU4ivlU8v+MqCvOCxyDqgNHUCXk2FhOVzugb0TPkEYWPDM5B
b8HLpOcQFMTxAD/ZPTjHZzaU+qY4Mor6lAOWqqphfBBC3rfLNBkeW6GH66jrnzdwp8d2z2KsYRah
Q+xug8e7CQ0yFl3tv8koDFwDyirqPQkbHsFHGQfzuQfgdeaF2+Q/A+CynNKG5UpcsvG5IRhInzvi
Fg/m8Q3ss0JzpJcwZXfN8ZeEnxmES/qos+BCx/wArlhNXvrW3W5TlyRAKCFAp4uECBqDX2UgU6Ov
P1EltpckrQinDU+cPgAz+hmZssDhWh6As5mQyNilPO8Fd0rg6xIIWj+gyzwqc76tqq9yxvHou1gX
hZi9znh3bXtgVYgGfEwc/6gpDp9pvOskhIFVCmBC4wWXMaJv1j/3RUd6O+MmlUlNLWrg7DptdAUs
XB+N4vthdHqy9ZaH4GVcJKZYu8noL6SrAgteWUw7O+z3h8rK8nVxZcQjsFHXaolfPqVq1T2MtxV9
ModvqhIgRD0zuqPg10PK0FGIl9jnK7gVlHX5SrR+8RbH6jLkiRZP5nLL0IkYLLjymSXA5CXB+Tg0
p7tappH2cJ8r86l5cZm/bPKNpMm6/Sh4atAFLJEsg3jiFkasDoYUWkwrVs2mYxSf6x1fTfrpPZLm
g3fzIcCWS5teGwuIyCfaWkDvi4X4V4gVWqM0bxVSRsoodhkly9mkyYIb5lvHgsTYEN7fT5z/r1B6
+PuNTi4vxwpeQF7596XxxxXLngJMgEwdO9vb9999ltIaHw8GDv+Uemn0kFD7HMjf8D0LEzT1NAui
3WLK+H4ZWZPC9FOtc6A+rrMbz+fH5UCIEdNoJPkvk7649R7uMAU8M1v/upEyiiQUXQkkYyyjs24V
60CL+aDT+WPEvnoz+YV5WiAKCeXKLeCYv7NiKVh8d6k4evJxvKCv2X3PlTmvVxkjS6r0IEHXDR45
zrB057O4EJ3k4LmBVYcFKaTcWST5vCUa0hzMJSTlsHXWEFzyX/lD2NwAdWEnzi5hesLWAwekwTs7
gv1KMW7ju9B3aJc546pUmXB4OEwYJEALi7sU6INTggMahV+Yl4w1wMOcwm/uKtJeG8tXCvc+MO/6
gmJ4jL1jnABx65LqWyZ67m+QzIaQGFIrLta4LWoNFnP71946YiB+UT32UsxF6LCYC5r6mLX0k/9o
i27B3aZAE+he22ykxoddUNcLsLzlkaIX8YXTrKRzA0qjrFLI5sc87HIR7iBPXERkwWcuLiDeAFXW
B/4RZN+i0BRN7+s/tENS9f8nN482Xgp3L2lZihS0IZQGpmBnuZ//dq8VINTWIY5EVtlFCK3AbiGg
bNc6M0bOHyl1RFWw1pDboqx/WuGmx+AwUlb7w4hIE+nNuFCNZmVrt/dh97z+KzPCrml6JbvSob75
EyvaZDVlskxUL0PzVioms01Oec1hQwj3di0FnpmxPC8Ns5K63j6XHRrmPuS7tZ2mK7qpPKXczJak
vFDbky9PfrM1c7/Frx9aDW1w0QyQo3TIFGR76qjl5db5f7TsFbdULpnRt7oGIy12+I4TO+VCGZX2
pICjb4ioP5YgP3EF8Hlc/BRywxG4bY/bOIf0sTTT4uGCWGvVcLy/lkSkunc3lB1JR/2lspMCK73W
ACkfvZRjZTAxwp8WvEWW7FUNn8+tYIB2R2zPXAAXK1T8XwYtBg6LqRYEQ2YLOp7qA74Xbs33mLGQ
hV+bB+iJWJXw5ujPJSif01YRJvgm4q3Dq+eWdwiZ7SNqXrbfMwoS0FjyucZZOTSyYmM8VpmxlZ8x
plfdpQaZEN9bDgWJu4NrGEmcDYXqIPVo4Di+pcOU9skb7Np5FUzs3EbKSztdDhexhyTwy6dlox5T
YMI40880xyau7bJkJ7gAbrucm2qyHDAKKBiLDpW3E1LIVnxW+WzGTmvQQPejP1tXxkst0lfpGYii
WXv5r49g61til5fKpabqW9jvUAIYEx36LaPCAEJ0FF7EVK7erOhYil7XyTY5Kv398GkLqfJ29yr1
r7rAZ38d3M+HPLWbtFJBdc4Z0s7VGA7+GfayvuwGojIQ9f3fCeo795RmMa9M9yya8GMLx3sJBEBM
g19H3RGF+crOOdbYqS8gkSbapGw1SefmVWJjPh7PWk002CMw7H0Z2OcYhXHQACKPRUUEd3oPBfbd
BkQqmlXaFdYnl7AFb5jVdVQIwHuipSTsp6seQJGiSZXApv76K/s/j0cXBtJYyG3Ud45ZObugrCJq
D8aUCqL6vgqLQVw8rpH4+M8KoOL0gQOx7gihgbqYB96ghI5GQarLbZK9I4OzsBAVrPudLT8RXH3m
RrsN7V8F93n6Ph2sLJpED/ATdKjUbMQ1gvpriFyPrptCPn3+E6Lj6JlpTGoNZ7cMeknpN8sxhGmm
PIZz6nRYR5SdZotgqO9Pp6V0xvhB/Njer1PAa7FdsZZkrmq2/xEo/erg/2XYjBgrijsbjETK73HN
tkUH2sTFTjN1RMIvtbrVIlw91YVQZ+uXAUyqctTW26cdS59QqwaDesEhVph6wyhrrwK+S6xWCdHd
dObJjfh7QUuHFTNf/ZR+CdrE/PZ+gqMZRDTqxZ1KwQAIF/nPGn8qfziIJVPuZgu2e9SV9q85wsaN
QmIGvzCRkSt8hHUFxyzavIiwTuBZIlAAkmc8ltKgrQXoqW86I2BWEtnxogV6OQf5DTgKDoI3WJQF
pdL5J8z+Du8c7zB/JPKPVUOGhj8k1Ux8jImjb5u7uNbvW8LWb64q3NU1ZNDywB/jicK7qkKo4DLH
YZHVDpsnIzblhx6fi5ya/mbqg6Tl1PzHjdVIy0SGMipEfcZQQB7Un9/9N3UahjDZcHF8St+lPRdH
XkavyaKw9SGJ5kK9OqwlGG9gH86UT5Vef0Xe9Vqsj9OxAFCRMNEUbx3twHf1cJXo7Y6zO8US1lNu
nPLZaR8dFyL1r1J2ilr6blcx34zSHtzpS1LORrqVZN4piUqlVujQ2RI+6Cz724eshDgYw0MwZeq1
YSyycy/vhnR4x1czloHlsnzVtLSPO63ayn6fF2iSQH4mNha3dah1nRRuqKKl2WMdyHuQOO2j5hoZ
EglxwOfzFK1Gg+ThZCqAOqIOJ3TaaH+1ENSh3w7V5HOw+7Nqeaxu2vj9kRQtjFQBDbDwVHwpEHAt
HzCvslQuOf0Mf6qTCoOXK7+4KSk1B/fWIVEff+/aUaqn6igSbPj2LT2QO9VAWFqNnI0Bpp1BkS8i
VLATYYCLezYqr5RqvGcgS0RctrtWcppS+pCvTR0Jj7vt04Ps8aB1Ma7aLiRnstNxRp19mUHYqQ3N
vPOWU5NNg4u4xmeujBtI9II+DBRJhtUwM3goLyBUqZ6L+koGE4bQL/SzoNgGdR4/Enf1FW+TLa5p
rLlLnVFnWEXhKxX24gYxijRrYQwRnI68/YPzM2clwpte1iLfSl6Gqf618CncL/Ky3IOhCfvNKWvS
egLABQZGxTOJB4C4W0idfZOyH6as5MEFnYJ/cfVQaNdQjxdvDDTNVrYFod0/rYiF6+3waQ9v2ahD
UCfIf4ZPlSgsvo3CiA6AmAYvEMOoAf5NpzhLzg+hthICjH9zPabZvNew8kaM6Rw2slPTLYpMRngD
x6v1SsjYLgHwZhkrdW4uUvD0JE5utCayMf/fM+Hj3QWnetpWVpKB4TX6cdtINUqA28fB2rbR4HhI
RMybHdvie68cd9WucPsMzEBhMX07Z0x8MIw6azHTnBziZ4dXei6Ga/spg9toYhpBCoVcnbNsohpo
EdoHVCRI5nbaE1qpeUR41kGx9UphAp7PmDUXWJ1Ng84jXESHAytpsq/qEBgcjJ7wyEh2aJUDiEPW
Qqb4OGALsSTgKvFXnIKqUJ/nzGMdLjs2P8W0KG5I6ktQPamqyY+rgAnU7TdfvcziFwR20EnNK5/J
EgTjZh+/ov0xlCtC+daZX8gmi0AQDkNTcI0HdjxEv+KA8OO4wLNFAwTv6TsbkriMDOxcFgo+UeHi
kuA2TGAoz3BtIbS/7QAhA7+10heT6/lFAxiBtr66JcV6c8YvvEHcXpR1bAQWABF1aejSAVu+Ge4Z
erIlvoOMv9bOqLX/4Tq9eHDcVFBJgAdJBa1PrE0dxMFdHMoLJ+mjBBKch2DBfzL9MOJRe21Tsoey
5YsB7X2ZhP3Nld9Bivwghh9BwN21qZ31bMb8gkKcfk62r+OcssyGCQcvI3AHjiV/j81H7ZzCfWeV
GZTkzu97uoA/3TVOZ14L3jYITDBSnLRPTyI3ZQTVzFM63UcR0RBv24QbLRXPTTnWhZSXSOneM80y
6GqzNaVK1Mdt3re/8zRD9zVA7N1fwdD7Lrz/In45T+5GXI/MGTpkuZIItlJ7tz1O9x1MZT0pS7ZJ
HxjvKFDu220wbZrY7lPjWGyNL0QsDQQubgsjMAHOEYN080MNnS3OPFrFNXrsYoLIRUlMiVVpuTzC
auP+YB14E7R/iaziHwS8ESNg193Gww953K4VZVyrRhdcLoSHGUMCAzwsXVOodU7W6yJbUTAnKEAT
35zO1Rm64mN9RrOpTaNBjYCtr1PPAIRo9qzW0BTEBQhHo59uYaEU+OQ5BVSyhw6P5a81VLdIyCBX
FwqseVNU+QaH3LbRqR8XSKtKeBTsRg9eAq8+8xUopttfRYiy1elK4u+h3cMaIw74V2b6k1mOGH/P
zmZGjCa+F4OfmpnxFJBsE3RnKsHZxDx+O84tiO0Sk/gMbFaAzueMJ1BPBVPrTZ8uAvySAHO126/E
GgZGZRuBEoL8NbmeDxIadM2d9D8XH/xyOZgNl07RMepfrezutNHbIrL2TrQXEaeh0U3H1Puzg/bY
YKKTVLYYktKlPj9Sti45Wz3XTqgddsig8RYDEQ0a4z9vcKw+ruSeTXGLEWeuNQt64Oq6yJahckk/
Cv9Jlg4THRdSFQsSnnB6WKsb3pNHPjNkDHukju8G05D+CI1tzNB/wKpXTx8BAjWgP+QQNQMyiYtI
qzr+xp8uLkg0wO5ZaT27CHghaZxtabyT9nKlr/FtItIWWPK4JyJd7RAwETYEV9vbymWy7xrvbGGN
DPODjY8YezrOvXpBjlkmzdMEETxqLEPrPGApM/3Gsf/Z4NIPOS8RvAqJw4eTJaJMsyifsvGZABZP
JXqgWbpqElHt4g5fVc8kosivHqiID0azdFXJUGF5qy27SMZSgQAGPGjC1hC/F2CCkpPDxdPTi/SF
MwPzqTxQ2XSlthHFYNNS2A3OLdwvOwv2yfjJ4tKiA9QCv7ulxhTkwd5nI5UwjiBc7l14aAG8CAB3
0ca5VnlgerAZCCMbjgDJxB+P3STInZzT8xewWFXEKe+c+9qR3GEDo2mCnCkkwGCwRB8bg6AD7yBa
/OZQd3JpT0eeedfLmnQcYkH8u6Np5bjuMdQJCXwpYJMGWoD6h4UW5JzzqYtBCSoKiVswm4PSDaDd
/oDX7ynxHjkZpoYvMulDgRsTKdQG+xy5GF2cJrvzqOfGI/sBvifFXH3QqsxFz2ZO/1dyGIVoYpKN
HllhItOM0jaHIDEMd93j5Rh4gYKQaaQxuaCcznl9zu5NDljAfy3thUkUU2y1AgtKDMft+K0d5v69
cPSniNgqpig5GJMrVrMToiuVo6B1Bz4A0V73Jijg546dPceNiO70Xtdwwg0cYNlSFw9hfvzedkW1
fG5bkENMPGmn283pvru6/x7uoIdur2Jb/dVDvDaUurfgioJ8KZaFCiKqSAmVCpmv1DpPYYr8mn3g
31C7KlLmBWppJ1kY5eYe2SMvzEshhNGk1lgJUq+GmDTql62i2/gbf9IuG0JiTohntLbqZ/JoKNbS
x1VSvwnZxUUlNtLce4U84jttU9aRzj5SBZLdGhstts7vQ9a9kbWbkmOfkJh7NXxratHPfvGmX/0q
mFUQCHqD9VzZ/Gci76g590XWoVDG5sBDinkOG9i8u6PU6PKoJ4x2z+KPVovgu0AlrCh4513eiZqn
rSIBY3ohMRzCTyR1SGhYhMMCPBPXAOb/7zmqrDjIVBwg1phnKHahABQrDVgCEOJCJUhMdlh7Jm0E
7L4g+Q7PRl4uGYgRFNqYazDVMjFnDaXKJR1aAxKNnVkCOhsPuo9bupV+lXnb3Xhz09w6+X7UusJG
G1CUEe1Deq9C7L7sQ1v5aaQDFbFhryaPzBzQM5JCfXPFQF6N1ve97fbc2egQdfF6A2eVfqdHva6w
Fdk2NWtDpe6wzwchxT04CZFd9Zx/R/ajp4RwaZ8gKbtSZdsjeboMlLsDWSThgJLJEMyv1zZrh0Bq
eZbqj8bXrzQBU/nOQcW1fsyOwFH80EcAD//yvIGhUjRdPYBxJwTv1hwlI0Kz8WvDY57a2sBrdEHe
J0xXRH5b6puJ9dod7Wso+kgS+VhZjeQXxeLFJ9b02cw1Kp4ySaPRouI9XX3OusUL1xUxEb/n/WBX
Mf61JNdyxzSGudhjGNu38LAYz9tf9C8yslYeU0cw8teqmQjHlI8h6WNdhtu4rFM6pXCg5zUHjl15
un2pBXntJ07xaSvPY+cFhGMBnIoRWaJe4TSo6+RzGjJryS/Ku53HDtw3dMczgaKOf9oc31QvbplE
E8MB5ptFe7FnEEGwZVQjunI13ggX605EUJKIUzQ55tsfO8hg28ik0W6QLnbWb7AzvB/sx8wTzEtk
c1JzgL0pQCviPQ71kUvXDzjSNR+jU9WXAKd/CPQLEhQbB0eQbwtsJFX4y2wrBkRwQs3sS9ehdG6D
NSzOk0sQQ2UNoqDD5j2ksAAY0N49+6ORjSBWgYfAMJpIHJ4R8Hm0ZY2oW3yO3ocLMeXxgEUHT4KR
S94ifFS39B1k2nIjabGfQmVzCks5aT0f7n1u5UDFOldExn2dKHcX1/c7q7tcu7NYRMXpxjyaStAf
fQ2VFW/lrsjvh1xSEn3co18rAJsfy8mCwRos7H22gulLARLEgqqTpYFIrZNqiJtNPqy8SvlKFSfe
u4s6axGTD2rUUEF9I5Lyr5s9PjKDSBeTfFG7q0cUEXbfaWdjSJaGRwtUSB9U+f56itd4lHlYYa4w
nZVZ351GaH+bNfuZgyag52I5qpp/aYYVEyXQSFmlizJMu/94w8uxBsT3nbpsXhr1h5Gte5xt2BiS
7iXQloeHK7ACbZH6MpmDYlxStXApD+fZiv4tyrIjbL2T7Q6TxmOIMklyN1n7Hp9i/bPMb05ieQg1
oYOG7p6shA8RHi4uYF+dOb3A6FHU8J7rZNd4PCJUFN0s0CKN2EtSFtoEoD/RkknkMaydhK0v5VI1
+kIjMW9E4XYmF2O8ErzQmdv4F2x8yZUEGG8ha+4yfhz8jbAAt4o7n5Ye5C0cAcDfEnyBDDSILeS7
4uDmacFUyzjuxnjR+NHwjvP25NQazP9/SaiTelSmhwupnRbRL6pc1kXoKGQ1WG01T0LUU40LuULW
PrcvdIaFh5aOWPbLoff6LvEuEvvHsZ+aAVfcM3nsgqx9MUPyTWDHuq8Co5AmP7BGTUUdMGbRzVZg
QA7OLMD2H1AdpfAqPRduS9Lq6FGEptIxpyhR0Uh8L6XXLtTfud3WfuwD6y05P457WK2QLCkcEKdy
s/h16Si96+lg11Rss2ti3tjLppnRl12kLVyDkHKj3ITC/CEwheY5Uukwtujvm9OLpORjZXMJDfTi
lvdgopgfm5pOoB0l1AiyQlGm1lPGp9ExgBEyzqjWcuCqdkwk8SLM2U1DC4cTqg1LZnPE6bpr7Aua
RBRvXVrAWa8vzzDqAMBQ/AHRutFUgjSIg/KAGw9GRbRyvthfHTFrNTjj6/aadFUJSli8oiqRUcA7
kozoLj2u16meAIqVf1wkxYoHamudRBPPu5HizrmiJVsjlmae5+lhfUqHSrw3ItfULWYbpK6+N/fP
OZ483VwQdxXgUA2PP4c13zmwoS0+bYBGczrIk+wO29XusETXUNtskzleDIvnw7zFHuYv3r0ZHrPR
mSRjqH70BxyGxDt6tWswBEXFP0h184PnvT5ovo7hBfXn5pAPTODkaubAaS9oatkf/mTqC/5XPeS/
FnV2KIiF1jjNhbR/d3zqNqoj3MfplQm+fOT2j62hSeXE8jEz6YIpLaWZkpWj1vt8fuf4dq4PpUWe
6E1ZfXtu0n8UgoshnFPgtRCQla1S4uRcJFxMwkVpft+Rk7Js6A2lWeGAwXMjqwGPHrWn4vlkhipZ
XIJiPUT5Iq+lQ+j2HBqU3R+XhkeeKSrMmB47hMe5iuDISs4g9eShBUqX9CVpgfNBjA7d2JuoOSGm
iISNjzjmy5Z4S2gl85Wm07IKdQZE6xgXCLhI+R2W/ItBecdkZiPeiNN0mp9WauZ/OzQH5szoD1kV
z5ZFy3S250J6NE5c036cNTnfcSy6u6b+peWkuM81ZcmtvIFLwFEyxTdpUo75aDpgLZXjsKwetxma
kY6dSBh2afD3ZXOD+h3mhMvZ6LoZCbjeWggldoWoGWXtUNkGrhjWcqwKw4iPepMOUB7XW5l9750f
Ok2Axt00bp4tjW++4YaHIhnOExBn8Sq4CeHik7eXZlMlLPN6biipYV00ph2IfUBgRIzPF/qFmgMZ
f71XAHQ2ohuvjMW61VEhQt3W3SKEa1a/GR1bf+YqBXfWeKloJBZE20O3qtRkAnq7mdi3VucNSVAh
EXUdp+tHV7wuwXVt5kfXmNV6EczNISww1pg8ZqIJu/5v74zthHzrYN6U3ZP912yBKZMeMHw6M8J8
42QLSTN2f0Urt1k6KCvjGgDxKEKlpfWqH0ZS8IPeIADbVftg/2OAZW15mtbfxgHQC8giiHQcDps5
Wt54NPmVydLzb8xV0Oztmod/wPMnmhynI3AwtLY2tysjm5V8CSJMN1eg6oosg3IFPlOUnOjpso4m
swhgtOThE9Y96e1xhAwEVKvXUTZyvR6Hu55Uop9t3GgvYY99lzhNva/og652jMplTknKQrQUyYjm
VHiCtPbOtzjJIBWsTPNVH3KVMdG2zv8N7g/r3Eamj7srLtOixG4sua5XwSMRIZj+Boh4+USHloYA
s90lYVODfWbQbuA7jt5wqdizZtDD5T6tSFMw7pDZNJdr5hTr5eKWztRS4JfZyW8VR3VJ7w+Tl33Q
deFjPDwo1VGSDTT+QD5EbNNz5T3jCDCQZek5LG7CvD07cfd6vw0j+oCaNu89pwJ78DEfNv6rSf3R
DQhnyggzOEI9qNzvLlGEXMRpGpHUuJh+DJJDvnfve+DqtI8d2+ulqI3znhOMNnhepiLs2tDOzxQ9
XXiqBcHQgALCPmLlx2uGyh7yXVeTK3FlZUe1kHzkqQHlBWxS0NHg57P1wjBffqG5ErTU22jJX7Xm
dC5nBrOCaK69mC3d99qhE59/nXXhk+TDO40706tNbtYsXsAWiEU8P6tQp1F9W5pTFI41REw2qXRe
zQfzgWJ6t+aBGdNVQ2Oau/rQXdDJMugaC4RDFhsTX4rHvIEMXNpnEvG9PTGYIarkRuP5IcFD2mFK
xMrYwslI5F7pbwG0T+F9sQlz1KB6huGvEwoaKp3DArPZq7iXwfN7wfnSURu/AxeDFRC5aKizuzSo
yOWNFE7NjWIBOS0Cn5JKVjNnKIEsvVnlwb6brJ3zCa1zD/AGYXqyB0yanW/HmDCwXsdUL3zwHTbl
WirZF/RApgiOXt8iVKGdmq4vTAUOjImqtvT9kwTnO/Xg0C5uGdE+w+0sXn4TTX2G1Lm2FZZ/X0uQ
vtw1N30MG4u4LPi69o1iFokZTLxe6AUkllhvR+3h71keKnChBTGzLHbl/RWilff09rQ/9VOlfDQw
gg1FQ+UZBbhfXUNRkWgXgqe1sWuTMX23rdJfNTOY9dW+8J5Cg8bh8X2230jSKxErSs0CQJ57lyDY
QyXaIIap+/kFquOenZJ0D4rxE+pRBFfTwJyzzyOAaKEuogtSGUrCBeQi34pWNcSye2M4JIfMhBi0
NIBP/J7hP6nxyb6PrxnFEhLXoQIsvbt1CjYbZrCH+FktErZEwkXIhCxvbuNZ08nkGL7fBxhVHL/b
kx+09QV/bgqchzWGIq3jm8ww6lb5CbZXwcPVdZhN+GvWiiVvzmaohEx8cRPaUoU4COAm4kKZOkFw
xweArdR9Q9JNKtFRKUMpwwXZ6SbLTluLLjJjJpY4udJrDcL9murJfJ/jpEyUnOuU54YhMZJLxhn5
N9wRetcLDOlKmE7hIiH0wEHwK7HXchabmK8jnb3c2vkxan7zH2YrICVncJiUhZZmnqEtwMLgJRv+
DuY6TZo3Cvhp2L4jSgSMhl479Ki6huRpULvapiLfCo2SpNzUG87GxyKvuwECLRllxeP2vKx4wsWk
LMO4psBa8LB7tnyxT5TSKffGPjtuo38vLa9jdDIbKGDDmEBGPHPlUIIBSutiI5SYe3ycDy77XuAj
jhFA6NchM2sPqlb/c4FgrEgKutk5kSr8kj3+JgjUHyqJEpxrhsP6O6ADwEUMc0Syiio2OiXsNy5g
vQzZzvZDqknp3T2J309PVPQnAlyAwfi1GzSreWlj0ow0zgchV8T4iBrxuetdC7T/gP6Sm7M+qqQt
FASOnoSILCmcKQlfBH4qVhrgs4XvKwkxmWqpX1LScTYlH5z/Pizcj1lilZ3lVlarw91q+1IZ0hWV
6y4lQ2GMcb37QPIDBRKX+Bep2IdGEKw5D8qIcIgaHvdhfUc1vYcF4n1AZIjKz8o5ktDoBFCWxt6+
A565b8xdNThmqAJhZdKJt5UuLa+QT4MkpOmta2hzkB2D5kbJ2hOtv+myBGPKpDbqTmScc48l2eKm
FojQRVwGL47kQ6gzgp1R8hkZZCDYskKePwdYJLY7joUbLHNWWZ0WYHtSHGmVEDmZfWjHggTNy/1S
/GwWuZxHxLZMjxy+M46cWuPaoxa5sFoDKjeRSmz1B3kpTMFm2wpFTkekYC3Gq//DENjc9f71WPjP
LxfAAyYI1EmKudNvZmQc6nKkC3jrvDQHT3iQdq/gqj+Ylz5qVcSOM95Ilj5s7tUye0GTSRjlqWgb
fXdiD2UA7vE4FaKgzIV8GbqSydFP0A/2kafSJW6R/Oyw1+/TXTQVy/n4wKowu3hAmC+1YOMP/hDC
htKbyDZRGmaeRztMMEyDJVr1te2Dt7qUsq73klI4Ka6Vzp2A0tCOwFl0FQipSMnlH7fuz9ueLErJ
wK/k9zCoh5rc5erPxs/NVvQagaha7ofK2jyHcF7tGxau4Xkscmuov8szpIDnAPWL8pvD4hmu4bAy
1LDjFWeuxmy/sBDBmcJhc0D9dJ0RMbCZO+jy8IA8AFuZOV9l4RZBSQjoLifbTBM+/nzlzCdiwo6f
lZ5Q+4zE2qmw7eXTgzcKMJ+bz6pQBCj4lVI5RJTnzG75YLGDRZ05908nsatLQXWzHM+/ae0iYaAU
rXvhMZJUG952vGRXoRqIX5sUkOxulOLF9EOU9okbTixLZrptePJRi+kKqbkzwqtxwGsDUlJdDgN/
0yvLOt1X/Uqs0qmrtUO1qvJ6o/avIDsLUxtCul7GmiA6lF6oKhVkVO0/8tJ2qfNUo/62OL/YdSp4
Ps9GlVNxiYG4edprTF3R88Nv59VvrchvmRu07v1/3VNspmGyXnSFUFyK+qK91bPJWElgB86BZFG8
LLOmeg0+u1C3EyV6QWiBusHyFaZw3cSd/w7js/m7maO5RADl5a5SXO63OwRoaMaxuG4vxwEBnIrX
6CttBkuFGrbsY61lD3QtuUnXGLJJzh72Gws9YtQGJ5ANvKc/Z7e5azWo2hgAYbosRgfqH2kjCC5Q
aiiA2CWhC3JozsvOysx1lcqeM/MixKs+6LlvQGgNQ9x1eHD1SasbLvqbnCyaZGrxDpiS7gPIMn+/
O8vavBL6CaSmweYSjfLtO0v1s7n7bqeni8vd5XGzFIGmCw8d+1O+MhUmP/cRLyE2TKhpJwfVxltn
rHR7hdxQBtcoMQhK+qcK20RDqeGlWgPS1VvSE8oeGt7liao2toazDWARr+tgdMS2gD223EzKzv+h
l5Veo9JelWepXyWW3aiA0McL2/7/LS8divwktInooNWnOYiqkac+TUL9AEmulrIYS2vCFohTg/DO
TsWQ9choFxbksbvouRkRWV2CZnCx/yO9wYEMNt4K0r0jGRD0Rn5PoCzKyCjbOobwOMGdilroOaW4
lTFIQW5Vl+xNn/OdXmy3IX7rHBjyuvUuVD1w5+wvnR51PNEieof4uuSuFBMNj5tLLw/uXDMcVCjx
2j/So7F6wFUtWI21+uMumDkvbEb1gRygrJF3vRji5v7q25IFqRhOWrQf+iuUtrh/h/fTr+Qwx+jv
tvFDa/sejuDI5+3+CX4jF7YS2iLDvZT+XW0wSoPQQY66iuFAbtoCX3zhte2e1zx64GOtYV/QnLmp
606+donNbHG2aEdhEEfPS5CA6zEPLnpB9x0dnYRzNrKPsLdjPi8K9kbUZh007fRVzWcwK0iP+LOg
avYbO4BUQBnuVixnaK/1I/4Xv1hsZIDZmY1fpV+AhWhQBbM6rVee1BoTz1Zi97mjQ3+revOeB+gW
hJCEeVDHSeg8JHIQGeEHYM8ZuXsRVij9hSYRVOGP1iznpZ3BZ+Gmmwpi/95Y40Ig69rzMoe47lEs
t3S5dgQUElt81MAtYepDkGyT7Hj9jBWLR04P9jmAu/h49mVFhrBAUaxK923CKaGG0toa84kv779G
60tSmDQWvhTT3bl89w9zeptQ6RjrxRJUTmJykj+Xpz6qNDyp/C7ASJbnHYB7S47B5NyrV+bFVYUs
xq6l4KrVfpU8Zhrf8rMVpR9t3RnM72FwSwxyBvHTpO5zhaHIL4vEtE7WDgs4zhm46+JHHYt9bXH4
fPUCBMslQEXjnhQgOttjHywQdPQsOgrhfoT3I03RfFu4ilG7H2VRcmEF4BAxFoJGiv6M3PijAiYO
l/6nZETjmEk8gYS+5zEUb44lSchTYLjHvxql1tjSiB/XW1YGYT2cLSnVw9pKjJo8v0JWtXFVkdnb
EHHwPjiMbFoCSfxJThanlYsVnClPSz/nY4ViYjVni5dX+HSkJSOuub/jeeAj24e1oUxFV0UhsVUG
EUq+OwhDy2GjVbSyqgmhoNjEIauo8CU4yobIhlLSwhtn+1xpE3sstzl7JczjgAarqotFuxISp0So
yepN1rBPalfDlr9LRheSr+N7Poq9HDch6xJIAQqaCIlk6+RpUIYQQ9Qxzk5T9QTWrBGorMZ35GSs
KBGXMUvnZgQIE3rTrvD1SDAH0HCzP9ANnOdTwmWsndp82SX2+M7zQwyO2alc6zVxx7LctvSAHy6x
zuwGTbcSoeJSV2UtDAfKMZc8RAQfUOE93OPoXsPBVfsm7A7UUcXeFrMCyP2K87/pr3y0b8pR7aVM
fdK2uvQkDM9GYtj5/mqvzFKx8HQg0TeuXwDnzq8ntESCF+QKv/KqmqsQ9kLtKU4/7CZN0C/42iux
qWUeaa5HdEnkybBC3hUkUIeDMbSFYGVZw9auy/HmhM1utXsK4COG+IKcR4xBi7sjY4eRNNr03syO
WCKa+Fh1/hV5t37s3i/eTuZ10iDKPcK8TeN69LUdfDGgAyySvGEqieoGKU3i98eEFO9nJOr1VOv6
Z4aCPkTF21cdhq8+AVyaPr+adRMTCEudZGr0triHJTEZaBcZ5N0JG162wyDXRaSyj+UBJqt+alOp
wCADyWU3nXi0O3OP61J+VLsGe3lRtk2tBvKBNU1fGFd0bIPzDSRedSBy9zWL2XLIq/n1kH/pFdRv
lJUpLBxaBznWtvqjqyjYXUThDYu+KZSIyZeCDqdnT0gZCS28TfWr0OBvGb/0R/7P3eLvCMglCAcA
cjRBHsS5F9zqWHxTrXgxNi06nlEM4GZy+qgiFDeZh+mwLePlFhItL9LkU/OMEu/3pgpoE8cc7lu8
CkbxVRjFjLHzA12S0+NBUkdDcRpcsMjGiW8702MnXs0tD8JR660cVzyDUnnmkVnCNt1RHKYEpfOJ
AgT13G1IVIs8O+wb1LPFt1YjnI5SA14UNZG8wOrUpWtDyZLps55mUa1fyHZvOes4a7d5kv/heDZr
5qduC+Jia/8Y60fYe936DcfforjolgxYr3kuLr1KSHlecwqPS/8J7mUb4XE4TD7zj+k6R9yq0MEO
k5hU1MwYcsOKJkhI1LnQQLVzAAXIufjhQikW+kB+b3MAUBCRL7JUCuQp2+2Uttrbkzw5cuiU6Jng
OC5uPDxBRIZTPnDLAfPQlxGwlskPUHJMdjM3OYtXDlQE0GQIoQrI2qwPnSM7qTihB2NOnkCD6+i0
iDtLSI4oL6M4Qd9hyBPeYC/CfMU+OAPrlE/Dx5KXr9+UNu8UMCi00tYDP67u0B3/LzWg/Gp+XGiC
aFJzbweEEiczKYf1WnVrSfJPwdNVAzsTG1wzHh6iGvbkD1q3T4GspHUqvMKLe6HAwtdQXXNQrAx2
g6D2rEyZH/UYFocRdg6a2gnh0MC6DiMjZSdljakH81iPbRBJBpRa0nbb6/rkHBQfgflTRiKeaTku
nTcNMH6L9XpFv/D9suClLlUTwG9wiFI0j1qDW7f/xI2J9Uz9fETiJD1TB16a3Tstfmb2rjVqtJS6
QhcUh38af2+BALHjGILtvRJImKvFkJqHzSW0gZGQ/M4Lr0vEIUCF+xX8m6GYC/1z4ZAfXsL7f0gH
irQqIwqYKmAn+ffIIn9qyzYPx1kWYNnV51l0YWtFTKhnYv/qPNLiWYH6v4WykH5QTy/DSyGChy8T
eaYM4iLRmAlIi9Hvag4F6OESQl/jjG8LRrreJ3Pg9w2Gr/700CEqkn8xD9+rn8qK6MJ6DMX2RqRD
ZjO2B6byMpwZsOa+JvaxyOnZw58IocIPWrPfxta5PaWJq6zUL4YqKTs5SIqkszYxFIas4e/ekLIA
vnTyFgEe+1NimLklwHDzAe8Ff9aCsWWvqkz8Rn7ENcOCBrCs8J6r+py3hkxP8WmZyr/QM9loCYtn
N34VH5YsfgqkLTVzmCYvB19fnI+l5QS+kZBbUQMSE1SMyn6o+BoKV2xyunEMUEx/yCEPQe1Epz2C
pp8nK96fh0NhcNC/2NAT0kHBouuqFG5hbHcxjNme8q9wNM2fPfdR1D8/xGwPxPEpkDy+pGOPwbr3
hTLdle4+IjMo3PscofisKyrqX4+gSeTQpkmhUbNwzP00ZxkUwiuzhb+ki6B+figU2DryPOHtbvue
ohemxQz5J5kNi1sOwJjb1X/Ht2/FBkKHB7nYIcMQxz/agDpRO7r2D/KqGAIK01NU9EkgQM4VE1LW
oYGEyBPWjvn3Pzt9njRj+Y8AE6P8PuQc2i24fkBNqGB3XMaSjV/M5vUo+gtqZSHHfG4FuRw+M5hd
cHvCuiilxN2RGswYh1HJQ/Ff6xKKKBjFsnEWXsCREdJmfOVYmpP+2+bhTk31VHFt8fBU3AZug07Q
w7qaeDwcDeKiSmUApeZboAeLpcx7ssGgK+8E/TX0nsRZ5Ps+EwzsIEXuCawrKpgI71lW9jsrju8v
8NW914KqNE6G6FHXhkMc9BFEG8jKFGUrdDfR9mQV6bEmapPM5h8X9dtW3AiaW0abx7GcYwui9Fr0
w2VWBtXTcpU6Ou1hL22zNwzSuHMzRr4Tseqlugc4XTaz61R7dc4F7xBakELCQFQk/neWG5SQgHVL
zJ5d7PEKtpomyOMW6YBvxsq1TlO5Ahrrno1Yp0pD2dFqoo5QOY9uZ0NQQTRR0Doch0BRow5G5Jo/
OTYYaHAQgArhFtGZ8l2z1RbsxipGxfKFmw1dT6MNiVjesKYmW0MjyNN7Q7FIlPbz+KB/Ep5T5xUp
g1eSSEANThV8k1d3tan7WOBXxhjUjVELaSU2lof4O2dKat8nxZG58ToI8TkN72uitci9B1mBeZzT
oDzpZCELFCAkaRjZ2mMZIPbqZPzv5/74aJmQTIxmVJgwf6NzA2GEPziMt4aCr3hOSPdWTULiGh9Y
ByDLX/YgGl/73y/y/wO4IHrXRXSQBDaeaqfl9D7dWcMunYSbZsAVPNNNQXfuIQKn4IDlGlVkiSD5
v9RasuxvJRUu6gvVzxkeBJKVFXdNj1B6j4OgIE314GrRkGl4ITixn6JPNubPO+wsMYJ03cg46DMe
uk5+nnD1qzolFS790Alv1RXUBqYmkdtNGwXrefVbgDqQU2BZ5vem4q8foRt59YhKyrfjMCzNKRs2
FSzVC1nhB3CjjZ/jwdpo/NoBnpNsZ9wwj8s8KjvAxFBPQMR2GqHR0JdVBIOypdqjADsLMo7GfGf9
24jdz/dtLEZ/qg4hI1noQnlhbS9mvGAwKAdSCoeJXjaLHgADLdSuJSVo52hfXEzcOfC12OGE+U3b
GcrMfJJa0j1jDGLj8C/NJ6AkPHzpU5r2Ldx9S01HVCSe7Vm75dRWRwWoIbef/+QPvNOlhjqYbJHn
oP5GB9jodM7hjPs4jt6jUN+QOLpS5TWRWqawy3cPyI4bQMfCgkvPXv777aY/r9u3V5t43mNI5kvP
8HRJnVxLLAhU+OYJDsZOFd9MTytEo5pnLGYboViFzHXliRWKLExFGsRR0sZ2uKiZmV9Ouxbo/6VO
a/iU/y88fEpXI9wGuEwIYyAbtkpdeobgOWn0OUuW7gwSeqh8HeqVzyK5bVqUB8UZPybFSBlCzPu/
aCXZjOEaz7RdH3c6yRtVHkDFm6N26Ujthigk1jJOOZJiN60JQTIeqwclb4koaExFh2n8ARZKYvn3
6sx6HajZvKlTgdG8RIspP79bCduYIAYtM/XpqrF+1d6rRqyLUjQIqTpKLvjHxvX7m9TJ2b4k8S4M
gW6EjWGoBl/Rz58jPjh8fF/kQVgtKusMGoE3KVsJhrpRH9ME9f8NRhXndxE9IWdMzkGrGS++aJZX
MJbPY4iWgSMuC8XwpTe69dRXxe5+ZU6M2DxdSNzSS5kq2RlvKCtuolsvzyUR8Bv0HH5qCU34JtX5
PF5gS3RSP8f86owUTYgKS4lsym4zdAO0h3qWSXKW1mb2F34Kyr+zR7EAcj5ttDSUMneRuB+2WDRv
XsMh3mthXNNrudQ9t339sokqLBsSPfEN59fni/eSB2JyD82aQawx8+7hYovIwNiOSOLjrDHPMufU
W9bJRY1qSfKlQRmRsZMrnucc+i0bW7EG3UC5qQS7NQXp0p/OWZITKpzx8tptI5hi0TE2QTJXqUNf
wOOyKwl6CMTRUXJrqQVAexKovp1MvrdtszwiAmGx+juflpVPusixRhsD4sbEw/1HvnrZyQ7yekbB
mJtDqPInvTWnVmxz8EPRttluJ917f+j43uQozxXA3N86ZHB1KZ9fSSAwNgCP836HoOn5AIn7juR5
iSL/nemzr0EO/zbTKzJdEBws5PdXwqqxFlGySvV/BpTiz92QcSwslnMC2w2/DsTPOMAFdYqotwK0
gN6fIXdktsXcHshqOmpzHIn3+2ujpVffenkqDhyGTvZHYzzR67g8WXoSOgC/qb6s612sj80ynqxe
MrjYqVSE7Sx8om5ypGe4UYAQdfteYr6GMNQ8yLO3xwb/0eahE5TQqO9t2wfOQRo1wMjKQ3mmwLk/
hmff0sw2LbcB5pOTPoUvt5xGouKbR9fYDeeR63OWZTLZI4S/OnmkhoCn1UN1bCeMcQ5Z11mEeKtp
HuUEg3fO2KQVa9ln6zNf+WS4NsiHh5qT5DusaQ50havur/8RjIfswNOTbnefcozbpulYOdhxx8mj
qQy8OBGfahE8BBTASnblZiax8qEQ6KKwdCbZzaN10nLXUhSmF1R7aicFgqKPQ2oGCZuIuqzwdIG+
SI3qcD5oMBz6fGvv/rDqHecg/ZUTfJu+J1R/30ZvQ+A8FP07WxVWOI/nL0yV7U9ifna+oTvcPZqT
PmgYXD2/mEQ56kdRF4RB1d51EVatkjBvS7tKOHRkqDSgbgx6dD69Lb9jIhGlHOkgFmANVQ3wSsym
uWlGxrxPJT7eA7ZBLB18Oy1A+v/L57R3BjL5WCkdz4di5LlNM/Oz5k0prsYdjBsIip170sk+XHGr
ahdM7O08uWWChJ9wydqM6VTMK0lnuqHKbAfJaVBFnLqv8xkGWQeAkOq50a47ORQRjItsHkuYRgQE
e1qKNvAOO43m893+jLswsPslIMcdD8+rKlVkjxKvC62LdH69C+dpoAqgoQ5uInWyxaTXXKCrwsGD
fANaAUw6mzD6YwtW4iUgSeI+b9gS9880Hl367IdARoyeXwL0QoPuZiDjpODRikzt2n/cYtioooRN
QU4ppySRvygDHLEBNyLGA3pHu/Hn87p0b9JGQveSnXk7jHMbSHVZv9OsEy2ARMHhxXAnw2NE2Leb
1gva5ECJfKdYljD4oewRNPqTfhBxmxdSC27Gpe+n9joFEONkIdbSDlEWjg/rdME1iKWq1naVtsa8
Od/pxwxTMmvooUv3FwWGBrZrDUfwiHIpaIThVGrk+/1dDKmpFdSQKcYET71YcG5r7oZV89zRuBlB
n12j9EkvkEujzpo+vbHcD4TwWFhZg+JhkeXGBMqkYTvHonvXck03mTfSlHe1ioZ2JUPRVDxfXUZV
+cxx2Zwir7nI1yepWqudovhdFvbq78EH8ImNVqb0LPkNczKGrn8mWp2hljiovQWJEPxtxUgbHb0v
Gexn3/IdUzmziRBnh2enCCLhdQ8j4rqM39a4outkPn8unNlZRlmaTtlpTMuUzrKGYilnEutffxoi
7PAA7/AtgN321xqasDsOFZ05kGurBb7vZT2GK8VXtP56ZVfDfJrjnVf20y80/TlrhAVHLffN4Km2
PYQmIQDJD3+DVuzWZtaKHScm5wzlBA05WkCpaK5To3fjuZYOefiklYT4BVyVxp/o62vy+CA0GIfs
326AU1qxqxfC6HO3FKWitAsY0Cv/pcwoLY/bOFuciH+pRqqYnxbYYVoSO5pVfeuzJNJ6eFOgfFmG
HWK3+dyNfpGs2bKdGolVp3Vg5ab4yuzCe8bkhUCeH6C1Kfb4/F/eyIHAb9EPx0c41r+y3+aVJJHk
DXSrnDV0Re4Bij//leBkbeBvGNmfoG0aeRToM4Vuo37Q2wnikm3QTNQk4Qcr6Uyqa/pFDYinILwL
f89hojHTDWZn7ZaLRPz67LAiQNUFfkQiVBYevGefJQMRX8M85MyrCzaP0tHxaJce42xa2LE6aieU
LQKmRPRzNihQeHEn1JZz22SZJQKThx6BYQMIDJe67mtTL9KlCC45JW7DH2raaRoYK9SkugQblI6M
bevqAB5IBcJ8jlpRc9z8gzKz1N/OO036fDsLx/Y9g50mXfmytRUKeicY6znyoIEJVA9KV/0MzCuz
Y+oOBCQufB5iDR2w5OMFtpOYtGz3tRYuU1GNmSEvPLlDazbcWBUSWE/nDqfRtgpyfG2+vHYgsfav
uFgyWS7XzPZKRz+jX3n2txT0QBQNBxvdTxP2hdecatrjbB3Ztwyai6JqFFYGdcTIH9lMOvpqY+OS
ccK1vIgU+CHrX7U0eHkcEJxjSxLV6lXzoEbz7xB91CUDmaKnJF9ackDn5EDTLrT+fFFZtm+Dyyau
6wI+fMmiaahIxC0L0jnIuPoQIKoXF9bORBCTTJy1Cejq3VP8WeEfI2QsIeLQyX6c+d7mdLr3/ca8
nnL6sPzIbEoOIoMoO80aY52HLLUoXu8cJ3w9gpZGD7k+BNbUs3723vNZ6gONNeh4p45wJrBA++yX
R+K8qeTMUim8KHHzLYS2O/CIe+DcXFOCzw663rGPIkGRULY7CJb4X1ZmmQSwi+bBmBplTwJH9Igq
wq/95KvUKt/6dRgA3eclI/odZ3lL9U/beRWq4xWnRhLALfsijpXGjxUhQBd6e7RCw+SzFXj4kof0
SNYy8UwkqcEgUIy80VQME8726EZiTVT/p0/6j/qhpe5MKxg/xVw+sAU7cpG3aLCY1bvhkCm+XcTY
hKn37kxjuo8YT97KLZ95DHDFgRLix69YaraqIxCiOtYdzkmqc45E53wwPiIhSoB5czbJiMUwXfdO
Kq2qH8ydkp7sBHjyNmprcxe+Tgv8qUtSMdgMdu5KdLQy6UHRdXvFq50Pwy1cORZtoSh7vXL/33Ts
51TXABOcwJGeLA27YdvUoJCdLT70+X2uIjAX2gv8/kCPPK5CL3S0nlz+iNRqF8uWm/6K5bT12fG5
y+CbwTNYDEPzhjBnDVqq20gMN/yAImTw+ojJmFB3WnqKR8CxVWs2rOp8ZMrCmxsvMaHgsmYzijET
GpyjvXMiZP6oOMOxD2nXAoqPiyKIQALwtfZS+BrVWopUBRvEl+1FVrGvOyv1Fsvy31S3rcfkqcSx
o4P/wO3wnoILfAky59wY1ZZG4i53JQbwJTy4Hx/4NkTxC2doXIuEFnot3Wth7WBLSEXTcpvqZkRk
67EZnardlHIsaCrju608K28LD4rqkuco+Obf9ucXZVfJxVxO4h7ZPzIweA+3we1qUfbfm903FAu6
fGiWILiV38PcVP3j5VOVxw3BAca+01ZUxFdrBDauv4ZmLc5JvBqLbelJKyU+VuL2EKcl8kKqZrp7
5iHq8vykY832xO7ROxT+ZLm9/CacI3i75eABQBEoM105DBMDY+4lgFxs70RCBtFyn8otizwcsVDH
E/7v7ekVrlfYVl3jszUe+3cl+NLG6lsGBZy0dCD94AhelcNpvfnqYjFkU00SaWUPON4GBC28J9LT
cGeIn9gIwM5l57QPQ9I+lFIjznyyA3hHYKIhBjM59ov+t9PYE43WWHVtNVjGb87+XDW0I6ePAu9G
2xa800v81FGCzDIbHi4GlVcCPuPNmpY2cAO/3iJK60k6G+Y3J8w39hDXLcV6ivERINkwvORBiX6f
yFJSA3Fjsf/QS5BR/+mlBfOQiTWMOmPdLUhP2gh1PVUfY3tF+niuEoDH7UWu/XI7JzBiEV4IJW9n
g8ebwSlhPgj+aU1IApD0XtkKKVIEM8w1iXR8/0pm2cv6DjOzI+MfxiaqY7Wu81W4QsHeFwkk94aE
Xg7kvL6pz7nbYAz3OfEreD+zoZSHVvPuwcuj6xPuEJWMNiBxN/jpn3W44pPUWq9lpgHZmBclCU59
2JIodEz7AUMvDi5G2YHOW4412nFtR5S345hecSrlo00m1FMPCqhK/BTFJQswKx+X+B/maCLEj8iA
6a27SiO8HE5XUCKhHG0A67WpZd9r3mQ2Ux3eZGMtEgChx7q4N0gDWpiOwlwlVgz+Q0rvCH4R7VTr
tcyqcIqzHKNuvIUspGO/5i7rpzgomCba8Qrlx3FjRrmtVEwqTPMXkp/mkxj59XNtU/bTx6CYfjM+
xfN9L1cl7FyYcMsaEL3g9m06m/kX6rCWxPLkT8qQtF2pOEZ3s3qGDvhEDSnEv80OJf+swXrovxeE
c6inJtKOw+YKO5OYd+b8MWC377gfAoEL6HjKrpsSBRDagCXPp3+PcezYZUMLjijqjnVmoNWhfX3e
G6rM7I1bDOFIf5+5ir7GbNMde2HHagL6RmV2HwkxFsXivBts/OYafgDL7GaKotCEukHZC1si8W5K
wVbk+ZI0O0R0nMnAr1iTGRZCs6Zn1X4hwrxXeeHKclfv+C2E56acE54LOq8jSbVCEfO2zKIh/pUK
ojdjyWsSphw1CsNlWqDFd5cYdOw1Z0rcuxPykgG4HC8W68JSvMgtt9ZbEoNObIuRLr+s8qsJchnb
p0IkM2Y00Wiy8ByK5rwZKksi+vpKrT3kP7zoY/m0EsjeDSXDdaDdWQ3cJ+OgEZMKEQt65nkqB31p
R6YlQOpZ14oRGzsKf+QczNkrP4uoIsIpAZ7NjyWbwrNcdLPa5Un0nMDe05yiczUM168OPr6Y51WF
tBVWzOwP56KRDy0KyPQPYpz0rmGro2aBeLwKjr8kfBdHaKAAzbPpb6wsnqwsYvma8kp6P0d03AIM
JhA4uxFHtjwXTHcy6EKR4A86Zc4TZDBWVBQatBIe1WmocVWSUUIv9gIhvd3nG8y45emLDVCCx61G
mraq6651uAu2rTNiFCzrNT/fStI4KgjcON7OxaZEDvkgfiQKw55mXeOjrpjgZsyCJ06uqPREg+Q1
/6olehSxfjEe1mGyvDela0N/Dsa9Ks9lulnB19MPM+0T/rFWRkVUBJ+A/euyY1fnB8bRvKhWqGvj
1Mv10mpz50AaROpg/Wusaq7LocylR/EKQjUyZaUve68dc1O6iCK+X5ux2QugPMBiBCs8staI5nt3
ckbaWCeHuyKejB6PkupmIdTrNgaj1dzCvIls3TZdZ5dfacUCtsl3475S873grEYXUUjQUl7loOfF
8SnqSmLAa5oucxN+8yO53JpWNX+RygSjdQJzhvg3jitfH4UIUyLtqcLXyqFBQV//5V54ESu9+zz3
T2+tSiFLiglJqlo9/dAkeeFvki3GDMvRrVKi5AKO+KZaj7fhZaJm6FPfloO1K3dl/pL+6JCfPaqx
UML2zQ7+KTqacpspDushf/EDe2M8+/x41nv/jXzXQEtlpj+fvKuH1RhGcVS+x/2odPTklgiahDpU
a9f8+reLL5s+c2vKzX6nSWjOG4d3Nu0x3T0ExAckbpe67s4IyyltAZ8wXWPSeSyfpglNkGt853LH
DWbNbnjcoROy4B6sqsBqPCQ910eTYHtWOTszieLVapR57mliWZyywIShykb2IosG/mdCGaqTFXcX
wT6xXwj3gi5T9zDfZAuE4lrfTrkkGt2MOywhHM0rfUs7xGVOHX/0LhmI8Hyiwo2L83LRy/58rVeP
SjAXP8xMsPgB6HGzofcOGVkarMUG0sSzOx30xorRUBeTRAW5HZp7FJNyBSQTsftzsa8Xr9ZIYr1J
b2dDTps1TycHJ4/Zhw62hEiMGVzKPJ+bItZr7YO563bwgyyBeqBqmfOUY9sOjTxRjj/FWAY5geAa
ZGsUipxujrWx9W9Nnopb8ROcfTEMyvrBVmYmm4DqO6m6BEC/jbb+MIGJHiO0rBtSa7C8t3NYKWUW
UzvcjIitlc7AXHPdrBwTMqOIpVUCF7lhAHfsnjwPupt1ug0LMrwi5Bwf8+VEw2nXZAqo9EWxdUiT
pTKtCqiYBzzBiHeZERK3K6oLS1atppHzQy3A1skVt0RPxr4IpkRJXbY6VsKAKDRdRfcH3eJVpPH4
IMEbw8FJFuQgVW4X2MQKTx7AVs5wpZMefNyvaTfdAwCvIGggFKZaTjkcaEf80wnB+R+iBTXzdYp0
VslMsxg3250V9adpiFvhoXdb25cFRmVSsztcjcYe8B5tA1yqrA+TsEUqwofSSIzrbksak2jm0U8x
JG3fxONoF6cvtPeIpI380iIOA6DiGFsVHvjCmmYs1bZ+MW+WTKoiKMD6FJxcKixg0QdN9ypJg1q9
0ponZn0E2oHIUb2DdIEubiHRKl41Xy6vpflp7+GNWFJln1d9f20Qp/IJBRGcoWn/t+NVLSpcKuXl
MEOHc+1Xwjf0zHf0fYTwI3Twxbwb1/1vWMDSP9CXVz+PexvH1PpcOECsRBSLRLbq/gKzBAdKpH/N
ktOS0WLPWa1jr4jGTA9PVtoMyisr9hZZVJK2lQPUfl0f+NlyQGesGwdbLzGTybbtOntJeajxfqgb
Cr6cDGnO94Y6AMPoWlSZHG+7XbSsmFfKSIRzC2rN3e9ABUt3h+E09e8N6sy9+g5+HMU0+lahvcgF
o5D0iDupqt4ecb9JvekKJ0xKmLJ+vtaNg7F2HCeW+yFHG3/GVRFdxTvhqqKPQ6j65x3W9gR98vqd
1Avl6dj562dW/D/cW44rcn4HYQkUdAKTvEqHoOYsJXE2Quz14PRJV6WVHwcVpoaZSPQR8HO0884j
2wXy7RX/aDBHGn2VBrgCe7CtZT5ythRv51DeuQmscjJ+QWtwG/LTpgPYwynRySo0t9SbCQ8o8Nom
C7gua0YPPkQQ+5pi6SojQIF+I2jLk/oMNqunw3FsOdfauUEg5fjG0SO84NWedHXpik188JzT4VII
A6LUOFt/1D3J7e161u5iwZrCeuzaFHdaT94zAujta9fwenNaSJbq086plzm/xXCnv/UW7aklKY45
clMQc05hM2eDlLEo3TCmMvnaquUZ7/Ln4jaRyUAPKvBzsZbzEbCiGy6tuSr8+BcUzjF3lHf9tDIz
ccQ49Wt4A45Xwd02CGnEbVVwqSVfBi6HvmYKRyYq6mZAtcCgh/WyMXMoAt6x9LwOnR8Qiq9fKtz8
c4z0w4wzSh/kdXFp2vYJFlM/Ya6MrRqO7FiRlbor6veIEORCKRD83TeDPIgS98aDsvvhhgSd40iR
/cuCoUsnhfWr3xzWlO4LJPVwlEg+JzTbbRgp5JUjYcKBDhTrKjHNeBuTzvpjWyujdrJ7mQa7JaXP
VAaAbYlgbaqilI44woxH+zQMXng4Ys7y2iXbiEqSnvD1IogoF9ZDwiHgQIKNnyQnj5shvkvfuyH8
Xtoz5cnd0u58IlOoQrFVAroCsUilGr0Y6WYFs9Yp7bvEQc5m7Xtd13foUzC7P721TOwp+63ZoV5u
w/zwRD/CjHC7WdxFZqOZFDTwofdXhrGczyfwlVtBfr8ruilyowX2PI3ynBzraa6SvCUCAMAu5qlI
//oquA+9LUr1sM1cQ6aCE6XFfoxsQriZd9rYlhswloFEzMh1MPCWFwvmRhXJwpNtbJHGuLR6gXcm
uSUOn0dvQjVt1Gg3LD4eKFJPYN5vyuoUfZRiskRAtgNstzZYiMvjVwo9uqn3bmRPJ+wE0VEeVd5C
l/kKWXHwJch+BzNk6q/CWl18k03ZgDGy6ujwvXJHuIJ5WjpsQgLPmhGfeIoU5EHF283pJPA5rhqx
DpQx6Xi6L5Wrg9ywayCDLCjPh8uzJk5DDbn14zOq0EhLaR8dgcqoiIgi+Vebl+3zrnA7aHfZghpA
FlnGnvt+das4+ueIvzLNoKn3LpgVteSTqHSYiilBNWWdi4gE7/Mo+joExiLlpQvgp1ei1h9jKGB/
DSDqgSvfuofc934iLhUVDO40vaxOF+agulH7wltIyvPJhyLjiQlq3k8FlZO5mATGnqAAdFk1CmGT
oD8iVZ7Q4GTHTPaXVYZGheNVtDpdsbGDMpqtPunXp1gHvTIwv9zSDapNDdz10FKRIZZdNv4HCUyc
/WttNLDwJD73QPI/1EhpFab4Hr0YrURZJ+op802YNCDevzMj9SK/0QQyXF9ZBl9MJ50jm6PAOaPw
nd2WmH933tgPq+W3BP++ZiYT34VKd6AQGsR8ZOoY2kKTifopndNVbH3TY4hsQE4NkesxlZMw0Xoe
0dfdb3+l2Y24TxVwmxiFCM6x3oExuBPX44qT0DSkasmzzukd5NqFLJaw6HRy0MXaq7SuO0smRsuE
dK2Ht1NeCPPhwNG84L4FD7WPzz49UQiiTJNmpkLv4dthudYHZTbEtn/hnikFfPhX/9o46VXzMCa5
pVKU0iMvrcq2v5nMI6Pn1/YdTLYoDyYS6SdIudZ2S6xyNCM1br+SVQHtewIW4qvvESkT3Y1ESBmt
HL3kqBwZN3Tj4WgPexynzENuSLW2XlB59SDYy6Ccw1rt5JwNQDnEPqZ4H/JjRO2RSg1C8OZAwW1+
lJrtbuJm8rzDCxYoiK4mPDRTs88QbcJNm6lbZ1xmdBYKmePgmajnHYzd4qaxOnnvU5VVZEGGCIgS
Jizcx8t5L+7pMmtd6P/37GZFQSScPAyQEFmXaRG94ehO0CGGWQZD+oAQWT94hYenK8y9bn1zXR3W
hP0gDSXYh0ZL7K1v+eYFjaQNNzX2mbPwByZYm6waZNNagg2/WlWy13g7UQ0jcRG+At1hPmzm9JVx
rSTQKVEl8sEFwqL9ALBcX2lDOVbTupxIoAlA2dLz7Vx+d8b9CQ/Ace6c8dn2wr2YFGOwYt5r8nao
JKv3UdF3fJBvsZF9nP3WQh8cEqTo6CNZH1mZoNgjr1cNO/bKJtesBHfxH5tBj3G5e1HwS6pBAjdE
RsYplXDy49C/rxVMihramlMz37IXqZHnOZKNoZUI2gujjTGjzsxANlcGQjfM5wjgmTZMBJ0i4KLm
pUr8D3gMAHCTiMGi86O56ejih8UO97h6oEBoZGQ9rN5zzVBAs4ZaU8H0nT48NWA6X2af8Bb+l2FE
goPHFNdgLSaLwdgJtcjSNzSIgb2v2/hN8Cj8gKRzCFsfV1YMv0K9aMQUrUqOve+OFp0T227EwWPd
ZJEB03m1Q3EdUUZ7DIQIOa2T7fRJCHAVHyFz7DHPeAsfsNL1QfrQTBLP/iKvst4En78cukspnLOt
NOHTx1IwxaNPBzMWI4i/k2jfkAu2LKYzUPwhb+jMbJe2GuqzNjZaf6NRaCarvXSZeXxk5sKijC/C
dDRy9wSA1PVANsJUvDx2kgxJ54mCsHwZ7xMYM1lQjrpknC67ht1AG+TGJrrlnCDQ5mukz7wLwoKi
EdbHk63PqgtTplMBcsOF2TOrB/wR8gObVYEOJPFJMuI40ft7XeZ9BCAxTeTKfPL+tGop4SwVdrv0
pvdlvbA44m5hJBj1b3wjPaGGv87kAg2tJ2BKodDwujizPTOnERkbn3BAUNp9axj4DYPeSvAZxEWi
WrpXCELIzHONnjygQFFzyOd1XyhDTlQli29oW0J2hpTid06phR/ckW54F2rqesgBuh4/BDM6MeGH
Wo8d5aRe6ZuTTCjrTY79hjhIaY+R0j5x8DZ7WBC3JNUllVbO3mkpWXWui1WigqBIoLW3k90TpmU1
SdWDUXtKyQjQsmiAC9/6c+Mc3meR+gs9tV6iIiqgx6eXx5kYC6IBosk/T2iLJHIXacB85OdJyYWp
xNpJ78mWiRxcPrT8i1gaYMrjECWyOF7mvHH+oxo0IqFBYtgIN2deo4F9SnhHFBY01TaMziDI8Swu
UUFVk9UEjOkCIc+FukuWruRfLSBnHi/AIg0SsXbNi1qhNU/xJGDtI/TQtjbolqgoFSIH5dxi//ZW
Kz7tFpi9GpXLtPS1tSaeX5vPMhlZh1K4gW+dJ5Z+FBu3ByywuWwHMzKGSM62yMsTVq+vf8uwVWiC
RORT8HtYmXYEo9TRhKGPvsi7KVwcDAb84RfZEJ7T2j1sn83ys2x9LJCOEFO05BoQgAxZV2UEgtp4
Tp57mkZctRFf3+h4g1vk5gpGxu03GtAx4LES4aKCqYgrLEXf3UfmYm4UFgKzkn267M3wVwLHaomI
l6lB4xvUzvOlOo+abUhWAFeAWwB33euQG6ImXed9G8sCEPe5F9WUULc1E0ERwudwA0j6flK99YX9
+MfeIObt5qzLdyL2u8S6kuZ0asewTeAx+73HLDI3YsfAtHBRa1Q+vkKRCN9jYGYmhB+gahmrxL6o
v7sDmBRLXMrRzC1VK0TcFjeXQQZg5bt9rq61IVzLkvAVb9uo5rF2DGP3oxSinR1Nssg6QMZ7jchi
Wnv0s8dcVhDj6XIzMMtSJ+HFQmlufEgAA2vhcXb6Hw2wLSx5ni6/PzJG0FBm6d6rJTWnLzw1BjX5
ZXR9lgitlwvs6krYxy/RoqayLVRqMxVCJrUykR4adPpw5cw+c4TNDSw5c6IJncY+8YlmopYdZD21
NJcUpwlNeR7FLttDBSGP4TdAYr7SGnaVPPBsJaMdlxEFwRtGTWCAMqohkJVP6ZQiz73ROpB9zBrY
fI80K7KH+kiVVfwKZvyYyS+8/pyCJKg1HgEBBYFpe3rQnUs1y+rdSny+5C/UEDe0CanaMS2ko4/K
uYzUTMOF2/GjlSyE0vm2iJBUDaoc8gEkElOR7cAR2NuB0W5r7lb1kYRCBzqZZjMPXmbMS4u6YDWu
/6VwwlWSK44gMw4WZb34PSNB5bQtKwBWnLAdLgtWxamzWYOUjaOnQyVTzAy1iSsoJPmj/0x6dkML
CQnVz6feYLJlbFuumm/ebPJKqZbqe9Y5QfnE5uyoYddy4ydN7ATbqqNs/rpjrJ5LiJDm/PpA6mLw
ZpW0RsNnjHbjiKb+l/d+feE9yh+q+2TkyWrISexOK05jYaNJwlxSqVm6F4Sa6cuD5UutsayRHviw
GD1uqyLv7KEGZdoOAL6+OZ+jruboiEV+YGePoYNVQGV2ys3KtQ8g95sCC+BNPwN0h/8nnseN2vJ/
XF6PCQhJe70ixb66smNrwk66tFY4mQmrRw15zzhZmrqJxGZj/SQWMK49D5YjcGlKEgQ0u84856aO
yzMFyBt+5FKQYdbeeZVtSZBRt1s81HRq66YTwEVuaumq+MXcAiV6O/vCZ/XRczn9ZXsHoe0OVQie
Iu+RWvGamtsN3QkxsHuYUEyfOCNBWSEa6zyc4NAFeB/iGIU+NIuezL8BxeQf9zyUPPjviFn1iM5o
cicZ6ViCxYgoPcaNyz5AmEvUWe0gu9GPzmGbeLMeBAGNORbj4OMpGdiMvQrlWDesUhPB5SX5e7uk
sE6phPrS2Fmt8lb/uOM4rzRhqH3oPiDMRIQTnMj4pbjnqTlhqe+pNej2EIIGwHMWWZCAhUkL1axW
ouCDRhZfhBdrmyrzSMVIqT7MuVn/ZLyFnCuERsuDkIzixDNQQStL8/FnhF3AmwNhlampAYP1VvDB
cPMZf6qx7mm6aRUMEPNR/AKSk8hSnoPSi7bts8MzTN4oiX408+Lego9tbSF6V7ZZNP+iECFVTeDm
cmtdUtuhOdp2mg/r05FwcQ6VGtZ+6vC8LGpXXK5MtHgD/Uc3RDjsc4LbNZK+GQe5i+OPf54Rb+2g
pp4gNe9n8ny2HsdUalvkz4p6kR+AYHKJsvKe5ODNTL9yJG7qkUr/2zoGzjg0fsEiEZ7z2C13xlu3
Y91UpeQbkaG2Sysfld/YXJDDiJSmA5lA9rysACiTM9Q+J1sfaSioq4s7c+BmwAauVMkJp0CVIHRU
jQSu3QcY41ygMhs50JgGJv+74KY88qxGyQ0JV6gU7VD7zw5VPuDHzGls7kGOZ7j62kMH6kK7grx+
DxGkUpyy3rqw6OmKJ3sqJMZLK7SEvkya5geBtN2Claj8fLpJiJ9US0+rm6IQGBPej7zg1317R9rw
WUoEscINHsCEy9YzagzQ5pzR0TZYPBx+Y8Zd+jtiWECVZ3s8dkgp0v1zTzbMD67Kk2IyWe7vwiRZ
bMyOK/nTdsjLxeWN8p6DXtbCS5SpTBcc0Marpde0PiQRRtGvp6HoGyZZ98smmMxsZqQweXY+GNkK
91KwPvcZW0vsM8tA6fe16tvWUYQNsp4wYExXfiNnSY7sZMhp39/vmcDY8fui0ANWIqCVdko7dWcp
P5oN9Hd9ifNYAUZL1Gn96RsnDyd1nz9zxCkSSTw2vA5/ByTIiLGTKpgeL1h5ketLHaCpOeUCmwW8
frjwJvaTWBoTvPeGHab8evQuQ0i6E0Pq0iU48e0DCv41b6dkwzhMqvT6PNRgJ7ZZZDInMJ08pyZP
+tb4qWmrlM8dWwZD+Z2NLyHgwPJ+vu6A0xuXvJZ32VBMTBw3ez22x+tS+M9ocqRAp0MooEiNodsQ
k3kDStU8kLSNmBw2CDfvIV8Bk1Xb6rr0Gm0CmkIfRJ73FuupDIjZ4lfgFj0iIFTsYF3B+u3BzW48
QZ3YYZo8W3mG2Ku+lJwsWdeUq0a+8WaLlmbNbtIuiBW2sFRo3RXvVV2HjgZehbG4p14rhvLulj8U
oyNyD43UzSbyPwdnW1BEEZt6jQdto7aTnbH7ACBHnE+hijxaqizN2oLHsKzlQ6PFQKy2s1MnCLIq
dydE6jrzq05DyzkAbYljcP0Ke17RySrnp12uoG8gkoF8Z56xbiWvN+bXIMGgQD/o0dWcY85r73Kv
rN655ePzwwmWsGFqI4Prm3iFh2prlQ29hkrKI3SwNj2RkF+Kwbowqb4LspJfVZAVGv9lBnh5pvk/
cBMX9fHkhsBcUHgnsEvbHHF02KJHQzpz9Noux6txNeS14+KnFBbs4hMH0Q6ftrD+pblOql65rvyG
jGmjrxDI2SrvIwwbQpkmc4WEe+PJu9rtt6u6zmThsitzMTC27tHOKmnn28BGQYAwAweOPJdRBYIn
C7OEq88Vz4YXbLkUGBUoUlaQoisdJxt0+zNxOXTT+rhPmhNASvJrE3++NrmXpV5hKmB4+BqLBERp
VcVx3oY30XDBTJxlbk0WBBjTeNcNUkTQoY7a7s5qJP5PKFtQIAfz/nTlIWeQKdVso2U9XcNAcpkQ
0MJ1ff//DmyhbMlCD1d6pjydclx42sdxAH6m+p4EdEm7OdgY9jFp325mueLWvaTEtGmOkWwKvaX6
TC/sMwzeh2TuZcG3UeKepUSjiL4cEYBCbFqy7EbdGNeeLfiR7lXudmrIZEVv/l0LUn32gNJOauCx
FWeYXungdspEGWqGDX2FS0bc8HvDL+lpbZH7FKtCaTH46CW5sI4dvbl+SkKRol3szP/i9o09KHvG
ybA4deZSp6SAC0EBORN7p70hEZokzsq0GOwdm+ZJqPujPX5b6WmxDxhIhlNpBoFIPAGtDe4i3PGP
jSYTcXyg9i2I3gV6m+jo13Uk5cjn0FYXQOPsJt2KOXuWsUFACc3GUyeNVGnY8jJdKbv+B3b0pC4Z
H2lRIc/cdOTaDI0Vy5llj1GZZ/pxTr3wQblja5SDgsvMIpeCOHFa59hKHZ7wvReEFseuvzFCrS2E
dw7J9fD9nQn1vvVIN81/tqcEpi8WEz++dCMykpLpHNpnUeUogFCVVbPzNHXIC0zM2qsyEdfP9vPf
mzcrSSvM8XCo0I73iwEapIAZWX7tTu3ej7u3kHtk5WARR8ByT3IYp63MF9N9n4er19aO5AQMXPHN
hIlDRhsINZM3J4dLpAuLhhK88zTFx1HbQT4bWJRHBAs0iKyrLdCR1iL3bnJIeQFm6ApNddJWBBuS
GyMsB+gA4KNsZQHe+RkUKKSVAT3iM9aqjkgw1vD+jxvCTJ68fK82KuVBbyFGe6HXl1yMI/+f54qy
7VOKqHzECjryyx0C9rHaPcoMuOQqERot5i+LNduUYNrrmBqewhFuKolClZIORJ1AnB5tJOKse3zj
xP4xDV+BkwW5qahkw18bb4q/sxT89FUHuSsApzFcV8uj8NwDWGJhiDHVlIanqiZDo4mhExe7Ibi5
iAJ8fZ4fkcme6+MCkalxAYfesCUoM0peLhzXrtHP/D3IorNQZHwcRold6cI6NCwob8qx6CcZMIpu
wmwipe1ackCJ3JEl+gDIxfxbdPOMSFD1S1mF7qPNMC/p06N17jRI57WKl0pTZc7e6l11mxp+nb9f
fnXczxw+oQBUV7LSFWhCZb0gMHRKxTA7yOEVgQTcF4IXJQH9j6t2OmCLHpXGaBQ4GxFxWHK4T9xw
v6sBGN2XkN/uPCNc1heTC0YQr7YY3hfAiW2y6lB62pnd93gxt8RR7Skti39f09QCcL1HmAUfXAD8
6a+QStYulh13FgBHAxFaSNnujymypC5JfPXEFTiyc1oo+eLpnMGS89dg7tEqvRSq1HtNL0f2Td2S
XmWgqzrSf1OXeaPsslY9AkGS7RLoMVtlFJc6byf6+/NaoVN6W03wuh4QpWNUlOc9fa9S7CjEGxJ1
axmucBQIaksLij4eprLXjSwimHJms+fY+7HtUfeW4c9b/318+VANitQTJVuc/5oW9aNKRGq0rVuX
50xKe7R9ytlIEUw+WXg99CI9UQ+GFh/rvT8dv1szJ6r5sZECRoRSfeVqSFuZf21HPNPyIKONjQ6k
WoH3TAgIiYhqj0vpqdGqD6qslGiaWOC/BKHxpzwDhpXM+hWwjZHvDnWqVKC2Y2G+jKXn8IGMTnBZ
k07WWn6PAWjhXCOWdMSSo6D9uh4J9pRUpnuSW5wqU89gbu2tau7Tpu/uc1wpiFe6glTRUG0aKFCM
zXNpO4+0xSBx8DTOHCahPPfxfB5hHzpU4bqi/IH1F1jWiI4cZQP8vz6PMHjLyUcsE93H178XO0DU
ZNdokk/Kmj5epB79TSFoLHchEq51RZqUOcuFmuEOnujh63qRu0cBJ3M1g9xaYhUlSFW6NugIhja1
CAqD75a6ivsW7o/yBMYhXGy5kAA5AH0g1lriMiJBi3PAPFfUpCKsvyN2OmzYoLsLRpbBDnIHpoKh
1PP1Dkn6dZK+6OqRraX3QlJcNJMJuVA88UldHvAvvqh0Y/diypEs9Jk5aYR7ZneFXvuWd7NX1/S7
jlax92zh2FubM33mCO5HR9banU2ecQ/EOdPfGG+sDmIKvDInt2zRw9nPkuJcq2JCOFyjG6sa5IHO
flFk21gcg8b37gowIn2cXfsZAxQExdYi+XsvCY1nKwBn1ufg/enBPfgetfy3A08PIcKyWouKCx6L
wLRtdYJM+sQ4q9Psu1TQSTIUiQmh6Ere1Swd5il52zZymydLZ+2q4HomWkJLTpALuOCgumq/KxyV
qkr7dexF/xpMJ54QazTxwsaIOI2fhkfMO4c+Oeb/+7gp0rWs7XrwhNed7ISMH12Qxcq1LdfjXCME
1Ve+GtBOS/xGw3doXlbrFWQSO3OSAMLqCIyENPsywi5ory5ri+eRqXcdy75Yir2p1kq5NnA00EyO
mX9eF6Fpp/OKC9rIzMm3V+5ft9PGTJENPGLjgMeD8ebHKgKnHxcq0zBkcWgNqwfCDn5zoBYr5BoV
N6ea/mSX2ZY5aD4VhFNv6GMOOceNoSjjiHFpQqam0YsKK9Pov/livyHu14qKwL4yCm0uqfHwbZ7Q
jI25DqWuwXXkSAdEI19z38wLInCm33XZPo6r76DaRz0MZCFVaRg2tNPmjg/NA1mVsn80wloSStvG
S9ZPE40RoMI0WLyS730fyoRv8jkLmc7311/rleE9tKSeFdcY5u5d0gLUrQDG+qmVufeLyRYgyl4j
PzY8itNKV/lHivTAIwi4e4w2DCPOImDBNb66ScZKWDBkzBInJCzEELWQ33imgz4AO7jAsm7G2SF5
WpfthYv3j++XfCWBzwyl3xvWHr5dAwQ4t9ghSn4pWRPQnzH7KvHCQ3XJvwCTXSg9xVsHMF6oW3+j
li5yj70lMulA8SomOLPl5E6LISb1X27aT95dgNrWHaZdmYWtsJR4bOA+xse9W8dmvpSZ86Cu+HYT
0HmZuYiDOzu+ojpR2VeXab/P3Hn028KfbtQGQqyfeR6cDPLe4l1o+v5gpj2PHiXB7wR3fKG+zvF4
g687DoGcrFFLq7HL+eBzH2ISXtdVfyinrOpjGE+973diKqcxCbPsxhtm9IcbZNTEd0kjYAVwU/h8
WWBSdykPdkLEY0WDSNI+FgAmNY76id99kqExeNg1hnmMKnLtXR3BhH2cDglTaty5K175kC/d7sPM
PjYk8vUt0PnOf93++lIoNiErjVyNqw29n31Xd4NUv/DsHaA/b+jcgR6R6AUtqXwYJPgjjmSls08q
SJ+c3Kp2W56VQ+C9j7+WdXsn9/vlUdntdVU3KkWUhkZh5UtuRnffIuS+fdON/gIXRUqlN57JVz/D
y01EDwnjE81Ud/VfRuQ34sDhINId6h9THqf4dCGLxi4SYZxvK/bGbiTbNjCuGlkejjf0zdxbgZwp
tDOAMt4kQa+XrPoyzNDaEflDY7oLvlL/uG1pSo7qSwFCbGAgqrEspQCwHBZl52CYpY8CA6cVMECe
NLvZFG77d/8wQVRCB2WBYBkw1M07K84piw2oHLogkciJiq8KOhYEOmrb/8ub0F4DGqbIC/NGfvm5
faZs46peANTjJdY07QwVvF0q0EQmReTL2NZ8AiFe6722K9Up5n+kcFEsjokDyXMn9F169rDCs7uZ
FeYPtADzxRDU2jV9A8SZGIGLY/yiwbYoC/UXLck6JUV9fYk8+TGZ5n9NAZSEawWWfH08tqS9lvFO
f3YuN9Cjsqjkmtw9EU8s1ztTR4kaSLZAyqWegCxdYdTv5gRFyIDGbkyeEFS8SkJjrZeh3SaWe4Mc
iicL5XAANgDBbs0UwytrMOyGDc5qRhX47iVNp9GI478KRyC++ZPRcgBlGmgYs0/CTkzMQ6CUUp/R
7PwkkbCh19ct6zV6FRavG+kgAM7i7X+VNOXopnd7CaTmD86WlPjVKn+uDs7S4QZ96SvGYMlqtdvH
1XzWyQEigkPXI7BToBygfyR5+BNf/7DuQ2nwlMsnWtMJBKYbUKKjKRhVuInAGPOZ0CpHmBbs+2PM
kpfa/HYI/NBj4K0hkn5lStxEuWy/1mSUeLJj1COGtlWNwtkrCTcbNQq0/nDTyx24M7Xuh1nWSJy7
htEhXkfqT+FS58RLaIKckwZhEZzUKvLOtS9OiSsJqE5TCIS7mJdI4vkM7T4r2nJKlCS1qCbaV6HL
1+Hqs/WEEhP6ZOUpxxPDwXN6ibUVEdBVLlC729pqPdATGBCwDQAqa16Kvv5p+KvApN35ZAQJZ6Qn
iJWHrGX0ZyGpfxxNyhXJaaYfS5GhZteBCZtrl3h1atosoEpA7d+/wJbHYdUWRXKLiFjVFCqZQ0iq
Oy/J/fLURdVtk7/3nIw6e/77TqXggH28uDy1LJZ/7IveaGQi9Tx8eOL1RPdtsEPKjezCX2E1FZDc
ZTjpPjKWN0CzdspuApr+r0UWB1PcCwtzs/xzw1ntqDRaLeqoIkjSl7sGdxLHjkZSZqdEnuP7ey4B
tZS1RHYJlrxS8CxSQaHH46C06UTZlKB2a9P0djfcYj4MPx9VEUb0YvHVVc7XZ9ivDrLK3zZ7CucU
sUzeExTDVkeIajLIlrfZIsxGYwsZvG+nWDhrfRjo/izD0xkX7z/FFU3NRXEWazwD+lWF4Y346SzU
e+jMq+ehuT/rB8lSuhUzEutL2uv8IjQZOtcQm/J1i1rYqaxsfMhxB07edhvrGcLEPBgnRmSwZRus
IoQytcPKAcOHf0C4jIVMm3rkqJdfccGSj9ivHs1U+Jnv4V/3eQ5zGH/NGXRIil8W2EVTILdoWltu
jHW1Ktft2LJ65ak1Ma5iZRg3VIlITeLn1eQCANj95bZu0v9bRUPuw/4G65YdAQRXw7HqbNU8oPDj
ZZIhKT8ooWvDhl51Qo/zqX8LD0Dqw0Swlr8Fs1QejTGLMLltrch1R8Ud8Ou4fI5eZfdo7YAoc3/F
9Bmt8xJuxYZqiKRSbxu3mTpxcfyrEgmaQ1LRRKFLjVa/qi9EKAZNMjS4c6PEvDk5Lgn35cxGUCGL
BMoybdC6bktJhH6iGB13o20QL0mWXZf8We2UWvrTi0VCYM6KeGcOonO3PwsT9OR0VMHOfyojG6oN
RydnekOkmhJKQKmEO+FwGZ91QJWmZo+Ns6eVpkS4P1qudh0yCBlUZ7l27QGWloNLaQvKoEccsxBf
wlKoOVeAU1Db29odFEIfDrETcSipG4GJi86r7oUy8jGEpqrUkTGzCswxR517D7NarZlpcwuZ+QZZ
Irbq1pE+HGdXr20kimSVwr1iT9UvENfk/LvwZGMnjHNpFZlixSqelNH54xmS42NbZ8D1d0iWgIxo
evm0wg+bQx58rzDI9pqiGluHTgAgdIl0eeXDmVL/zbSJUVEvXmgB50xcfhY9TO30w3UMjDi1wRN9
0Jb7RIXTcSpGTM4kSBaBPnEGds6DLyQEBP2ivQI/0pnnO62bTuDXhllrqokRNfIaOqZdKo7nAAns
L9bBo3llF22JVydjwcH+UnIhEuY0RubUjUH9Uvr+szwiwz1n3ybgpss8bdfnGaDxyxBySMJlfZSr
KAQ66TeeryuV6gaiJs3WRKdDi7TAw2KEte0Bxki6ESV7vJp63RGaWgEYhz2sdG2uQ3rXiAfgYtGr
x7XAucrbW1TQbp/nZnIlJkx5dRY3gkeJL3kC2A4I92pFOGGijs30l0OXbrDsV6lqO1Y6twALKXp8
1KJrsciRaL9haEtMgc5n7JvOHncx5YFYkhXRyTZePSa5hg6K9Qxkxs+sBTB2DTV9z6Disx9X3Wyf
dODEgHKvNm9LejZqo/v0osGWGcagtx1I3DMUX70RVdrPZUnM+8jYcybrD3oQch1U9RhGsXEBgygT
DTkrhyAaStN0BjaPjPjNcFLRyQ0rd164j+SYP9pokvEO9HCc8L3T8QiMt1VqZ18a61duxUAM8y1P
c80uSAKSg5P3fmN70swo7OcN9jVt3QPfl3v9F6iDD137Nv3VI1qbwK/PVJdmkXJDsULXcFfHCSiV
7S18uxgfwJFyJimpxmLAmeWeCHMq5iKnu/FmD3ZTJMJtE5a7VhAfs1KBTTw5qMJNhca04t95iEf4
lmfFADahyT/CsjTfPZLQCwGQA4OewiOT3PdbouxE4vzeoQlHl6RHqbZkVJmhSr12u+jrEN+/km5u
Eu6RbVOOhcQ32Yp6v9TBz5GwzAbuoLfPM/vUIf/pRh6+TqdltACApxSJIaHO7oVjBTjtex5RMElv
JSVzJIq0aC9ylFGBH1KbgDc0JpzEeiqdHi2g8KDzycoYWqrsiXSDEhCLfbcA9ZXA1CIEF7xg/1xW
Tdr3WY8IRQUrgjAITwh+DgdeAADJ3vbYvAjaCEZI9zvA8dSWyQ3tA0a0rNAUnulHYivVND3xH7pQ
5KGzlObZX4ArDIZG1mPYN+SDNOUA/CR9WjQJLBEyiFkSpfBsXE/X6kYU+ngVFno+hQbamQLtMlrJ
nlVgc1bNfv9WQdAcbxKoooTPpwHJ3MItL0saNtvi8w14Pix2y8ZHMA3k5WxFooJpDjhwV7Rt67ah
ICTbzyD/BbA7/XNDyScDdOu0UVp/SGacazc9IFvaD6txW95xkjDknR+27BuWMUw/G9JiUx7og0fX
OrDEyiZmvGKnaejXDJAQYSVobY5cjPFFfufulUbLHyV9qHcl/6vV3Z0QZUAK6X3Bs0zKeiraAdxl
18jW1T713NqyUNLsZd4y7fPoll/PYu44HKf/hCzJ1HsDvTgtB5kJRNfIvTXusEu6sdmPF4F4BVXz
Y5Hi2Iae2tovVPsGk7O13euS+N3bZa4oXwSK+FgRuu3E0l45HflF6oBQVnwa1wxNMSypiRs5s+iw
F6OmCINrJCPck48fcbkUeSkmOe1/2pTIJW1F2l3xspdVnZZr9M/zif82mUuHVO6yDXp2st11j6Jl
wqCh7yo+e2kkPB5FsnoF97Ysjr4TEcJcL78x1VjXcZS7dun14a2lzwszU3ayB+pq/KS84ZNwxx8m
D9/PBIEq6wmgPpRhYmmP6LKS5DQkOX2DOh3u7gKlbv3ftSsVi0joqzh1guaTHDnI1fxCOB9TmnRX
AKMDC+qEURvt+LTqRi7reSN5/atbdocd9RDhQrGFuCBAuxLr496zNef5IhjbGOneTyPhJEg0oosm
n8aJsF3sQLnNU2xTZwRBEfH3pyG/BHPaQWZe3VnEBudfa6KHjOAxuDJdLULc1TXoVAUj4I7R16FN
DmUyq/0d13YWeaCdivHhrzZCfzpaLedoBd77b16JX3s0Hlj1siA1qpZoKNIlbZ+FkxJ81jVu1diY
CPER8zRIiKf5cJMeP/5cSLAMQfC5B/yTwan821KVHHPHYLq8BPUc5shqllrhnsvDUIbo1esVlSBv
SickISwPEk7GxC5ZVuQAMDvxEjV2pnsWWPLOfhVMR3dJ1BPmhhe5jCw4qIfgol5XfZhYiQp2pgIg
1SDqLbGN+g8vozwOG3TVeGk+3+NXXIJNPC4AnQblhZscT4hFTZ4eC55zJsAlfSE7hAG1MoTpSlZI
7+O60kVYtc213NMJfuDTa5ZkbKy+7wMgBv1QAsv6OcWP7JP3UhVbSHT6eh7TklGGOlj1BbT2oBjJ
VbSU61awYMirNvJqrsq5zSSSiovXWLt4xz29UIBcqgT8ktUPzX3FZ22moipnpDPJhceAo4JNVUE5
5ApTt/apbVcgl+Dc+fI34mdapaV5OI0Dgqa8XSfJ4MbocS9qX7nzUZxUmUV6yKohWiXIqZ9gOx35
IHRffyJ+U38mXkp5zkURTAULXRvz/AhTGmMonQO/5hMnkrTuUVd0E53ogL69j1+YA66MBafLn6/H
n8M1qPE6RpkdXWgt0UKvKuJVKYTdLN3QDtz+kcyHyGzx+Qa71RmdTblOU0DvAszlwxgjrsB7D/ll
sJ48bagXNXTmIdl9YG9YLC3J4F6vKYAjA1nqqIrPMNmfxJ8oGtkT9jQnpN4f0jJBYZhiXMqi/PIj
JBKWwyHVADfTu1JDkF01oX1mejCy3yqefVuun5tqLH4DuRHxJY8cq0mS9Fw5Zt7OJb7YN22V4mAM
pVgIj3ZujYTjBL0QgxYER+ct2GXi8K56NJ75sxMDlrX3T+HSslHC9KcSpcEesvY/oqGLw6e01/WH
SiyhHCs66xbEZHtz2IMPUlHWhZc5ozp8BQUPbPxFYJOvBqAlYS5OUTfUIE67pedrMRrw4kzAr7vE
eUPJhe/hR39Xzbfs+X2P0NMLLXDPaVkC8KFT+275G2RqMI0pHkyN69jTAWW7cn9ttPx/6ZB23CO/
TdRhsF3GmvR2IzbUijxuCAvKn6r+QP0H0+JFGLOWygDYyRlH4RXjrOl2/MrNN/UnWsfIxrxUj0UN
5UVLCXnVPTRDykkMOU6viSea2kY41pWa5RprYkOLp/lIxzc+af8T17YEGm3WZNo6mii20baUvFSW
TBBJA7CqR12WavdWYddWTKKgKjrdauM2zKWMGQFTpxX0qGHrLcT/q/BXM+Ec5qQWyFIxyg69Ysu4
Xn59so1NKSFmEtt4JS5IuSeWP5MfKdLqpmRxc5ynrmY4+HVcjM+Jz1an5EU3xyD3qRMYMeS0WtP3
X4/hpW1JgklrBgokuO4b2xNjacwPlpvT/dVtWgYhKFGEVY9K/SFe7+LxRuJ6+9ZLNaMgXUgYVOBi
T7BRpoRlY2Wf64hHC+JV/sE3QdDNyPQEsmb9NM0eOv8tez0HpNYNKb8cwToUlUxnyoxBmQAmszNx
/gUFjUh8hS8BUg5YmwdoFXqySGeHWxXbKgHjNBA8lZBrtTZ/OAY+oKaTvEom8SBV0C4t1iU/ZwUw
uZxKiIvBKVhYojtIhdLOnjMQtJBTQrmd2cQBvPI3UwR4hvyq7G7qGZ/Mpusy3x0naeGCVRZ0Paks
9cP8Q+zrfurZ9iyqEoTApzOj+nGAJesZUEEw3UApFhYrq4o8cBQH4IJC4KUZGH4w6nOAMO1T3rmy
p/YpgLkEG8HLd1HiYXmqdCdZuUg5Zic2sW+8wnowcV1bK00lRmM5ilRv6OIs7+dyZR/oMcvglL6M
dKEATRI8uPQETJijE4VKAwzsYnJ/focqJLAjvbECQhqlOmgZOt6fu+avChF646bahkwFIqcCzWop
bqKcck2DRng2VQZwRdJVJ7K8EQbtf6Ouowt+H+/XIV8DThnv9GehZZM0es6NqQ7sgub3WiEdL7C3
T6p7PX49WoBqZrNoNzY69ZzCR5al5CmX3uHQsLNxceD+HgnpTT1dX5y2hooCKMbNo3R0CaD5mw93
OZH0QXj3MT1yJRY2Ney7I7aMuYJAcz5WpF3zyJZ+X5YoYuIv5/Hag12K/mru4z2W/jcvsVZz9WlP
bZqWzIHoumnTdBI041A096uHZDk7m3P9/wzhfaoqRMRJof6EusekXzZ9USwxJId9iB5sFDegbXM8
vfBRUO11lDs92aOdeGfO9j6SmRWKMNm9B5zBwU+c4dTQhx2z9Lu5g5+UYYbDiWhUm2d0EnGdYcKU
mXaKf2UEqIsf+9cgCpviAEYM/auvei4RwcCQ79KPIcINHa+Sj2e0BVnc/aZwrBdk7EltF1uo7eub
C5gLXpUK7HFNQX39elzxZr9PcCa90QXXorWSg4xT0cvvy0Jo0oV1DezmZrE6vkKF13Sv2TV18Db4
6PQT2VoDDLOU6dZMH/YY6ChW+5hwVjSAPhvYK8IwFdb15mSIH56nVgFOC4HQy13shy/xdh7HR3AB
/OUf9z4cdRkN6zc50X2t6VotrmdTlFRuqqXFxqrFo2sN57wxEe12TpLMwBTdLm1XXGxT1UIZXts9
OqUYAGFYlaw3suQA9TUiDIqShq4kJQMafUjnxxrkSYo94gRt4XSYJLn0j7AJBWWifh8DyIUxPchZ
iblQ52ra0Sfze3fEhJOU0B3Rm0edKUttflv2xMZB2obIWIxevED45LTgOfoXFPuGGrxkP7bji5rH
AnpmloAUKUgTYc3VF2mTv0RAXsLPb8cSBtcSqz46xBNvPbR7d/D5OUkMVRcT1HGeo7fDWm8OaR/x
5/Rl85Nz8RJAjPmdb0SoD0P9G33PeINzpJ+Ny6sJUuqatyVLE0BT85qR3ei2YH0M1EN4f7UT5PTS
N3P9C1KR0dgF0GIT6tKLOl8EmIXMxnHp9lWHUZ+KJCQyMsL3wmsJ/O+wxrtQ2phXOw4/kP2lX7x7
OXXtbVo0f2zwJxbOcj8q4aRQuLy/ybKfQo8uVcLm1TDst62fKYC+z5Du5RQJIniHPBUBMVnAwkwf
opSEs9iyrh0j/E/phm5rX5+o9Cklh6UYyTLeUr8RDCeYvMMRKqI5Y3tX9qrToEdS+VWAq29DXobP
MlF26Z09tgm/TkgikRMCfIDvkdNm3obHGYvRRPuwmIjKoWg0OioySp0E6tc/mFEPgiAGps9AUWzP
0BA1+F5CKbt5vP6lqFJWAv5X0ciuwn5F9JooKovDg7nteDtzabweGJqiOHi9rHJKY4n9wvbee2/E
s8un18m/2878MOCndSc8+Fk54YMCUDDAfpwggboze4raBRXuRak1esMPo++EZ9TN0gKdV6t8E/WH
jPmke1qP16/uhxyw/TlMylPB2nAZaFDkRtKK3PKmGcCKXy2ih1dW66MmXiNO2nmAQxj9ayjiRoMD
R1Euals86L9b4JyIfzA+zEO+BLaPBKqDiJ92XrHo0cKleDhWSL/oMGq69tXWkHRbSvjZscBEKy1R
XPR14MjHNXPCpdhM9eb1kNkx8kRhz/fWHiF7oJVViWoq5omzQSsgXbeHBKvHjta9X3k4fakzz2X4
4rMShvwgM5ms7KBIb+pDrpgpKwqgSDl2iRxsTiZAYO+yYEVCqhZXz+dUTmyWuRAPYt0KpyJSNZFE
DO0nu6ygizBf+tyGCaOtPrI9B+njjGnKEFn9IACmfX/UDMpT/0L+vI/NRNlHTm+5wKwkiVXoeiYn
vC8KedWHVP5/6AMUpiF3hlRHqIXiXvr9dPeYy9flaCAhsHgv+aXBUVitg5l4kQpbHb7OxVpsE0wG
xbNH4FKLcsbUF/utmhSk0E5UIN9t5AFIapB/NxR69i6bYZE6sMef+6wqzuMkd/L3THTgNT2EdTwr
Sh4P6WWfaMrlknIw/d/Ky0NozsDyVVOBy5bnxYse/H3E2rn+KXBPL+nNlZt1tgYcCOEFtL84Z8JE
Y6lDdRe2tOTf7SaKDYgkVC3LnEy+1dwu3MW4U3fgvASXoh7AJVlFRuAQpcMxjt65gPCnmjd6Gfg4
Z00effM2RYM4ljGPMh6Rin/toLcKJhzw3JhMJEwG7zxTuhABzqva2zmzY4tsNp7rOi2Ax39hGBAq
olzgkUpy5WxjQDXjwXDYzlv0miaKZgYpEy8SClX31Kb+Yzf8dKQeHsrDzprraS0Rz4G1oJVStaF/
8EnGJSLQtsv15TZygrmiNmihQeUh90FycfOo7/g3SsI6I43e5wgAy7sITze34LNhEzkRtdtaoHnT
zuT1zoYBHlGnrv1QIxH9+RIemadx3FRzi6MksrVSVm3gDh1vqi9JGBEHrzS9hGaNX4x18eNofuIo
ad/ViyNemBIezUsDbP1rw2CB1w5W30I4aw6CxnS8qFFAgEeNsHpb7Y6b4Bn3m+bEzgqWtqWcRMUA
Y0OqOlPkedl4T58DjtWmmLOl9+reCigmGZtSnQQt+I/dITKpJkaTBMFXkZV3yraEd/y8OzyrTcye
J6rAW5W73R62cpSBgsMTDHwSR4223QTz3rrXlvMnYLeEzar9DqsM/HIIAfRmbJVPCQtLk10M95mn
mM41MkhocqfQHGzchd76rJhBHX29C8G05oVDz0YjVE6kHER/yQFN3MH+tlwTmlU96nyIb5kiSTDZ
AqNhLNq5Crs8kiNcTfsOBN9rJDlgunGAGIe2Ut028fHbN1VACV9qgXuVuNSGuKEydeIMrzI2/dYO
t35bv/502w2j+OF9N0NoLpN/00/iZucB54BGJBCo9qfMJEIIkxGGWnLmJqnGI6DjzCIhx/xGbQun
lyIHjCXag6soqscRyyKBVx6J0RuBcXA2/sQe2COrSA0JTXQCjqj169O0yaHA99ESncCQfzP9CW8V
5sVa3ulj1qWe8oLu2cIMgSUg1CuKL13jcCQT9xhQCS/Xp19mq6zB6Mdjhnf3lByTmRRLKleYpEXG
OAEvikykUv4cTa3Eo6swJC9usSPB8uCjSf2nMC0Xawm54KlCPSt2HhqKf3BoCTtxLw26uL+e3bj1
YmvCjCGfIcz7QQ+xQWhiK6EUDO+z7qUPgvi6PsV7TML9KOLsqOnhbyUl9P9EvNqbfSS7FCbFkIHz
QgNcnUuuzQuy+dPUOD0kAvxJNmZxllbf+9WRw2X1hHGNbYdvCpNQ/S912/aM5FL6273wp9dZc+bI
JFAmLkmYx6cLDQ1z9oLF4mJDl0OLgNwTvjcmSdWb+Dn8PcGvz5YKLpGxZfpm7lxfwUUTlGT8LNNZ
UGZB+GsqfERVloU7enm/ghiLlD4Dg09PETRnomdggzTnRz0Yom5HRMEqaOQHFuXx9sGn8ILQNUo9
eTjZhj1dqkKJco4OZCof4xNP6W4m/yuZktEGJXXzgnBREnJQFywf7D0K5YWUVwUFv22JeN+zws+1
OVMQWWSpZJM9uCXAV3MK9BFayI4GqHjSYggK+NX5+OJ6Ep2/9o8ZnxpBPXHyrURjDRMGbEdhHNhe
F7yYbX7ZFvsZeL9GNTw8fI20UmNzjbkJ66J6hFZ+NTM7gZdNurTfOdxo32SVF9Y1Eq3rOOfIO/ox
AgbdlLPjFAoHUqC9BVs8tNaLrfsjBzKv/AVq2rtmNsBnKnm2DliKv+E/foxY0xY+Y1CuAGHrCH1I
tH11RcpQ920eQzjzBXes6CJrDCtVaucJxP62o+94PIDSg/uFdEqofPsKELllrY1ehTHwUx/dvJy3
oyJhQf/BkAxVuuG0fZgUg/zeazG7xWu1oXbPxvTptZIQUYS1IRomzS9dHwV5ESJCJoKvDKLUqrIR
RFGTdPBX6wXielCS6DhD9fvIR5Fzhe95XyMJnzmP7lGyvpws6xmS1ZHJZ2IFFAzMcNHvGE5gyXQM
no1nyyYdlamETufhjtv9WGrjc/AMlJtDuzOX/ka+GODyVEyYWvK8CJOUPOWbbPynWE4uPr2cEF3L
czttqXbkWR6y5OXXFO2/OQhMHCb84LtWRdOr9wqCYfwuUIo2cCgUSOJMnBkMalsMyngtxbQ7Ugu+
QGFkKtoTrrQhcvF/egJg8YHWKZPx1xzj6VOssTN/A2Xv31IaY6R/DtQiFN/y6C6c0O12VgD4Swlk
dxR0+Ho5S2V0Fm3YqnGbwvSM6hA89yhnYqjTPpP5v7aYO+90gr6PJFlnZzMh6Q/XEx+2uaNNP9vc
6wfgJWApW0mN9vqAptvWdLATHx9SSPpb1NuO800oW3eseEgKYuWf4jHTXm3an8ZkmA2iuECCueBl
twdyEhZ1U3n5PXykTXHa126I1tJD3fslj959Q1mkpJ/jaPcJRoYqOOkNJJJzyLlvbU2hcPXCxuKg
z5ZFTaDI5pp6YLOvmUGeVrFer2aMDkd7b3NbEAHNpWjNrgSFVlGeRIAF7IeFM32qt8jRsskRIfZa
6sDZ0klQ0B2YV+aoZl7T45HtzXJ90sDPA+XWeOuY2icp4ayKjYsrUQ+5g83CdfgB0dfOoXZ8mDj1
H/5vhl26O/z6dKyeW31UATJ+0yY3x07tBsUc0y6Wb1eLmPOFSieBolqgzktjBUaO9jEJnMgh+7Vp
Pnapdv3+WBs0H5SISDBvcKVJBoDU6V+1wJ2LTuvb7u5WYfiNv0EeOflems93lflD4NwiDUEMaQRY
XXV4n2NfGD/AKOH7kEjWVOeDZa5ivq1z4BgThbob7IkZv95ySgrSmx38NSRE4aN2nqeV0Ob18UXH
2MGmRV7wxF7zA7nKeDvtVhSXuP94tKRRw0JIFHY7vpHmXSpR6CCvpFi7yYQgrfS9D3CTTziVGZR/
fqflA9PRxCxVvUaBtepMPeVV8bN+K0bQnXSEqK5soOpt0GnTaK1+9pk5Lb0cQMGOunAQtfFDz5Ph
Fm32LK0516GW0sQyOqEAjnOd7KmcPpkwEsKiLQx5NONe79q3qAasfRHG2EBaBtlX1rXPP5tPcqHN
yoHXdM8jHr6WlX00NXbmvMm9V/CDm0Fn+Es8bg0moOGN0WS2vjDlWuoeuOM8wKMVUPoqtFRnjFeZ
F+EgDPr9ksoqsjFK+gx2cyU7mAIRtoT6o7TWmLwC9ClTFf5zLqHWjY5TpiGnR4aNkaf6iork7wJC
5KfyhVbX8yhqfAnghDJI9BwQMKI071qyXDgRL19QTaBWQCQTnQYY6nl+rcvIF3U6nlWCUxbg5eXG
CD3D2SgtkxGDgUEyL4Es+uPe5Lq4n4hJWDD18ey0qYyU06bfrQg+Rb6hqvoUs+T6XwHQN+VPWhFQ
watNb3vrZX768G2gBNZdUh+wbMF/QWU4Y64DVDDoPOVCroOPZsKlvZWKyi8cJ3Ne4WXawtbJEJiX
86t9kY3vwAlMYf/EpgPwV3q9KMzT+A0vUydopW6N5RPDhonH4UCwSGOXcz7f2qU/0vocESvi01Sd
fRNupyQ7SEr0P1lofqTeWxcF2TGqsySMNAZSdfUgaQBedId26S4zMt5jg/wdFBaq4KT0OHzOUTEl
Nsz7KC6qg3gMQqk49pT6sNL8PTHpo3gWq+gUnX3OJvss2A85azOKimgsFgGEeEI5BPUBu1BHLb7z
+cUkOpRnE3HPNvIvY7B4JwF7QlRdpOsl9TI5jt4TuX3I/Zuigh3UH0G0i9pzTYVPizEdGmiDSwnm
nLCv75zJfymra/AbPZ6QJHDLDez+Qz4dpDlqkZm4Pj7WPx8lRawVpIvoyNwiNhB22+wdtBjN82aL
DiYTmq4kKutLEQ0lPJOCfVATi8roLR61Y9fIL7206fQYPGkuzmzsdGMNMdA7sbV48/+v0i2dKI0t
m/A7+gsBD3QLkA9T4MNyHFQnzVT1W2lf4uaKsLOBQrnwXChFzPH2XCJD6fuxClP1gVqJuTKVY1L3
QScA444Kyc/v/wLQaGiqnuYEJP6fd5SV7HYKmAw0OmQBr790kI+RQTjSVJzreltGLAgSZcIERL8p
Broa9nVM4cL3LF9bNeCLZuqebzDGi8O/Fd4FccFbzP22Dg+fIHQNw2KDg+3bq1tScuy52wlK9JgV
+AcQgCKssebDEm3gPpsm1HH9irNoBQtTzo/uWYl7jUWxFEFLBOGCq+F1soPWxoqMyW+c5UudKTtF
hraNANYUYBzHWpWF3Z0xQBoqbYv7oiq1VJ20HYZPQ6Xo4RowYGnRsnYtoev5C231ONmHQ2MdyaUU
9bNzsznl1A9JHBydCvk7yWlYLvj2c4FKHUHuyuKwsQZWlUT4Ov38j+nKjHItErfM0Cu8IskpIg0j
kj7/CHlEIif6VuzNPcr9PV/3eDd1sZ/NanCjfWldNfF5Ov5o400FNtZh9++/McNt11SLrLwRtYtB
ZYIEEr2GMSiBwkxOxzyLSWRqazlNStr6OhLwlTmk/rT1YCCx2YpCYz3BPj51oq243GnwkolOW3f4
PmDc7l1bmsQdaIjFrrTombYS7BvX3O8wnKjSih+Q6y5I94o8mpsQlwnKjCdPhfsJf+ZE5nhL7ykQ
mFRbo2XmAtsnABaQpQAMwLtxed3bQ5igm8TE8nmcD9c2l1xwkQCVV9YQZKkZjPmpBrnPSH5dC/Qo
RFAhFIy8CAqvk3EsepkGx/XRdZnz1q3J+i5rhasPFbGKbfDRhs5NkqB9BYwubENOVvtwY7PKKWDN
iPkOqX/qMBk7z23BLuAD2BlLR3fjnWRRlmrF+K9JCNcbkwgg/YDEz5YnbMltVwVSwPvC+h41E4lm
OUrz73+yGgJGBBTDrL0sfPNIXQeOtRmFci67yq2jDcMMpoP2I9XUw5Cr0AGjsVO51DvB91a8BIZq
yDiau53IpFjX9OXcgQHD5SDAke4mDXXYuJjeQuVF8o2oLZ9JEyymQEvsvwKJzcAFHWXAurtgge+l
acNZUhWI3CXTh9tbkgex/TVzQEp8m9gRrgBx7a1jA6gLIGq1OICuP5KhCrsDLekNYWiWk5+7PHbC
dKLmghFioiTQB9po9X/dqyjAfQw3AxLsjzH3cCtU6PfE6Dwj0MArJu72CTvyMDqzdtEO2ADNrNaB
jWUzRWQpSQB+G5yolutvXjfMSiygNIL5dbSynC3wVjoxbFibVm2n+gby1KcTnLo4WaP/JSL3VAyD
i7nKteiUeFWHZJhd016uV0Qvu1AVFTIWNSdkP3rKqqNl2Z6p1RTemVahfeswwCUFOKBPDoKHePts
kmCOgcv3KUv65rWP8qlwyaJOZNf/c8QU+8ShwSw/fN1MQ2es2BP9kZym8kVTQ2KRuoUz3B+u+V+0
qJI0ixlUak51RiX25oJKdqnuSMYwXJSP0y1cqO8L878QjFPk/yXZT3QUEnzETFoAZB5zLIDOPayX
H6nqvmiw4ITi7c8k8podmiPP4YLedxUE8NzGDoE8dljCL7kpGY5zeKz5bvOC56Lo/j+ZbHpa2Ef4
ZhNRs9qgLhcxtU/+HvZN4TBjEy2pGY/6DLkflE6UrWQlJacUa6+6Fqb0Fkqnh9P585HmXBO+lUNE
0jvaJBMYRI4QdutPrtV5+hkYxciBsKcY5pf0sIqkZF+3X7gbpfeq8ONNeWjGFT07tdiq6MkTbfwa
8bQbahkER19ETCF8UmTdoPsWUZxfK5BFMrd77tx6ckIzjXaRtOEZtbZkcM2qQbUonaKwtu7EcFFp
PJdSLoEJR/B07Umpf4xMvgv8SriPfkcm7UQ2DmzhV0X6grY5hm8iXeeM/DkHNXv0OdBPnLZK2BZ0
+IC79sFsMC1W4qtEofLwDHMMnVDl71tq6EwKcrz3Qfj1Osm4Qbb/bkTbXEKheTMxkGul8qbGZS/W
reDfSL2XFwAlo3t7s/+tG8KJUSLYQFqRy0hMYCsVhBbqEGqRrNAtkuFvnI0ULFqdE9j6SPTZ1uhR
JTOc6p6ACoWAQXu3qAWm56wblXikY24DoAjTPxxn4kbxa3un/hEoTqwXgrxvTEYeXdhLxU3IN9Uh
7mQBVwoxGRyrC3dRqxrIN1iOIoMqEaRAWKTIIIClPhH51AmVSSi8oDhNZ22o6n9L7SobqsUW9ca4
sNu8zBwgn+ysKtMkJ5QFigHKPtr4AwAm7t0CbEsLj8g6WFic16JxVXuZLee+YzJn5eSFvjrDxn3S
8VbyAfDeOuJWFnDEJ9vtbukqfYvuXbRRRj9aEeFTHfZpO/hFGu0ciyFVzUdVxSmaNAoo0uH9Hwpf
rSpNcuUbAzhcy8HK9eG3eANFVzCVkMFO9dyt/C07/Q5EIfwmb7KmB45GqkTfEvI3c98oYSt4S/bC
uVAT8J+L3gG43exn8XXpZahjqTlpilZcGAvJ6wSpN4xDWgb7Ls/YptZ5Rkt8lPojpxIIYdvLgHUi
jtH4Q7H798DMpyWosvDuYJFbXT0+VKYB68uyoHrqGM8jNsolZ1v0OqNw4TmHnKEKR6vYqELW19Zj
whPAJ8FBVGcRYZi1RDrpWnpbHEuansNAOOdo0vWLq1a1xO6D0yPjq0um6Son+eSOSG6uYkdHohBY
iPqn1sSW/mE3nGeJghvGlYOgADktRiJzrVU7it/Wwyp4iZB8hCKQ8u57f1vCMms1lflDqkBq5alc
/MJ1/QaKlTjid3hnKJhYqAeh4QVDXiraPdmK8JSw6bMmNtDtWJcgM9ai+uICAU10vjprAMfqF9c3
owBeN42zrDJb3t3CL3ap6HzZJ4wE2qSfjAQ3SLne1tsgduhidtEVckzAx+r5aFmFXppx4KbQvwSn
zz84TnDqPAacdArgT9T/HexkKQJsTIvTJvQoivS8Tp93EoAOYeeP7hXEfTRwzurIm08jsmVnaqIc
q7Vj4MDlFfr06JwtM5FJmENAax01FbSUPw2m/pZvnfOdN4Atw2BkQSVGloV9yUtIE6MHlBoicxUO
r2sdQ/E36fANiCuS2efsxfmlokUykaFuWTlGWX8hNWVcay0wU6uAxdLTQ8R5UCKyKehJj4sib/8W
KM5acXb/bk8O2v0DdQmyv+WkIM1iu24wpz2vODYZu3af98OgVbjop3wabcy3nAjKyp9nUt/kTXdb
L7acjtRP+cnofWVP7ZULCkoGoeW+Etege3UVmXhpzU9vP5gT5yVuIUsQg4kWIRkdYLgAJl+kkSWW
dyVfNkIkAJk1gI94vh2393aGxH6SxyTeRz5gSYsLAmamKdBG5vUzfdJd6WjK1WN2s/J+lc8x+mS2
uJg2Hc+EyANzNVzEdhc9plTro8DCxz1Gr37CaC/SrA8zhL2JUVaDpZ7WRkwi/Cxt6rXqVB69WoMA
NqumZjYoShW8NWo4SmAMXX6ln62QM4stFBy8MZnJPCEcYYxY5me/vsLzjrH9OdZnzVVjOwN1la+2
KfO4XJBIaEKSMBRRcljqifbZq5AX41IJ5TBHaophXEnYiJ+pSfBzOEQJyjRnxxamr9dyQ8hYA2Lk
INPrR67Vfi9kgszCo2YSS4q3QEDebXhvY/TTYVq/oV8coUMWJDbRIlp/Cj0Lb0PVGm2yzw+sD/AS
BCycqvZe5aszbkmbPLVbgKtIU/KWsQkMGwyMM+qrDhdvX6ABfsDU73ReulxWuXuoTZkx+Cw4TsHr
Ixkp30/PcXFDixiI5EHnH5o3IG/Ss/iQbReRGinTBT2Vmdb1jf/4HAmPKwmmhNOCftkGWRiT97UQ
FKzCAqMPL7zynF3FoH0lJwyNP9WZCer74gpwAJgEYKPia2P8xTPxL41TBzwI154Naeow7mtC9cj+
qs2OH5FZSsxNGGpPqkx7aUa6KFvp5sl+V7VtHRN8F3tjTtt4WnwujBnuUujYFqdBdOi5MBx7d0r9
27UU1d/QeHim69kUJyglPYxFddSIiEEUQspiG2T9jBuYn3wPDHG7szqNLJjLRHU2WmyLGCbd5DLV
/kgXeL0Tuklh4c39N2/VQN20TSgDdCGhv4YI1/xHksMxM4GKJm55tdR9nJtQJCTbt6NgeXxC/POt
70zv7yLFM8HR+zUZO2y1mpBuK02tNhZ8L0kZThVPjtqAWr4PHpiN0Ub/rGSO8C9u6wSLH91evKws
a0RZPysQgZFeLvJRyu9ZxJf+1Lo1lxhXZtjrvChy5eZ8BXlxPJL/h840jllI+xs3xnr/Y0op/GgZ
N6udjmsUns1y88jg4RjPV/3AlKU1aVCiqSJL6u8abRPQQ+cV5ASxdikZURsIhN839/Vlafihft7o
NhhA2XCPhy04MtlCPozNp2BQNfWVIEpDRpTqvUt4IvoPYoIrrlp+ZcXURgIqg4uC5rCBWILUcEwK
bh3jux0dLv2K0d/A4i46cfnJ8fHMdsOjqS3TZka0HT7X7bzNGeAhF5KR1e1wpcJrwz0S/VD9CxA8
H/cuo6JugjmvEigdDWEydmiLOCWhRzMqgR6SF7qKMOHH+RoV2grdfp2ODohTweUK8lSiY87wnKnD
MLtHS93CsFCFzrPOJpcmJAbe/9NVMmT5rQ1uwAUazrb1zOfkY4g6gd3sbTfu8RvhjaNUjeuvjVyb
nNtZFhvspqnGshPZOSasBeD3JYBpyhewEkWoQwrOWdcnASlEljdxSRtMvN1uXvG8R7zDQD4rF9HR
waZ8nUsnAH0p173Q9UlQbvhn3OHXnhlJn/idv3I9YF+BkBKwEcX9kHVRiWCZgrHMJRQakzcVIzNO
10eJxzWdAKJcRgep2jE3RfLOpx8kiXsAFaGWA9MXhQ+ya0DlfPnz5+l8qkHXyXDsb6CPleDho5Ot
cyQAocaHhk3W7d5Tt85+fGxiZ+CxnRYqiq13LbbSt6xoYNCepJoY7Mbq3LFHBJxHqAttknIJPMQp
caaAi15A5H9wOrjzzt1HnKvBwNFoUY8aWRrVeBInpDTU7m6LQh4vVkvT+/x7rdE/T+mO4GFjIBcB
1Ogf43sNyxIMM/ROfw+w0jLJyNmV3+m6MbPwsRpMZb9I5BjMNrb2huwrgSSkAgOD1hYccZWMvvSu
s+EAL/QgESeDPC7u/KdS+Hh/lYoGWqGEhcwGyRTIrXSFLEgYzTGDEKr+sMwKWMe5uexwSoevKyAD
62XIWTOSjxM1YcmBRlnVOl+p0RnwnCoja05K+FjVRFcTtlPa9C6AAwDWSf4bHTa4BjLav4t5NfGr
Ck405SHYq1UVclrUWowIeW6dcsa/4qIJhv7WjVtGvFA0YA1j7iuycdEIAN+zPcV+O7S8JlGYxhXE
Bo85U7K/MPrf0j74DjjcC914rndUpUGSU2QtuIW3ukDMce9oUmDm9K/ERBGXriizsSd3bvXFs+GT
yF6A+6cOzwx4sxwQbtA7xteZ8CaxWt6lrz/rNUfWqLQaD07deK2iFkC+fMh3YsUsNgYrhIZGkgDq
YhxIgWAucMs2MzYGy/65iQbZEFtnecTfFt94W2xtbSMMdQyicbJQIcHZFXIrVmvPVoUIWOmwi6/A
T4JnnvWJ2p6ugV7WH7x7sAoSArPc9oKMme36yU1QINn2QyMXkr6MF81VR69iHOfGo3czxYCH302Z
Jbv807ho/wkFNS4WFfzhm4FM2gZagZj5FGGCScdobTAHwl5CIguboafjb6J/x+OrFS5Rynab2Ia7
qJtclBIEZ6XtB9MdknZiGwT4vVDG9KYkDzntZ0JNdptTsu7C+GLNJESx4zOrahhnvp7AZhOQVkvU
GcRPdqzLVUJY+nwegPMBGwZwQqGb29GYKDX3pqEbRI1G61Smrqta5Z2+8LLx53OvxdP82S3lCajf
SnYzUedFeyC/SQMOCc3FKVSjzgS6AXPQ6RsdB5bWs7kKqneybEFtAtOkxQ9eoyJ44UpUA8pmDssy
tNzGI4cqw6R2Ttg+Yid/4H3OIVI6/JgcBIJEO5610Q01oa3S+CuEeqiCIHn/QJVfFYIY/ZPVvyRc
cQ5+gf+8vFbfifQwe218jAFq2x+vvMWA5a7CRr+eIy/Xumz64aVlcOXPQvOP3wVanBVbwDVLtU68
oLX3LhGhfm830kSGStMaIPbXM7yyLZVH2qEVVBHri8dX9TXvEHX7xf6Fo6W4C/hlAujoKEP9bTmx
l+a+47vjcRPE/5JwlRwzh+H3h/DNU1mutt9arNyCMOb8f8kvPwCr+duDQXvIzbe8N/wPfgk5muAz
HfZDi4pRYFMzCM/9HmWChKM5MCP+luxqSuM6eqq6B7u1jTvN8wSuh1tI5hYhwPFUpiyvvIZb55tr
f+4Y8MP9rIV0nK1ewF1ck4ymugJnwUp72PyZpLfvpOhDrkIXnlIBEK+7GU/v9uPvggLW9j3w9YMp
4BU5dUMJti0tkPZz/iTAWrh0k15mnIM6sMIvzOVsA0NwJft9HY5M0pFjckZ8N95Qv4J15aMShXk1
jSVP6+qL5X6GkQCyV93dbb+KB9RfZ9ja2RySbOOsATKSR8VWAY9CrZSE0XPr41WUd/UCj0jsUDEA
s73+KBOGkkxuggIwSdbwBJ7wDy7OZJ9OCWlAFjqyDoN+ewnfGi2ybTyCvPap2zh6KovEJ99bQYpM
HQ66Ub05T9JXxRDiLWIvcFQs8YE7VDGEgSCxLmqnwyPhsc8o6Lq+WgfL6LEAaX+v2o8ZAZ45DQ0F
hZCA0AAwqPGYc8Ci0BfinmkVYUvT4zxb7+Ey2koSZCdnSYM/l8FiPsMZLtynOIHl2t+Z+ZyAdHjq
07hVBb0dzGfKoIB6M+EKtOeRKNbcJkyNd0tpWNP1wDx4xNUMwZ94X4HajvZWx8/2UKXuKIViFGqq
+afk3hz9C3U3FKrr9EPThi2nIrUL0ML0nlkI3nEmd33u6E3hisxXGUXhlNcUMGKI1j4xj6G6F3KG
wd+VK+Li4hoD3/eFMK2/Pf0bjcWU3dC7vAFLmGmYZfofasqcaK9w5hxx/T/qI/Rfmm+8iovuQ1MG
ALCwFHcc/3qoDu0X3q5TWQ3OMt4hblQffo6y+1qIMAPjn1B7nsZ2fGhuiMjRlsT7zjcZI7vfddJn
OAyB/RD6dI/uwa7UyO7ciJXG0C/AcViCNGD8S6xUcrEJk3cRhp1STcK5alXoW1UdwI26IE6SbBGJ
+/URUg6rFk3nPMcagzYI6R9uaOzO4a82m5WzLa6UPKH3s5AssaP20CdN6ab2UNC/QiB3fLsKDxEs
/8G3hNW9u+s4FbD4ZR1JleoIsPQEgjXENCVcvVBbBhBqGLNYG9ULixlRoWwDznZPtZAHH1b/pFTE
Mn6zimqtXiugI9OcZQZZMeK3nJ1RYtHkLn29hq9CTiYoUgKypLkQ2iMUXMbSbLrdlvfo8VbLWrwB
0mvfAdmqoCdi/73g3L3XpX6XQIdTANy83aUnSwsMak3TAy8RN6giwjpDejvBqIJrrbcRiv/Rjke8
U+mfGaC9v8WMIoXZ0kg4Eaz9nRge9ydyUyjRFb1zHWFS7Lxw0Kc+LPLNigYDrAH6YP+Z1CoL2TY+
dETt5VTm4LiG6GlCdDClHYrWH3EOR8dsz/aNMerhzRV6TjKucmKHW+TeaPNXYXiqIn91aYMXveFT
rq95uwQU5/pWVvDlfTZqoX2sJpxWzR4bsf6efewp01+NFdLDvr+o2cVMCJZSnU0g/P2IznIz4f/x
0FRXgGA9v9i9ahKWN5ueV00l+pb6dZANmhq06Lv/jM9Tm9Ii5uI+jJ85YpZ7+oyZeGGraQFe3Tv7
aXES5MB8FP0sXlI2CK2M0rmNuvCRgPfNWPr5rpIXS3MqUhNMGe3NWW1VmYdswdyNtWPa6v/7vqe4
RlgyHKYSpBh0O/JMSWL+W1S8+UjJS8QYEqvANSlwrqaqpZH/QQFDYVo40qV8NfOivR2/tg1rJ1Ia
zTFRS7f7QnO2SbbUcwTApoCwDnmL8q/Y81ZgAzQxdO5/H1taD04PcGDNKUEYLWcpGVdxHC7YRoEU
MIonqcVNOaFHdHRLJn58OACLmxbFmV0HvCnV8zrikN4LnBS04TUpYZjxpaQDehTuHh6ywJ7Cy2Dn
KsIKb6GUJXD6LcC7Iyq9btzuWM0zGRxpbqEzWqP9Ku/9I5cF1PcoDu87h50LC/JimZBHJWMrm5M7
4dAGEcrHzL6vlBb5RqRQPqBYrmi2Malz+Ob9liXp7eSea6fG/b9Zlt5wqFBWnZqs+J1CTyEuanY4
cvM9msSU1wJ4z3pgZaUBeYskBjLByfPHAOLnmDrlkJMADLO8/MI+werTpr/GJKAcM6X1xN+4khCH
kiPQH1aZ4+g1R44ODSBLqgIoLmw4EigylNhfe4A63bu9KaE77R2G8a6w+ilgWFqfF9VTnuitx8zF
KFMZuGfBICLUPDaUnhJHw0HNexPLtW/Mf79T07B0Jnn3m0aYVPyv/umFAbqQJck/qGNkrGsz2BsE
dVwmaHRLoAXQ2Q8REGd2wPjXrcTuShCucLEAjq/4z5y5JhzjSGmtkWJhZUdn8Pe4t6a83B9A67ep
Hzg/HZcAB4Ag9UesA5cp1AXjmLuhIrt0vhdeAip/1gyeKuitxCI8fmBjkyjwYCWtgp3y7ELsOzwt
xYSqP0lViI8t7uKaO01cUkmXELxHoG7Kf/+09BWsGYyAk/RnTARrzq0LhF7Qb5JJ0gVyiNUoHO2e
RSVuHClWo6R6tOKQgc2A3g167M+r5pSa0ACP/IOjjT7SHNEBubybnnghnJR9qxSTZbsjfyIGc+cZ
XTkeU1eOFNDeVqupB3PKJ4xbWvYJkG03cBGcrn5WrVx613dDSJuKFDq7vgM5i+L7nCFQedp+aHsK
w93CgosDyQR/JbGriDRf29gmkC4xacLPs7LrFjOSbq0tNGxDcAKgAYbWfX2BQ+ex+8y0WPeG0gtu
gGuajCQp0UoA7esyalzbpYciywuIo0K9eA0mm/a0HvXqtfJokDoie0he62AuWBgGd9uXs7uVI1+D
kuS0jo2JIawyP25P0w2Ut7RV8ag04e2tAuqsudCq42WgX/7dOMLHwSHswgwFQWK+cj3243PTCTdl
z9+Dv7dahpPaCDiHHNareiDEaR0xNDzyapwDviIFFyZ5e9jP2xa7t7qADWxJiGCULfsiysZqpYNR
sIzJKZldPROkhSbVNSPeyB0AzZ7b5I38nd02fvZ05FO4WqSErEW8OLa0mpUM5/QE6jvIln4lC0DQ
7879um2elu8o4etUh8sC1UulpOQVaLffjRgDzAw34aUwBB78jK0ioCAFlVhonbfcx8KEHl7Wg2De
/xyKMUtxDGvxm5b7KC1KoNHRu7zkBIAvr78VqZeO1/ts7rUUZsS0tIMz23dmDPseAX/iAAyUuvQP
c7aMIVKoqmjib/at6P+WKAeSYRmkCJl6YCFosCEeX2pezAQj2Vx+xBTBMNP7+35pFldy2RJCSxho
RyPJj/1K9vHaToOqMCUdqkeWndfgONvmwoJdoxp3nbUyeh1ZOjxxBgHqYdAJkO0H4h0l3JwYDkcQ
xIhKj/WuYWsO/32VSwlLT5HGTWbFxrnvEVzxskfJaAzxmZJntZJtTndtYXzSqKGJgJAZZI1xYaZW
r0Va8+GFPKAug9ILZMoNUvH0ldXQAKJ9ur2EKth7wnUwC/t1WuShTcAfJmOzp7HbO6y/QUmU7NWL
uGAYBSdwVnzfvZIEn5HcyJ3K7JInNARxainpb1kfAXJPxoznJnTAX6pUOcTsslYkXhIIeoBf0GKL
qm1utnKhsh/0RI5zmXToKh4ohVUSN+V2ymiko6Ivzcsu0q4NwrHjcCkqGWUu/gy1Gbwel5SuPFQO
BSAO5Le/BorZg6PCSLWD045WvrASGqC5SJ5D/DZsLCQsN3R68H9Fq2VzYqwkOibHr3PQKMDSfKEW
5vlIQCXFlzVDatCg6/UbOJa1WkJMw1emtW5WFggIs/Plktkb3WNK1lcyD1VC8Vuzng416e2D25eI
ZeknB4md4FIivs+5byHWLFvcHPBSywIV2baEgQBsKJ7Yyd9UgVYUhUDZnkOH0dj6N/Rti9RJHe0X
HUdhuA546TbLogV91XK21YIzqoWXNDt0ksPnAjFkjBqKpqwtoF+CUjc8A6Ov3HPKH3cKN+jPgKwM
EbY/328BllhgmVNq2LhdT38uTUtx9+r7Tgqc2ABDEJIZ0IktRby5YpwwNiTm5FA0RewdqjSE6Phd
F0E4h/DB2icH3yduFtplJq5uSbHHwyCJKp3wv9pH4ULz0443tmYIxyMcQY+naHAG/lFlcqcEAeHv
Vi4tRn8WhhYkRnmT8YDPzbqWVSledqu1qPqGrHdliCo2S34nYm9PE96t4Yl23U2qB0WN7rDG4Wmd
1vt0aBnhrFQfbtRWBpPrKpwqWLAAsdPoFUecQlxkJgPiIjeH2NtQFEd/Zev3zQzpQngN7p+85ts5
0ypMSYlLjIKmEXA18sAw4M4v8Km4g5NxJ6y4UJRUiWzRBdaz1VUR/Vz50jSgkQkSfLDmNrR1jwrf
c26BQNGvq8TqtOfORk8bjvGdMYW53sfP7KuXlQeeNhFJEtNSQZDvVWyBLp08qib5GiJA82jZY7KH
uwGl0F7UeOTwiQ5c6nURVoG6Ic8kFPkvSnAhaebDaAP0EtDFh7AnthWKuo352y3au4fRRY4BBmD4
g7EMzLo+XGlgo9ller4rQGFaB8Bk50OsFyB5VK8crZHSUP0zps0fB07eMwMSKdaz3JQiJBpxBsyE
iwhFTZgqQUtgwmzA4Cxceryxebe83i3JR9CVqNNAaxByLetUJZ2kQo1/zZjU64m/wOnFWJzjxqxo
LlFtjuSdbb3LgBieWXBPP3rzYp4pkTA0cxqjTKAeJehvYT9dB6qvzQlG9w5FZUjXCjflx6a/nzI5
7dHShb323JXZ1ftupCZyU4iR8NJ0B7KaEeTzgoXi5D658pAbVO67r6dSG0Yylottfph6FSuRJTZP
+PJ1dnEAU4deSyMmEOZfRcYWruuyMUwQQ42ze05xrbbzFzZaCKdwWWj5tGDgZcHRzkWUsfuhmUNs
OMjn/lF3Jq+E7xZJPsJ4GquqNRzmj1eulcUifxNh5L8nuPZaE0DWtM1N+3ysqf7lk04R1ei8dZTz
Z8y6PYxo/1+pIGVV185LV6JEeXrTnaAfPOjHmoXkQKBKWQYfTo1IV9JCBfiVg68NlpJsOSp/PzJa
3nRSCyep7nk/hWoU3gVXge2bp2F41WFP5yWkTIqN5DlALXP8sMJBjs2D0/GzlJpGQSh8S5pHT88k
qe1c9hb8mWwIC4Mots4fX9VeW5KoonhclHzOKVOzxU/LnRhJPZ7eT8BlCWkCrsBWyOuohdby9Wvg
ElJk9m6z7ceIcWDQN8bUf1dW32HBdZrtfrVNkFgwa4ncHNZQz1M+xpvjVeRQJ+6yct315BEm1Tz9
lM8lM/iEK8T60rs39uy4KejyfDOj7hdWlM46zqlt7wSaD8qyIUJelSAjvx1/4hL2tK18VuQvw35n
qQUDgz2hPgPQ3nsLJKYcmbMNUHknQ9hGzS8LUFtB+3flbt00n50fMLSEAeyN/NFHWX7kruk9Q3lG
RkVYusUYioXc3iq4P9axnqIcB0fNy83pbwo0z34MovsFEkrt7RdHVpmg4vfiVo0Ae3rmImaJwHDc
7/4ZpP8bhOBhltxk6nSaJQd1/2V6O3i3TOXbmE4017vTyiEs1ngUue/Hs5FGjtHCugDppQsumwSy
zDsbylfDPGQukk+6vm3mHcbpp26qPxzf2VAVyemG6AfedZ0w8oqVxIEo7tB2J/IzWtGmZnKbfKhq
t30vk8YFx30Y7QYpP0Io9pxB68QLYuHuut1YOW4e8hIUFEQFD67vMCUMqOD94OI467qpdZHnSpg7
m3ep1jMg3bWJyStqJBv/TQPvRqMlhIBJTb26LSH3EB2YOHb9G0xuWZlO4qPZw43Uj7SN/7lU9fne
Y7DC6j2BZYJRforuNx6cChDgQ4UOqrFbTfFza9S3Pq1Mh7+dAzxkgztGzae4KGgbDEbfHxd0h9Ti
wL8HJVvczCektuxQD81uN3ihHvqnYwp7Djg535S3189mK/Iy8LEatDNbxYn9w62tVqGHptSp32gd
wt9sDAgLD9odlhrm8axgInHknDUMyj3uAymYbmpOojgrINUBZ/2AqcMBTR1qX9LyjpxtRYudXel8
bZw7nyWOUIf9Oiy3Y+WrxRinKQ5+ZbOANMncT1lx0y3FJQJq6HFpwlPYHI54pgb2EfWmPp2SyZRh
5SQ3vzfNI6eD3BUIbz/UMyx6XSDrDoAGFDrYy53TGuIZn9YzeX9PG8K1ffjkhDikBRxyze+hTSUM
4KuOTnXYvem/kCiVssF1O698lB2g18mqb9Iwdb0yJC5vtGuL9HKIfpTMCx4M3OYkVxNuOcGpHHHl
fUZLJKPyt1MN5hA/ICjKhkoKoJol4zgUttMDRX/g1jhhZ5tFLkFUBzIEqd3p2cByfNlSABIrceHP
9WS5aaTorfaGMs4laMvmFYcMfygIjv+XVy8fIBHExiGxLPuWDc9GJQtqPH9Y4zDXgei8MQeNxUfE
VNtpRF1bndFwmGYSGkNKvdgq7aaVpj8UWST1Pou5+ccFwWVCZaqLCJAMG4cyFt1da7/Y8SBxxbUe
sDZY7Z1rVjuLzEzako9K28kfrVe0+5YDhUPEbhL3oZXu9cBoirvVrODcVL0Pd50r2TmjbbUGwlf/
GvYgFRJqupHrmMHb7R8iEx51gWuRmkIPnnZJgEuz4xqd87zv+416+7GG1wBFItD7EKhGXdZ+5Gpn
2LOz1unHAok6Rfvz6Iz2JOHBggnLl9FCdujHPEjwAAhJLxqmq2XRyTZbjq0SLFsvtCrjBrSh2I0v
zKaaDin9SQbDeKtVYVJLm8Q7dprKa8xtY9M9dJwMxJ+a6pjiD2V1D4tdKilvzxvSE+W4exAfPNCp
ww+BBOLGf9Bec3j1OmOLc75TIpHQotb+kTGDw6pENJ3ynb/sooeETyTDyNDqXEQTseKRlzsFLBGd
iR/3SUZz82HAkxbSmjTgnYlB8Sofl+D0MBC/xmxellVqgmLNnAeArK4zJVrdFWRJXVyeAVIh4Snn
3ygVjheUXOOGkNf+bftRYTjjK8K/naQ1B4rAViqaKiTgRkfr0uHmWkSGI5G2HR02v64m5Gu7LGJT
aURAynhx2uM8jBHbJhDKvma/97MuU10L2dXZuNftBR5Pv465FhOd7LYTfEpJQTf6QqzWoahW9A0g
XQ+KvjHyB5PxO8Q+ktLlFpMk+yEXl6h8L7C5O+VKVXgNfjwrcSVXjOOr9yNUAfXnXdLM7RMIgKys
rTckfkHCciy1ENBulkqNm6mivvXXCwx1VAXGSYCPO8yAo+LuIm4Llgd/TyDhf7Q/EqSGZopJvHkM
7T8hgizRrbnJArb20h+4gkAnWm0FobjUMN034BMY6vRKaeqxApn3H8hKZL9gxgz7Yvn6IY5Futd/
zJ2dtGvgar0z9k0V1Kb5/3o8j18TltUIilMqpgLU86hevWRLIEjpHiNpJRFt8G8V6C8se0qCRW2W
Vz0f4+Bok3djPDSitKVazr3nNEHQfKuEkRs5cGYC3473FtW4/fGhwnglxY5jt59BM0GzE0uwDi2m
JIUFSb837o1WPU4YlKcE+zIZotwAV0eY6IB2Kd6BbVMwJt135nsT8+oyZGA6gBDbazavi7fbRUIQ
EcJQsKdd3hVNGZJuwTIqZ4QP/9M7CBbEXDAQhVBFZPAFUX6AERsD7OG7vnHCabIHmg4q/iA5jAfo
2XF2DGr/JDLnryDe1OycWc7UHqDta3jdUbnFHzhyKB3uBXaY83KSqAPiROLb6w8nHhnvmKkS4gEh
yyB4Fwp8qO4cbiY0FVMV3nRvZLBvefoPa1ERkLL6iFku4St/fcNZgnxK3pu6Rx5UoBPafYsKyxFx
v6c12O4cANDX4IKbytjjUM9yj7MNWXuTA00N3XUoIN3W+hETNNxz3QCsyokNQKsWsGEITaxne8Oy
OYv7toQZ1aSD7SBpqBiOBrmE87PctXfol1cChXlJbZKcJODlFZY+4n0VPLwSRB301mu70b+/j4Bf
jYpPu5X6wo29cSA0YhCUns1+/TgzaOPeiR9MxwnISUpTJlDVXl6+/aUryN3+n4dozZU9nC4fKere
YZEV14uhawzUtsuMG/kWeOTWKDFVkaChWPLtvL6RrZSesf/FCvn0NhnuQd0PmXNzDf/SNl+CUYd6
0TciHZoC1rBxGI+BigkISIJedMMbodySxyAdLPY2BEvqbZr/46eq7Xx9bgKm9lYLO/YV0SIehDRT
cZ+N/Qm8+Ccjq/ciJiwG+GhZ8bLD4q0y5Sqs5jyktIbuI6Ie2CsSeXO8uGABlHgTN3M2+GAagdm3
xl5QpDmYdYfP1aq1Bck0pOwd4cvzx82KhhvRsEihDdolbQHzaMiG+/7ooIFUVhmNnXU2U0imC+fT
I7UORFnrRGstrqRNw/s6nEqWcqqdNSU7+10JsZ7VuXa/PkSZgPwKEUPuXZqTNNIRnHeZ5D5Dd27T
zHDKLzmY4JV3GYO7UHtd8idueugH1YhiKuq3NGc4qdbyasc3mQtr8G2i4vu/gqnRip7RmO+ka0Sf
N8H9bI4yau/olyC7d69b8JNEtdcQDZL7VDmaT8VDKfEntPDe7HbE+eB8jdjKhTWV3ZrQAjB443dY
+mHHN+cUJ6lOEaYx95yF3+Vyj4i0iJPbmTr5Z6izGkzLRyOVBoNYmVZw9UsOSZuJqGJcby1dcRct
zr0nxyB7nseKuaQiRcTzMW2v7QiiijnvwVWcqaOErzUsAsmm38k6MIBixoamCD3jZvxNovrpWW37
O1Mj9DVrDuIHUM5W/ro8qmclmyd6q9O4thKSgZ3Dok6lGmMgrj4i9/z4HO8yH3Dzr6qBW1YMDLEW
8rcXxu/Y1dB89JPIOMTzslKNXUpMXJ5vzx07fpiENZ7hYANYZ65UkxoQODDCdPtBFk/5DP8uH/Ku
led9LWngF48L1IlBeVIksRZRmkAJbbyU3vr/YFg7ql9rxJ9UEM/F3l6NHKSLROP/+VBZyY7IzCGe
3V8PYAd9t78mnDa2SOcyzwI670GgSooRIR2h7mPm8ySC9IaFlsaKMQosFUSY205Yk+dE1cVAbOjA
q8/qfrR35nPVXy6G4S98NRBcmPQSfQx3rM1dURlLST5EyEigwG/aiTi6Zc55v1hYxsY6V+Q0cxAC
v4Ozdmy+FKI+XO1VPpmazebxsE7c+9EvtEgzTZCs8wwiAZQd1yxl1k3WsZ/+aDIayoPQkY3iv3xC
Y2usKWLUvHEBGX4OyYQbZpnBNhViGDeXGvj6whhHX60QDGGfjucnyOn41yWAmSI2Q7DcUBKR5sdt
NqhhtFLhWH6p+5M04BXcHfCA4bN6+T5a3kW5epamF8zrQI5pjVM0NwOyLzk05ARA8qbnZ8wiBHY0
678dtpzfm6GCVJwcRUCgAIQN8Wge2t22IETk0jv1RxeFdTAj8lhGmdFnnamxcwzEGmFyiD44FIO9
p4B5MLUCb6BZU/sUspf1/pB/SJXo6SsTk9QuBBDoBzZkqX8BOmoP9NWPtUGy/wUPi80QsuTXdI9T
FiwKPWKXYuiOQLGJ93w9LY38EfRb6jIQHeqwgoVKpI5xSl9i1t24uoap1uYUwXgrPM5+2cjAww7q
P3BlhLOmPEP2XKqSkZxWrxfbLZyuy8O6osFVmFluQFwzMuRTxhzTvTxnkJqWi6iABypwdxQ3d6ht
1yF29ULGDvpyVeHg4RscpZhp/YUU3IrE4YcIJ4S31TWFjFP0OVQHyDfWxwIElZeL50+uOuZmiAh3
+D3+tUCjbxQPfYANP50vnJv/TQA3JJdwLutpDRSaA+rL1jJJV0pYVLccS5oSwMRZL1fR+jx7yiuA
KqiKlKlQiZiiHXWxDZpm9nCXmCEHJxijQqCOucvxmEh81WBnKaH/8Ozjvak5Dp/k9a/+r84swsia
Z5MTvMgREM0U84EtJTr0y+owvMB+IPQ5TVWrlE7ZCjFx8rl6BDdlXF//rSFnPTtnFgdxCL/xe5y2
W1ZKIMP1YS4lFMXFw1UKUBUM7gPRDZzxm8bla55HrDifEDrFCiNoh+pPDNpCyQIlI0sE7V9i4G7j
FzXJccuAtrj4BM0J0B7sHyo9DFmeSNHuMLwBvKA42OnVWJPoltg/O96/XIcaNliBs1uID+TbDhWg
5tQrgLgzyuda7JtCS/WNfOxz7FQbe/d9O/KB/gPJuY183RHawj6ivTiOEwX/7QRW2IMaSwz5hs2h
dXuJOA/EKWkES2zHW0vW/7jMUxolck8Alb7s2Or/Qx1ohypM0DaPxSNMFVNmAqOvJmXHv3lgc4L0
qyvwMpimWyi4FNrMzaR4UL/oIpoywDwnCSyJQYbinGRKdg5rOD043u61782T+M/v/LkilBGnWLhH
7L8kv7XyDNFslZaQc/SVkcW2hgC0eX7QaLPUoEG6L2+vmh9p9WQdPYPK5bIdGneSMlYNjQ71MXGj
kh1pkwp7QlUKZ8W8gxWgULwHYhPKsxmWn9tDRD+UOrMr5JwtBzVp1asPtW0lLiyi99KZz8c+6Ewt
NveATEAKpRDxDzssOn8rXJnre0bb22Ulh0dfqhNURLzQ925BSUh3RIb+0dva+teRD2owM5OnJa+j
oV7W2ijniopv+GyZVERlNgSv/WNdaMLsoI8lC6KhDrQ1UPwAqjOuRnNhVbgO5JUkmAAUiWmrZjox
sX9Xtmea20UsEmP8n7uN/oy71xxXgFrps6C7i8ktU2eUiOY6QcZfwIlBsYkGjveUhkuD7atsBcPD
Lv1Nwc8ZKDX+GUar44IMqzRNsP/Bi6sNQBIsX2Ox+8mOeGlWUmjuY2tUCG/X5MX3NjWXL9liA9AQ
+LGEKr1G7/SBW4/6bk8JO0IP8iv4Gn+GEzcOEG7wscmFk2ApZ0o2zXuO3q2RVtu2FZx8Xni9PVKh
2Kae0sWV5pbsRaZ6cTg4j214OeJizjJjtihkCL28Ovl99V1dcjgwbN1OfiXKXU/wveuOmAPCblhW
/nwfyE74KYFlGrs8eJtHWiNMXNYKX7FCZGmfhQ5T9pDbQg9ZpoMExV8NIgLi0fS9AIzEI/6zG84N
HzBAV3RZMH0FclFNAKwBJ6wNAnpu1dNFmaktJtjgwEzFT9el8jz5fSjIZJNGpziUkYIgMKWuL/Uk
SpHDlK7jHZ3HHfQne8askb99uU5z3K6KVQQyHNb3sr86Zc1k0DQujlsgFWXsgKqqMMZx5tDJ5thb
7e3DxhDqgfR7/v0jOgd8vNEk3sjJ+S05bScCHSGNfimCloOo81AQ4CQ53JZIHo5d9MDrDzBqP6FF
Udr72AuY28uGdCzuNxRKIfkZg/JTEuHToTNM5NnJcAWkOwA8dXbAy4PmPRclXzAsgEQXXNLsnUg7
Rkdm98+u4BNJ5UO5Oee7Cm7ZUbliTxuufdJQ4R1xX/y8bPW/b9EFpFu6Mgp07DJ6EEf09O72mlrL
7bzZppbuonunSBjfo8l247X5rsoa7/TmL+3MJVVwvAARAbItOL6I4lrsU/SSXdXOPd3ala32diSZ
EdTEYHW2xV7jJXT/2kAe3zlomPe8i/g4GfLrOsRqJR3DKwxlcY5pn8EJmBLHgLsFAQqde2dlJ5Be
Ece1frQOoqpOshgYX5nKFT7maLYoEo+dEnHX/JAXorse7PGe6gWs4+eEAyhjlhx2AhcOx6mZx6bj
1j0+avoZEgMajoD/tng6jwh1ZxNIp6GJoYYj7LPURw0u4k4gC7QrilKkDKsnChFuC0ectV5G4cIo
Wsa1FENKWpz7n0W0/Kw+tOtbJ3xb68WocRHfidE7U5WPvCPUCN+zgkKpo8qcNvQb1z46ppU8r622
bkWcZYGXdEEeEbjMHg3GXFGl82EVlhOf2d9Yod2WGwJPF5EPZ/yz2JseZU9S3oYkZ5i/kA8/1lzm
SneA595m9329caVlItCr5NdyVRfvbZtMjCCjEjT4bOQ4HnUKk88FEksFQky13PGcVCxtzGhE96i3
EJyNZPqcQy8BGTqx8iDjgm4quvkTCaL1YTbg4QCeeFn6Wb34arzKRkE2B8DVePpmiRvHDfOUKP9f
g6CVRs7OzEq8nC/I9ugFY8/jhNshwVZcRK3VCcF05k0TT/mB/nlYIeU4BP3lnQV7Y3rsElXUAhsz
CuhUZRVr57HHMTLWbyDqG2Ar31nGHix1UlKwhzoq7+O4MekiAdC+T7KwV1J15VCPVkTaex228D4d
2PgBWRVMMJePeiXsBeHIRUPWReWlCW4YeVI6l4pumAF9ddW3DvxfuCnF5h+67Rlrq5MazReXPO1N
Y356yAHQIVPbfgS4JTLNvlruItz1zUcZXuLzRHUO9RZMajyiBBGHKd6sfOAhEQpn+6PQ8MRVTj4r
AAuBBZ2T/x17uayR278o0faeIdIaTQCPJ0P1duPgWgBcuknga5cTo1iRn18VCxNW3mg/nyKELQRm
lIf828SjdVejiYNe4u8mlNiPTRuI9aUlyWa1Xiabwk6eFu1+PuJn+RK7uezmGUB3SZMn9Ld3U+qe
k5wfvjhvwJGEXayt8ytghpO2T1nLuGvTQ02w78rCVyW6uRPsPfaLHhbtbxqFsgCGiCP1crxyY/eo
dNZpMwjZgDxjLK78C8dvWTNfmWRRZBOn0yVIcs2c5XDDDmYMTOJ7j9dUGeCSOYPOSgCblg7+hwwi
ztM6AbLpCFwjQ5TamWwaqNkeUqnJN4+zpJjyjZyOKkV9N5+abCbXJU6DW2DyNgvEmphCD8xfJfYs
8aV/E7H2hdUcEojowuDTHS/dTeeQ+bfKu2CctX//eS54wY9tFO4j6npg8Jm7xPmic+xilsHoBjHM
CJD1hPxHIYqLguegjcLkv9LuiQgCFz2j2snPHE/ed6gc2Wx5UJuUfx6Enr0NR+AQ6FeU7/c6r/3w
FFtA7StQv/Hm9DVVo0rSzoaHaieJtG5vuom1KyGk2sRg3eYYrds7RgUCc1Mcj19TEBW/BaIafs+6
8bz3IYrJLVdkOkLjTAt05e3MZ1bjo9QkC5YvnhPrtaxi4PRTRzaEZpB+nzWgobojBRwBWXyl2ILS
2I/wjaBgsLo+i6l6lKPja6/l308UK42be0O3ixdyNN6Wl+vNKTw+0GIF/S3k7wJIC1yC5zIldDi6
zXfkrEevhNjoZODrWqIIpJgMdeP1zoACiMDuYM52rnTSd4ToVAhERkEarvTv2TRwep5FTY/vLols
ZPDeNHzt5/RIRuX3PpoodGTiF693qf4fcRGCRzY8Vdc06FJNmztM8UqoXZSQ53hC56eO6Z5Vf2u/
RdJcpusr6ntFXahpB9X7w/jJZ1WmMSZvSvZPpuLQMZByzJYtq9b/yMyI/MCvO8Dw62NsDoE7ktmq
LG4LRhFFZ1N/rV+Cqm9kEFHcZNREZwJH4TUpCV8Sdod+v2QyXNiblmRi/NDLx6ZIje30UWBa9Xtq
JSbL+FJJh80fVkyl/3lIojuoqN8NdXQNDBszHN/oxVD9VhkrPtB6jrezeROOycsVf0TLZyxTp+yW
cVJrvGrTcfaoEmlQI4ziJJ5qKFrZW4M3uotKDpcTbWUc5BWrB/ODD7MFeo+Rf5g0KQyyfws01Ay4
lmy2y+qVT5ARavoV6Cn+3pdhyK45b1wJoOJuLOViFh/hLbFSTnal265oxSltQnLAorO3/DTo8LiS
WTkTou9T/bITbFmeC466mjV1aSsGp1rm5cUTAQF3BbYJXVrAorw9lL4F8zrvdNUnINk2AHSK38d9
C99/5oxM+4SEm4b1geEdIbNhSZzGF3ZVZfHAiWDqrlxqiIXEq/hekOnAdokpUq1K40jePdRWkjEa
lr49M1Y6NR1CLqID5sgu/rvRqkT85hR4uwyNdDBinad9ewgkBr+o81PqxS5RCTvEl7gxOFWwmmTj
Tu55Muh9opLG0nHxi4+cWYEQS5qXVO+E5VzQ8UqD3ZIfJWTH9hxCeQqzlLIiw5z2FzD4RqPaFJ10
PZAMUG8bRBrPMGf12+DCDZZUYra/DMA4e2KuqI9ABhNk05LToL4aFV6ls9nUK7XjfSF8YntoHlAh
81IpqMkhc2NqfA+ksEaeDz0jixLrvFZ/HDZmVWn0iwEr7ScwiibzOyBhzvTDsYaTBRvrxCFkJ2vR
4R+okHB/QK6o5UzJW1P/szESCW3vVJq93oB5ugZoiI3Md9YzJ8F0M4h8Y3eajDA6Tj47eJuRQRGn
dGQ+F/A1hYltu1YXfxgGB0FKpYActsV3ESvMqseYUuV6mi4PaH3dwC1fKnnRimgR0h/iGOV8y2ar
VvO85ZrdEYm/Pn0jA7p0+LxOQRbMIADMpwuLg8hrthIsvcMBH0jmflHCSoSqv/WrWO9SFMl+dSL/
zWW3bf/5GI00vw65pj6e092unFRAMp3+i3e+GyRflmQM/t6zp5+Oy4WRuCiT06bZWEtgDr/HvIa7
WYOwv7DN5SRGW+0B7/lY3DLysYbWo+6WcK0r2W0haXBw7KOCFbBftJMNI8bZvZ8z/dpIp3PzO/k0
/1mSce66eZjF/k6JZV23adXyq0qotmCB3tL1dUgIy16/HeQdIy5qVnAofSULH3cRbbyiOkkvXiYF
GtsAngxNa25/scAIORWAiTUwdIB7AYh7+WYNwjX9R0FxnHsALj2ea3C6ZoKpSIVwf2RbepstvDEE
ftjeOhrfamQpc37eiZPwWT61ZGeq4G5fYtlncPr9GXSSy496VfTZjhlwmYX/PVEGyICXosyBhmAt
GSPikHmoomaWtfLUuHBkvUZy0QvGX3o5d+nhOucdxNKPGM0Ru2x1JHPUlx9uf9r4jI678BSRoPsm
p6AKqF28QQU4AAeR+/HEpvsimgiP+2DMDVnwScB8P8Jrx08wuCF2hYbrB60DDwoqZZGqdlCDDgCs
+5+E7xuebqIdrvFsDAmRZu3D96G8ecuaFOIERpnfCg9SrohbOt8mnOkY8rRz7kMaRKUttNaYbQk/
bKc77289Z/ovMHNciBnKb70BGyovE3gyhzf5AYyK/lHBdkQFOw023LAcHHQPEnrM6DXf4gb3o0fP
pePWGi7cTQ3M1gIvOG1MIEPtp0bRR6yLnCBUyLv90DvvhW+k9T5PEw7lX8K94TZfLKYUeMalTPxP
bi+i5bGip58wxklBTWfqWFAadMX4mCY4z6qXMgPpZngMIk742yzPEgVmVwAXxp/OimXm9lTHszBL
oIZmARlCurafI/zLxW39uZEvaiAalMU3eEblj1rtpE9by1cjEx7EdzeEzd1q7IJAwQS4Hk9Li+1x
eHVhmlZU7/wDGu5BJ+OgO0MT+F5bwdRUq4v6O1w12slmEVEaLGCM22RUAFNotPAF33XsY1RD/ept
Klk3T4Sbf5I4fyvCy3XevKawnrshkdBwfllwrXYoajVl5rH0phbYcpzKuL1ANNHq4e1KhMmdyb93
1bFinEWfI63R6Nmod7K6qfzgw72rTqcCEyVWDgDXodZEipnb8Z+NgjyroOmZVJPgO7J+OWP+Tw2j
mSM88QAREAGtLBCukGLCYcxpSjm0mndPscg49uev8qHjGJtY0V6doiYWvxsOdCr3NkZ/j0wqNwvP
bf/KiMQHKV7J0cMvgjHQSBX65gdoomUY9L3VzlbNdKdKU8/obA7Qfgfht3EwESwyyCdJpE5geW8G
64BMqc3PTMxFpr/kPpgpLvOXTDCWYNJ1Xh9Nl9zFEFb6ClF/EWy/LOnBpO7Pad1fyOWifL/bTEvq
fw5sTrB8gVCrAH2tdeBiz4V29m+ytpZvH8fuoT1NmJa1L65tD1BvJ/EZSKWHax2ozClXLyw/5DyM
ZspZjPBMAoBp8yxfdgPH8CwEaVf4orrTuYrmFwVzA8UEKjTb9L04wVhuWrmtIauMKUtgvA9A2oYS
PKdL/t8ereo/sjC0HTPRIzEoGL1QqEtE41aHuElSRvBrTE5/JC0bLWzojowV+JPKs7Fye6YdDOy5
jOiNilayTSujsrBsC5761tf4Fdrs/Vs02EAKUDaO0fpw2FlBDEt0ZpZx7jDl6X7dH0mQxeHMd6pv
5i7hTouYKh/Dpwt8ESbZgarywx5tCjCI1c5PCI5Vid2xs3AsvSKT/l9npLD5m5u6PqKfF8HKYtyh
dOaXxBJEDUwlCRKuNIG1QkfC30q1J1EiqSbqmu1+zapPGxHhXlHuxjApnUXOAKOQbFDOv97LuPPM
M7IgWXz9LIGLdXnkQM0X3xmnHPVQM5nJUYa4CTC7wMLEWGTt8aYB7LvSM3YtuOffT0myww3T4XHf
/sTbThaU0ypqhE5agKK0/In1zoYQ2yxMVO5i4/y323DGA3vjG8qO3qYOqTHPKxw6Th5Irt9FrW4n
Ak8DJunC4+jHe5Cw9D1Vpy62PP4kjx4KAVQBJF8Ixms7ZpFM/hV5+PWc0MWGAeQ6d/DVd26t8NQr
TvfFrenAWGHw1fSRIDQjIO/JpQ8LR1gwJAv2YoMpNresYgnTEJILveeZQAAFaxY+Ft/8st+BUP/v
beSC52VLNJ1bHnQbfScHSrJcL/SSQG8gMg147W052FTabtijPG2RViylb2PfvUc2C6rfbb3EU997
Wyt+9UEJA4To4kYzIEM0HdCMNrLGsLAs1C+DmSRmzKl1xCNTXgYxqfQBYRnbvAamZhf/s691l8nD
pswINCv6vHmfjDpJt5RFQOVcA55uTDkc2wE4xSmthLEvlRvd3uKt7uaGPO84umrHQ7kDaJH0XPpv
6hjqcRsMePXusnaA0x4HOFUVmlm8E65qXT1cKNYiUDTAySLHLSt48rljk0NzdVhDA4TTL4kg1LMB
4YBh+Fih3kg7/plI8GG2BhLSdW8KzBqoE6PMoYeQApHJTEyhNMk8GUAL2VoBNPPCb7erYI3XpqZC
3cW5Rlqk1duQXcjwlvocq+mBBqhDCwQNO1jM9boQLdOERVIEvO/1Rav3weo+oVhzQZsFMNYViyFH
FtUIkwVlSs1tBwCgqtil3Cf+lUg1i3e+V0wv36+6G0TrDXfaia+sIYYnH25wgGEtFotN1URtF0JW
R18Ihoj/gASkhoQ4ZvZz88ioVM+7Od56rpVmxBF1NcN2KxbneeGW1wOXr25zFQpX0lqwQZSc6Mca
7nzTpfDaDy3BgpknnPx+Iib+9CMv0ypcPrYTysD5qa3WSddqv9rKlYnwyy5eQn76ovwDIAmh5y0L
FbCAE/r/MoEYIsW2+NtlP/53LlAUAcjS8BwePVZWBGLl3vDowffG9Ebzp+ZXOAisC/g5kFbXUxF/
ppmHqvVSY3IA59x9rlWn4E4Xbn3oaZLtHenMHW+xsnsljoX3sNoCkTnlNjJEqImLQH3bT+lWqoJC
7hwumqniv0h7uLC2PVi33Al64WbofU9v05cpoRypsKr/kTJBoxP+t8Hdhl9zeoS5pBfJFoq+pNs3
eog/OUV1gEQNTegbKVwx9yxgEZckDMa1ZjCEHCvw/iCtLH1OAChLpbtb0xpk7fygkWDKjQ6Ds6zI
t1gVUHF/c+nNNQAmGC9cncYLyIn87Mh/T1BqTlfCxWmbx73WVmMyT6Id49o7gYHSNoDrlLgpt07v
VDhvVv9rGTzLxQl2wQDVLnxJWFQR16XoUnJjOS3WaR8Ez0Bqla/zbUGK0MXdi9m8REM4IKp7t58Z
LOvKjhPj/Awpfomu4u+4QeJ42KmqSnurnI66mTdOjWBduRczeVVMbvpuX7hcNmvI1KuvG9/v0Tt6
FWBK1xMxLByLLkLJXwFb7k89KWLQB5BOx9YMiKSYHP/sfgRHRV6wzlvxcWhlwIwyicQnXuozpTtb
vF16yrLrl58wN1nsBkUZGFkJBmnKhmLf61Deeik/gXnzT5kfaXEjmXxkVj+bFt95tRmY77jT+7Ed
JuYjbDYY2Chwg+l2f7xb95dvBKiCYak3oMF3p6iBeMJ73Zvi8c+KhpxPcQ9FomZB1mJaAaA9xAnw
k8UQSD1CQwPer7v3jLGrs1/JD5StzC+dJ98PRpRXG3SsihvrrbFQ2ZHnTRtG2YLstXxdLTvQAb7Q
DCX+1NOnkVLq2YoS6ewwNMeQSHvGGAj3h6MxfsHQKUOVGfZX4sbNRCUf3KUEDLVFWhZPFaVzk4rF
+Ltl4+4tfIiHcyRu41OOAQZl1SrNCxSwNWzYaLbEOL2nFMTDwr1PkYq853AbemLsRRVksZOz29Vo
wBmKUIbDffFSgCrwXVjU+nyQPGMewJewyIWvbeusYDoa47V5zJwvWgWIe23Nd0mlpnN7c0wZx6HX
Sk6Yzq3SfMfHL0+1tjm7PnWmcSzGAP6vD5UEaXCkyjUpV7jNVlNwJ+hSE9//S3XSWMw2Qo0PyiwU
15S7LH9P/K9VBFJ8Ne/i1LWa3Fs7vtdr44SplFaZqU61bk65zcI9c3N3cEVn437OAdqclCxbgTjr
rhr3AxoHAwhHlXVW+SDYApjA48M31s+PU/8u3oSHdRA04i68lYOTFCU6KYCP4vmkcAraSCmBq0ph
4eGtmP5ZMwaV+UR0fcyvl/TPDQN7L2V/Xa4JwN2CgrFRv4xwALWbZQdUkMFe6JOjkainTJHICZ0b
rSdkikRbG7efEzdvxBnJuGqmK5MAi1pBzzCAhUUMVMYynkSaO5xyCpEpojS680lgYqjxj6JXzHPr
Vu1TpJHMw28yq0NCkx8/W7r+19qrtiFH94jfnxsu+mK+3vTE7sepjBo+saGSdEH4CDreTjrlCSOP
YVA4T4xTMtTGIGKgUEuT82ypngHA9mlpB72dw6CQkfeWMb/KQh5bYQ/RetAohUi/b4iihnPH32Ob
oLWKfb3gvTcVF+qPDNlFwltCIiE1RmeoqN4rtET1deEV5LcKG6QYBwaJS8Z8mNGUCXjTelNzdIH7
6dEjC/+lYZAw3KNH5Cm+bVklp+2fuNuylvJYKZVsOr5LwhEBJ6zP0M53PZoKH1KHRkT8CWbKr3Z9
F2sBOgF/WoL6M3/fEsSecBjIhWHp9nW5jBwZVdSvyqNpZ0paPDUPgPz8Xo1yw1eb9PZQCL/DynW1
Lxk2/2LWRT5RDmQLWBhOmfNtaLRT8y5kiLiFo1ywRykBGpqWv3byEEwei9uKS6LsEmPdYzsO7r57
hRtkJhLlnba0a3UMewiAHFuiFwX85bGmuGAi+yMHkIDJBr8eyubkpT+Lf5MVr4q0YwuPILejGUpW
fkgOiQm5GEYn9BCrzDPAfCB6FDbsS9+tqZpRDhvB9LGbApMICI9MzaAFcCHC6qO6w7vIdWkTkEmI
zvBNSfDba//RV8vSZ6yy4Xi0uHZLSy1JiHu23gU6O//wyBDhBSqX4yq9lKT96/TpxQDyvzllUkRy
Pu2eTVNfEfTzBOIoujNFCA+yWdjboJmKT8usjXTnajjzbuKKvrci8KS7+tvnis6BBqCQDyN2ZxpZ
reqrRY8zCKsV46PM833IMaRcx2KGeIu9zZUKabTMOdl2CfZiZWOYdw9R/3vNNk9HQaNc+mmiz197
+wf426Rtlx5i35cZzCkayPO12WHn2ek+WsQXJAKPuXhQ9nrwozSnV3waXTBkmpih5mmT89N/MRaL
t75GjGBNbiWOn2x0WKDSvqSk0MpcQDVZ05DdZJC/8l9GJjAIpwjdAFlMAjK2532YWu4nngOB8hJm
Gu44pDkXTapvTZPwAO3R9a0B2wtIUiNsJJPp8tFTnucy6Smjz6K6VQ3aGW6elP36Sqo9PlZ+rXxm
Wja86oHBGpKU2eSppcPtdXIK7+yb+HKzU+nHOOfaB3uPqDll6yXf3oN0KF1MvJX/P+EW9Ir5VbMb
NnzBdWbp5PKQmBM/K/uNspIP0h7Dmbhu0Vij+RGUOunKr1heNNDbdFGic6dUYEAGFz/0W3U7/Ons
JxMvmOwScC1p+u+ctii6O3BOMMr9lK6BoWqveHDwo7RvCxuzjxUa0qUJLG4lG9oDb6z8TvGuZUeS
jbjElQ3NXpNpWHpoPkQV/0xnVzU/iPOoFV59EGiFFKyjUyOlDdxrT9Ha6nhXTB96hFPZ+wdYtHlW
mAPOCs3gbw4UvAaV4OdwEnTS4fyiONCUrtbp8QEqrHk5RO7UEGUNoobZ3vMeDrbQPXtfVRFnkpSq
JyX1sBerXtWi3BmkDQaL3c7vroAHdVc+IK4LxrTQbJNIU0Z9SyhS9cZgiLYrQac9A0/fJbA4CTbz
l14GJ1OqulRszRHB6LrPlf56Ge4QlHtOmn0FIJbsgn66S/k2+pkye6hcvaFoLD6H1Rilf1dLM4S7
gW52EUMc22gHo95INuly/PjCy4G0LjQZebUvsqApHAgIrTMCR5nHNCVg9Bu6SsyG1+zt9v4PMnRV
FVRNKZi8RdEMHeCDOb7BgIEVIKhYPqTnbHNKRwP7w9TaU2W9UYOoqGiDYb32vNh4XbW+3zqgRNsG
8l7re1F2B1u/2plq6NsPMzi1yZgSfwkW15Gq1hrimLRehnTtXoY3noG1FPPMt4o5+xJ6FVI0RjuI
LFmJWLQXGKZx6sKYxyVXLgaNVpIBSIPkag4s/MGyHkoIzzXylUWokMUNrINjZE1ZKqUfJbm58e3h
JvjvDqxj6+3k2VjRcAneuUVvk4QN8+nDvSAbH6nOpiEYkN5oCHnU8eB8TWR8KNcn2dcHBLmwrGeC
7ZQ5NtzLEZEUb4H1jhjaXran71bzlcNZ+6he39OCsZnQ3UmI4K8L6fDZ3JIc7DjWWVboKHg8EE4G
sAG7b7OOuYmLCZ2nGlazl8ND5Vb09SlwTjjrIjwNoYIYGFX3hFVIGfENsuZANbuvLtBplZMa8z7J
YsN5Vih/CNhAFfC6m6FntCyn65DXd97xTTTPlI7eRxtvmm8hKT80m87QgVvoLm5ElwP/6gyy9S6G
pQRzs14N/QPhH/74YTKKDmpvRKGtU0Ilg+G8/MwuiCAM+fI58QgVqYaK9iu4JTkUVizK/vkqgrso
xaqqNKuIqZgq2RX+dzZPm1E416UvwrJyb1sZ3JRs3v98zttOyBVb/J33Vydb4CicHdojfORESKYt
Asbirss/NVhT1AtroL7Xp113PaovLVIvBAV+SXXoviRxbnmU3Ik/QcZG+3G+h0NJFuy9KgYKAAUj
z6FtEg+PhBzddAm8cVi1nWUUf99hvMC4aUH+hdA07s0OaMt2lznEzS4mtdDIYhtdHawTU3ti1TYq
hk1APRqsn7Mr3HmcISWUcNHUy9DefnRVjwWjUeSjGtRcgFr2VP/Nt3sAL3kGfCRmB2jdYxmLti8A
e6ndUhoWjpRu0bIrSVnJU8y6NR9mhrnEaxUjpRjrVqp9UQOBOz5eHrmOWnqQbS+ZjA7NUytLDcOO
Qi5XZDCSCd5jJB8fg6cfEgrnqWHDIX2mIkYVTc4mK9Bm+QvCWKJDTp+JQM0WkhVGvo0+1hv1vrIP
csoqsgYYRas+HhF2TzhgAkyDzOCO6KrZEOpT4Hd7pjYRCbLUBS6ptDcLpTedgdHWTQ2mjHqXrUuF
WBZk5iLKmHwFx1WJRNv5aMyjJNaEwn3qCqUQ4G+7tRG1qjnvpeYRkFhVPNJD6AZWA+6XDRTBQErM
Tpq9avB63QjI63UZzvH/Lj3woNQOVQBN/dwINaek+ExuZI57Dk/9yvtcll+tnuVCsEQ6QvUE43/l
lhn5WOUdAWgl9nXP4MbuxpV//VaTFHAXLQ+2e0gEwTsH5S2qytlMMjIAURtzV+1OElLt3cnzi7Pw
zq6nR5DX9c/SmQauftslJuCXMwqVd9BVhuZgnrO+eEI1tPvyWt7/xNcx5AfAPQrUtESbt2jOt4NM
G8VWv6rbcdyuQd9K3RMIUt8S08n00UC6wHhoC25VmUhFGkKignF4KVFetXcQA/kPHKSdkv6t6Rv9
KKBBCguwPIhrO/SXUyJ+uZwDTynbszIjtInaqiL0tEAabldwS0xz+cE322BalybnlDMrgNJL4/L+
mN4GFC3OILd83BCltGqOLBTRCHdeyh8VLOY9IkW/aiRHkcdnJ0Zfikaddenkyx0V1QeD/LXUwaB8
oGwPaen90RDMGh7/SwV8Q86GxKpIhUj6uPxnYtCUgQJKy6TXmw+WUIoS/KOQZLle4eW9t+Xbj5kp
Mf8A2429SrGs0bnub+oU5DLZtbqd+DmcRc6Ja1lzUnlibOn5M9NJHNU3T90q9K2zEZIVDiWt5oVu
r8WCSFv3RXoe3/5RmcML2Tz7ALq/5wyQlNrOCqDaiZMlUTti3EMDdj02dRU14klK7sXGtazzzS3x
hkSlsA5AEP9dja+GnxLpoufNouIa8ieH8T/PQiTY9yXmH2oEfOPsTy2JxntMvUXqAwvS4rWTreAS
6lqqbjMpekwfL00yNrjUkwOFZCk8PIYSlfa1VkkicIVVT49FwgpYm1HofKld8uzQewCm9gq8ZZ0J
RRwQyWVYzY170MVZbW5tSlL8TKVe9kLUY47GrXK3gBUXYaCzm8pPuWFJQNHvA8nfLQkEWvKECB6x
zLvezzawxa3kVtqj0/biRihAzUXEjvM5N47A9IFzN6I5vdbMl1dwwYLGhx7ede/HLZB6/u8diarU
RVYZDm4m1KaPhArkLmGgwAfts7HN2/qeTc5vBrxnlDrkBZ7Lgqb6+a+PccqOnYpLYs8K/ZsW+oTH
C5OMJGBdPXxpJbYnaZI1j+fFFpRLVbLL+6scU+9xFm7+GvXUZunVW3sR6211oD8QgpfXIDJDlWEP
wJo8GxZgMztgJ3lM6AQnBJX7DYQiLRYDM7qSyL8Ow7BRRxU4vHrqCYbYnYUaI/hv3A0pfUqTL3KO
Cy/aw8ABjml+s7fUQjk+tMm4+09wDrOIxmtkxDurG75k3MxBdxcCvT9QHF42BiJI4H60Jt5Dz9Fv
JiFgN17cwwiaHQjSJ/TqgWuTt4lQBRc0EW8SYb10Pavcg187L1xwsknzgMwjVgIIAAbjPYtc3iqb
R2fSddU9DGd6rt84FtZhsQbNHZPGV6fTi0ks/SS1wPpHv6s+uGqx7GhieqOKNhl8Xt1p5QTVkYFu
CiMZ1Zp70ZFcsRdLgBUFLQkrVPh1aKTVfTwPMEsCn/LgKhzz9A0h7UhaxeZKR4pmQNPlwZ+CrXeB
/PsP6OYqdrkF7bvbAHeMSp7e0jh9U0GlWUnqJrvdMMM4LjZZy6BTDZESPPLFSLvbMWZu4CLS7q2d
4vTDyzM0RY7PYu+HfVAJzdw49NV/XkEUhzHfFItmNRusM5gl4UhP7fDPn9aQzzCiJrPpNmW+4mX2
Pp7zjOk+0p0OpwLMkKSOv1ecBpLiZ2IZ/JlIZzDT/qJbMi4qkBTva2qpbGjno6opVK6TRNesZTR4
hgYOJAhENtzzmjDQea4cPVeXFBkACkmfv/lIzdfh1SOK5WgMqAEyvkVvswWcfbnaf6sIiHtIJQt/
YkOcu65ltuzdmwMARjl9cWOqGAGwzcuxI0cpsUE8bkfWsMv2LEJhH41ZDTlX4XL5EcVYTASkAw5p
BZAPJ+YNtkm3AiHO0c6wCLIX0YQey8oZM9BPJtofy3ugBCROVTPCJfyXkT4iSCJUQN4iajkyW1WT
YSSpy1p79T01SD7RNa5MGzUKfVIrLG8ipEhrYn7caCwZ4PupqMF/CET5Oxk6T/PFb0n/mQGCROJ2
neiVlwe9kbx+4hc7WDaZmNc4erUTtQjnmmET3moedsfItDsZD9PWi5hEaHCFuyI3uPWwK4lR9Ws6
4SiaQpJE+BkERHURazvE2q8sk6NB1+BLRAdST4UApQL2dVMCCl1eNBtELtDthPqwt0IbUufdY3Ov
y4k03MYeAYWUIyxGOzgzjNT/AY7zBtM99zIRvrPCXAHiForGQsv9KbVjXEnURg3KrTd5euoa9r6z
PnrhnBXSawFS1A9eKfWbuieT93RGxnUmtMjMNKh1qWZVsSGGHhVPF3LzMfZhqitv9mH7EG/wl66v
0VSLxu0sF9DyZc4eNizRdy86jMzigT5jCPz+KjJ0Z19GsAEYIqfEEbrSMgXENgifWAWuXgY0v6bE
FJkqqQtQspJuwwKtDL5n2iakcOtPV6vAHth41xhEeIF3e5mXXyORnLW/7rOfn+7LeUBXdwBzgIVe
DvN9gABfHVtwv5qBVzN+iUW3Lwumd9xXdyo9vHbSa6YBXCTkq6P6vECDpeRWNmZRLMcOfciQVja6
G6URBjWLLfC8nOMhlrkhrJBNxfKVZlUB+seQ4mjrddXcdbFWVxzvKtTLYTFfPjYF/VvqAvevKZB/
Jo5w78iGWZF8SYrycu0psQqzNLFXj2XacfUvG4HGoEBIi8Pgqo4NC0fqB37DqsllB6kOYwo67tvc
ingrfMwcAK0+5uY0MeB3hcuars0/3Pmhe1abPeHjn38Q9P1VVehDqhudjp4x2H8nbL/ELmpp07PG
yOCLCc7KmiFy4MPRHzRoteOesadTWXnwKopDkUzzKn+de96d6+ZycTHU6hxjg+fLChpQwmBBldAt
0/TQ1O4NwdXaeU2L8R1wOWw1oqWoJNy9gKztGtrCxCtchLYrlkV0faJ+8n/0a9BvoW3DDm0O3O6J
giB+n9uIOXicnbKdHv6xtP2TreSwiBZd3BJacMWoTgjHQ5ozngBVFGlEI5uRM67ZX7Rhz3ho7B9y
XP3oSlj0LIbrrDy0bU7N/W5mi1JR0bKR93GXAF2hE2Wz13HAtqZQx8yK1QZ6ypLGRUaNKfwoRBCx
0uQ/c3QLH3cBj+4J6l2ndN4+Pu3sZo86/0lmcxbgnFRPasoIBdxdCWVFL/6i+azbdOtdqgniC1h2
vi0TCX31NR0qHjJnH3+W1CAQkbDTlSsLZj6nNjc0kcXY/DsuUytLm8mwSf2MTecxAwn5k6rqzfmz
c2RSRTXC6otTtQ6e/p9n2YlDrAwCJSmBxBspqOYbYMvO0GherOKeu9cso0lKFr4t3nIqzYV7+x8v
X70kaWDcgsezMuT9XJ8dTn67sQ4LC17Szx9jqvkrFnyXpCaAxYJluuWij+Fawsz1ItqaXW7ylW8/
UpQdm/8jLmsObhLyoFjhfstc2puYXLe/167NEEZMkSlVV0iH5+NEJqKc4rUA94YqT3w/ERWYEaZC
RVl+tLqm+G3Yr0fJ0KaWbJjFH7Iz6sUj74aWdbiIFH8cMhW8hj8fYxrTRJPB0w7i+J4tQiYfLQX1
Iq2SzZCmWOUATiD7/5n6Mcuuw63G2tqFZsASqH1oiZK+6oZBrKJzmQTw5hvuek/MOU5R/H6eFU7J
y4RX9UmzgsjqfVoxZi+wO+vyicRJmM/4o7CGZVNcpB6+ccc8zCbBKw6G79qfnXNHJQRjbMWwi2c1
nrIAd+MRLsDE33Wmc1L/3doKM+KbMYBIN9yBwm/XsZVwsEk1QdX/Uan7S+3fQZShK5xpIZ2mKYnd
9uXLpv33kxZaOew88lFtYw/IULKw8w5+YItQIupsrcCuTFphexYaK+SV+MDLahCnbFRk6+ucxW2n
rqPDTFa8iQ/WHPXFhVY8DC3DdRh26dQ61DnNmeBecCLLTKN4jl8uzHg6oLaoPHwJmEt1JdirZXMB
761UVcKjCFlgekcvLtX/CpoPNOJSChvDaPi/Ami0vES2icyW6Oq1dawOBwxgJP21464wTObeViYf
j8HjUyhG81f/f3GzLI+hzahEQromwcXQz/HElzhin/AvSi+XhQy0RMhDUd9F5DND5g4kxY4d9GpK
ucZnMcpWGLTVPVO0ZjDlvjEzTgNmywvzxuQ+HKI5b4gXbsXXmrJt+PcgDAMJBiu2rNxLiEiXEHPF
P/Sfgtrayo4zBsL6L+2H+fIeROiaiewnxfwX+VxgIw+54rHJ1RFhoWrW6OfUlevLOkgF+7FuwshG
3765kyTvvv2+yPjk6kz0ilrDt3FycoulnkMkqR+LFewLXqwuc4CrUrQeuHrVBfb/4b+FX7iAew36
uJbeyJQEI7mv4h8gBY9pmIVKpuqGbZKobkjCfrDAqR6FsqULk2q5VmcLJP6MxJQMgEVson6PXMWX
3HM4ltk0VZMFDsKUAG0Gl5l1uQ79hT0nIzgqGL1lSnJjBtbPsC+/HbdSsLWsHfje9zIF10XVIoml
A0iGIVSKiblncRMHBBRGYwsS/6a2nGs0lJeP48I2K6nBaN+s1Jyxgoaz3hnsQ9fE2U5ypsn/0weZ
KPBpLlElouEJusi1ypGOb5bamRkaZUJl7/KD8NC85OeDLL1pEdubTTeUNdSCshqlYTFtF8hzuhnu
G3rqtdAQlAnc7wqm1dlW7EqRvZXMoiPqmpjR9ONsDqBzx6J4g0j4awq3zNsJhFWBLYjNCdF3Htnj
CNDFgpZcwzb96TTQS2r4z4yewK5G6igMaxI5xHqwvSSI+LcLTnNembIzBiP7Ba7i1O7m/wkun6HJ
6PyJMfZE23Pfvcym6RzNad8yF/EgkNxl3jcery4wKqAg3CQeQHFWgcUGjyBaeMkEjo8Qat7BG5dU
8XGMkFUjZvuE43nWOVZnBfjtvL0Z+QQdchP3oVc40XfmcAQMeeMRC7PYDh/bXX0PuOLnFhPuZnUE
ZluCKA1PeBDmEQGuzWnh3HJFowNb/L87nlPj8x1/pDppSkQMqdgB16y3AxU+nKXlNMXv2MCcG6p0
M82Bds9eba5GKynzBvOcuovmvhSN8Cccu3OXsRBZmwg2P9qXsZo7LSGZ1Oh/YyJALW5l5NokJNpj
9uUBGcbs7v+AqfIqltM4KE0vGz2VU72V5iLfitlgkAhVeVzm+3G3/dFH68IBOiRc+NDf2eWbUebJ
Mb+C+ZdjyrddhCSYBd8ilQHTSX2D0mVjE2TczMLQp+g7yzEr9PSQ5rHS414vuZ/9umfn6FwJd1ZH
p0d6LlrnBQ3lTCocjOFLdEhbGlXifNfYbiy4JeM+LOOXKHRjhNGAca0OzafRiKsBbrKSUWuoYQft
YNspO8fWmWR4gTU18lTAYEIxd8coGPdaknMB8AIB9befoWIUT+vdi1AaCe3U9gLXypWq8DFtO/8U
m1AAR6J7XqvC6qqNFv/lW0Ad+j6rACUB1kyJZGleDhHvVWOBOr0h0uNedqpb4L0lgFSvqgygiJnZ
JHeAKeZPif5vgUVDYfth+vnr+KUizGciO1IzjnXkFcodASqy47PUgVgZz2f8ILeD7jrDWB26TmTp
FTgyU2MCOMpsgcBVeZv6Ujghzv2Ju4b2yv0GSAGYQMTg1MiTW/P3lSPrVOjazM+CgBDI0r+qdEl7
FOPJ85yawBhcQwykBUXNTlEd26HhzOwnVvk03aG9naMCTB+L2eFabXG1Bh0z8AMFyRzPo7tOt8Mv
g96N9ki5S4WcLqnMx9SRq9Jgm0F71RzLo5Aw7TKU7oqDR359UAd+kezIStVnGLkKOoQVrr4QN/f0
dxVIjGjmLRzkdDTyVDwUH1ctEqliy5iWb24lHGhlvohB/Ji7wo7jojf7Y+eBG98oDB5d7F38MfTC
J2O7gtQOztE4azv3UgdJmU+iVDotwuXOckR+7dxD5tU8hYnunuYqH1Hagby25272HOaPYkPd4xHp
BSvRtlaFQG1X4eW4VR8Fv4crtWwuVklcZPWH9FV5vaEyzo3Mp9g412YFBjEL6puEklKCMNuA9OYX
nZHR70uYARl+Qiz0Hf75ucufTo43DmwtTGJuTJdIFs/ayE1HNrqtNTyJpQSRP53HqVUnSu8MZ3/0
rJwRHLvnBs4emQLRb4c6BOImqm9rdZWGiJF80G2TqrfRjOBSXOPszd4TJcizdzNbrnO9exhaGLlg
gmU29UjWkQdGQ2FYCTo1sLEyp0ugupAt7+9sVLMu3y9hpecZq9gvwPFbs4o19LzwCaKwWOrktAdG
uVSkg2bWv2IZLo7DX6GCjhNsrDO6HwyV6YMAlvh8bL17mPxUHuyuNrvf9LPZbqd0dsVv74qgSn0c
SdKRfZpV4jMqRpIO/tQGxncmbCFqphsz+2Pn5N5QBRCiDBHfaF3NyWQ2iCIDfMylComwq1Q7AAr+
fLcntT8LXv0OQAhwmu2evkUEGjtUlsjmmeh8Le0OMqR7+OmM9YT5dBTraVC/YvYwQGz/MS5j+HHm
+BbKX4mJYvc7TGaMwz/s0RQeiIHAt5Q2AFcIlppro73aqHLXjJMoFmvppWVzUTgkSfhvnObFj6eS
JWCn7zNQMLoc10PlGUAqOhtW44ede8byK5o7y6NehS4bziofOfxODDapxrspQVQ8oCrdDWNAX+YK
rT9zFwsu03mFyjygvajeG3jRLEpMtShewnpOpy0JqwndMiF0VFlFhwAwh8BmvivCRGEDoVs0uHwR
Cja14nvLdDlqbMU3j9yRuRqtyGXrPGFjWVJHi4tZ7hqxj3sZCxMqpG2+eU3ipslOHj82hW+KFyMC
MIT8gOkovOo6YednPaGb77JHpcaLNID2c+dt6T7dny5/EOlC27daC6+vJVC0+hrnZtdJnWWbAknC
CUzDLpuok87qg4KyAlSctY8cV25vguRHAhCHeeTeOhltnPcIIBEhpx6/4duQV8PcvrIF4hmp68du
dp9fGhLS7/F8sx2ov43IWKgW4Jcil7quotTskV/3SjXUr7uihgQpMpjGOdSjzGDGee1OA1+U/1FU
sahM6l1Q8aDi/mSIcTJVp6KQ6dd+B3IQGQnipywLp6i0fM7QELinhikLg2tZjhaTV+LBLroTTh+M
sioj4GVJHYxQgf33OWx8AEcQIcxTCE77k1kbCghOb7L9jhShNi91jl8m0n6GZK5TUDNptg3YzwSS
8/y+/FD7W3HBcKCsjVzzZQdy9LpT+ZOV4//baGoyxiE9i6Dzazrlr6kE8XVV/18W2Mcns/CcgVNF
o0skzHq3rVLgcYsmEfpAitwGtJFSPEeDr6oB48tZbn48+EtdhqPTslKHWoVZZvgrPU4qzTE+e3RR
o7esnClRnVj9cDqLnXs4ipjzvgw7Ty21aX3QnhoSDTMeo5WeHYwvMZHL9t7Ipi1h3eF33piFH51k
XerCxotVf+CYYl7BcoMYqPlG8TlDZ38JpObhi/+QZrNTR0x0+4woNmp3NQ+7AZgxKlyzs1M+OOcb
06cXMHS75wEq4Qriy2IfILIrZ44huiq6loqjGCwcl0CMtzVrYrGUjoajCUn1kJFIINaCZcJUauEB
P7MYFthiNdSXjHNDLPoDEjDkuP53jb9fX9T+cPJJ95frXiTJ8pf199aOz1htoQr31d/+QWYSvBcg
VkqRwkKXh2AdojHw1bDz1aU5wAxCl9PQ3H+Cr4uSYc01FBUUYGYw3Gwgg2msCQ+FAxouJ/QBegds
U9018QPsz4FuylHcETyCvpYEDDZid/Vs/U8/mJjtnTuanVGofMhFBp+rEijMIDQs71RhkzqZz2r+
hATQekb6HcTV0R0e3kb+6wEAjBnF+hi9m+uiO36dhulC6o3xLQktQiYiXOtr/bUlBx7qkib/FHRc
7WQg1qhDsJ85/2TViaqsQVHQ4JPlHVhypkiwGSorSUHzYwwsJitt7ZzBogtl8J2sfGgJlF542LOE
jFuxRN8FXiOeM0ex4Hsf2hiSv41qgPtXZ9pr5Q3wqaNiGB2yM3ho686BWQRCYqw2KVmc8IQ3YhHr
rBAvRwjSTNEgxEXLyA8FVzZvdbiDL2Qhm+di7C5+x8iQ1x0EVzkEKMFLHL5U/wMPCjgBI12Ak4dS
3ySSfwEitptvk0Yrvl9g9CPntjuR/DPN4ov6z5lrnHdaZNwxFRqOErzFPgM69jSA5+B1SEfek3T1
MUE31xP1KjX8jz+0l4fiSkwKkyTUUftpnLO64T81zaal/qf01T5gn+Ifc0Ve/N2ERZsmE0DbdDI8
masH/gvRh7VOO3/fymyCiOpLeK8adaEUj1NiHMLStZ+JZDm8QHjelsAJQRvGcm86nBeSrRy/AiUi
ti1TLIIlmV62IyRDmGnqE8aalCFQN6TskOxyTgPXZx2oQjs5xKeJ6XiES9PLtP265u3XjulcBcPo
fCXB8x/iayzVGhmyD+KKRFavAs49gbDGvKZFaQfK2dAGhZf+kDKPyPWd/x0didE6uNh8+boiO63L
YkFwOmeLw7VFLeKcj/eB8ciV1OFTGmygJuSrR3kUmlX3ICYziJ9g4Jb38EKZUXSxodVa8aBqDrXa
AxPejATCpTBqqOyympe37qDP1v11XmXzl+xmVmI3YNkXE4hZdxzMxzTZgf7PFOBRlDU+Tm7SWDXn
0ZETr8w98ltMGIluWLTEHvtD/xuPlby400nutCgcEZAlHcIvuBQfGCAOOgkJK4O4l36Hfu7JUAmM
DHaIJTCVIk611Yfc6Qpd6UCLUtCtBeiMD11z31JSWxWhRMtxQ+SnQYL+yEOo3BDLjkxJRsqJpvyC
tAktkWKpl64W5uIjxkM+Z2O8ooZlzmBaGf6Dt2uAL09YaI3ZGvUegWUQxhC4tsKSI4xzlVgOdnNT
YtkvT8Zh1OPwmxZoStXG9nzF674H0ICV4D5eKuo4vMW5nw1dXKLZ7zbh7YRe5Gt+oYyTDta4y5PD
GxXM+C/HDQHgDNPDNWSrXYKnTxG4al8ovjQ3BpQvG4KxrpX2v1BNrnyvRJ9XpBuRwCXW3LP/X8dq
4vvrLeyrETyzppjIjtmNUL0PuEi/4P/GiDEIInv8r4ehq/hNPZ0jn+VCOoMuPAeJ4Ccs8o4pC3Pr
XfXy2Uww7bM1anPA2yBdhjTGGynvNWo5XHyF24lwVqf+VlhDbMJGaQ8+bM30AJF66LMM9UN5GV14
2g0UAWpwOr6zmDcEg6QIOfY2BHkew+fKyAtuk2Jw/qP8uTFfnClCwNOKZAGlCD/pTwoirpQzlCbH
QyZJPkaZpUDjcvQN2hKM77c5scGJDKR+VWgCQ2gEq0rol1XsbWhMbRC/1wrBuBq89TUH0+kLDg2a
cSFfYM6rbBSx/FjvwL002zFrb0d8HIF8qcE6kEqZJTHVrAAnJmi277yH85bSKdmkRWa9ItybjQ6N
2FQU+et8M+MGystVYdzvB0JlX+JqndnmO5AWddEFglqXY3WeVMWXL688AFL3/iDU0o+fMSn7gDI8
8ObNhzTyMeHvc4bQRgoYvMAsR1NY7D9IclOx0Xu/KFfUaWxCoNaS11UulYlZCN4QAB6iRJvGKPkq
V4vxhhJFTzf+2laYRBW+9YVvDqJYYI1V7olmygcASrhdKMVAdvdTTXjUYoG5fxJa1kscoe+L5k/h
8LsTbksILZ0mDJBLhjndWlcktSv7kdFq0hC9B+iv8qaNTs+lBoWJvU/sHlaOJTPbRIbEF1nEZePV
tFtbyChTJM14tbn8DqIoWKeFlFbNcvvvG7h7o5YLAOQCuiqTlaNWOyJA1WmWYMJIdRko+CQQnGro
xBtzakUceS3D0mubefu/qEo0O6Ib+z0fEbqT+rk+YzQB7lJmGo0QyY6w8OQBtzsdYxywBcBFSr38
LbdmWR/nldi+CSIVc5FHksS6TElNy5348S68FfS2j6t34FvNZI78EHWH9Gux+vfHFv1Uy0qMM1UG
OFujI7wqIXCHT6lbJzb27IWouvlYjEQXnt0EPyuo2uR+/jzvJb3ST6HVDJBStcg8tSRFpWwY/Noh
pHQmvPXJVfzMO1ZgsCOEg6Dl3vuvNpY/KglJI9FHjS0CeU1/N5f13GZyTbteTe4BbD5nNuQg+e37
ny9J3LsXol/cKGU4HN/M4hFeJagE0QIzLamUPf/oNZ/2mcfDps70kWGPK47OX097bQJsaEkRzTal
KmHBHXpZxinb+CGshf9w+7liqyHovR4fH8/oeC7z2y8wSN6ZNVwt0K7DN5dhEu1t6zyRJQovU37O
9R0lb1xvNyfpnwgHTBrBo+SlJDEbafXTS36890Jd3hOxBmHFQaRCcLCtT5djlkLvOt/sIS1Xkf95
v2aq0BtdiBYiA5cPpae4mDqhnbJRWZQ6xrmPfqqB6T8WqzuhvTtPCsoU6HZ9wgd1PudkCIZxfnFp
7EVKf6XYq1QRZoJABnmGFKIMEpAZQYCDFMiUPmoFzhPs5LhCbQWPXsFIWRgSUATWHw7Y0+qZPxBl
OS0fAFQB/DhTtAiYGwS4Jizgswd5clrCAPJw6DWyuDqjcaK4y06wvjrPOy5uVWKjRJHmDKYp/RKq
CQR78Tv6OuAsw+Dbiv8UPcq+GtKVSW4+ImRapmG5ilJPIouAOmRBzk/qDcZwQ8QPG+zBAIwabPTJ
v+wpAprSR9gX0MNgrUT1JpO3KnsLuTWe9cMkQ3hMQXbNCUcTzn77ZRRrOiGbRcx6HvxnWEwhossJ
xB6I3E7LxIoV9VhmfJBtzIIBIwokXSnlJKf9Zfr7ySp+5aC3ydHWAzZvX0Kr66jFAYDxmsTtr8g2
YCN0/catjFbQrzMW/F2gPozZ94GY0879uSV4UZUo0utnyK2UBSVtK5zdSlfhHaYUzmVoQm6gPlW6
+03mQAi9JHfo3hvz4dzGvLtYLd1J3kdOregnKRFRzIjV7mqjVNjIOvrVVUFL/TtEiidryHFvKr/d
9f0ZL3g/i8flv8J2dEa+jc5ww0e6tH83bDfX9hjgX0CkJd8DY/jy93uJpa0Q6Aftcx8LKQ/AhelS
HYdOa2rUsUkoMiMJYhFXCORchlu1Kxc1LW+iPe/4+8oQCeITMSB9nT11g0Lz9px3oghm2CkxoWxz
f4/ful09FyYSgY6Z0mUSUXBddj30k07H+3MiElFOmf8NcIuPqhEpBipM8sRiENZoaWh0vxSz2qXW
Xcmku6huojcvnd/KgVHTTL9IOzgllThXxgFWQ6eMpRIBGjVbeMF9iybZp4NyCulTYskWfgUv3vxN
OMxkLoHzksRiHQE/3/ximG1bB5tc0+dg0JULl2YWM7gcZudGKen5h5+nuVO+9QLBTGx+q/JkLmsm
UiV5/tThR8xsEqMfVcotqPQwENCVaMfOWJhCKHOSCZG3O+5nwANnByUG37VZIgSfZ2UNGqm3JnY4
8N+KQyrFUut3hyUfOpyySZGmXIPcvVuFPY0zTZOKE8+7GAKkJGdw0VyeJBsHjk/CqTCCsZZogqqF
YcFhN2+SScRXmup4C0ldm5rUpXaNJlesNhmQIsnLoqnjwY5sJ49alZNH8pzbXPWaslj80P9jkeE+
PauQfxQKnAoeGIQPT5nCqfV7cU1cXeyzLYaVx7pLfCGnWxaj8D4ZbDJRer/n5cCp7c6g7xuw+l1Z
n6Zb7MQVa73KpCmsQGPUqx0jZodyOxplSIhxQt0msT0EQ/SBYLKWQ0r/hb31gRKpeUafe7LTKP54
qntnVkjgLccK4tzna0UXBVNHvvcInRaV/CxDRBVtMdDzLHVfnosKzT2CfKwT9WRGEQ5FxfSsApsO
RKRGc8zedtfVPH7/uV9nBfIkezkUHjml1JJSFyqsRzAte7SIZ/6tXV105Fwn/xeHFaC08PBk5thC
Yr6nXX/AiR0zNGLP+FD8aD3F61BfLnl/nQjlsDoFcaZjjM6x3spxKxfBtliEAMI45LLBD83pgUuQ
DHRDigeXMyUC78rRwIRAMIqdgTsaDO47hQ2eJV2VsORRMJGlfYfFsQb1ty0G9hpnc9MCLgGXl3YE
SM+0xmqrvPtP8meed5rlc1gQBaayq8vQxF0+pAFW2LHIoRZmz6ESrDQFbN1VlTUvWtSU+05Gnzqd
tGYFvboaKbctuAs8fWPvGoRRJ4TgkB9lp1pt2kS2zjZycvsgI+fve7h4lFuG2O+k6MX6k8rdiVYy
S1Dhdqra+PjSYiEZcvRkBL2nicx48gVR55sZuoVgV8yEM+XeLCXVfASEo3NLraTpPpaOuUUI7JLa
zFvxEsY7/JQRriPCJq8j9B+nheMfPG4sXWc83LPhj9hHZhuTC1soihyb/7s/Kfg/AoJ8g+N+G79j
WyZL3Y/uCTMjqn3EMUw8pV0IaaFcnEhRZL4K25/UPOIIsl/HhGi+UC7ebQAlcmHPrBJsFhqlsUn2
W3n5tic75lrU74x3BWBy9F/OLoUUEqmg21b/lG9b+hwHORAViyB/7+cAVeP4V3dqkeaHDGN6xfI6
mdqcGVbEZMp2S0SuT8CwO7+i87cAUlTfbEEtsF0OZOQhRkupg2dRPOhoglDO1T/lFtUe4/3nAu+s
xav9lMfDjqTuU2+iXESTl3do6Q7+ylq4sQSNIdQ5PWZHSTQmTtqk5cEWvhMDcmJIcYyBid4XhHn0
usQ++hvM+PQVSwxbpBt0v51v1lQgMI8TOIOOcJI6oD5lR10UNKU1NNuKWpxLilK9uZnpVX98pbxc
W3NahPcv5jQU/5CGyvfJtDeLMhhDVB/sIpxHz/IXWjecw2gbs9ZPOMdpd08D8LZfDYV3KSh3tb+H
ZIupl80ddurGWnmcwON/eKeYlR2Wj01WYNoQsaNYhAugf9yl3lRnqxSftOEQ8px+ti9ZpF1ivtgg
pcGU+KOkm2w+/xu0vrbGw1GkfYlL4lD4TwddpthAz+pWnRzjzcYuWX/8eUliO6F/ylEyhUpULWZ+
0YACWidaw/CYt5QzUxj2AlAuRVXAQzBJAEGoMRSZ62EAiNGE6HioJrWoFGfayHCtbawXTSJQerib
5x0//NHdgZ+htgV5IEs6mM8vEpsRx8Y3ZCUn8FPOAwzjwr0d2vW3sZXOEWn+ey2g6WFoFXEm8/u1
acCHncmWGfoYySeV/2SMIQPgmmjQEcPZSF9dL8JQPVnii5Vp57x5jFALDKsu93BVgTUKm7OaTjYg
YVeXeT+LwqfDcS+oWkWwdDttsReL5RiFYHkzraTH2zYwdqsNQc3vf0dIW1iMe47kAYbKmQN/I6SY
meu3UvOzX7+Gzd583f9mzGTnGZs9ymEXuQ2ru/vOig2/B7TYdAzwhZMkiCpHal4wwvah3EYIK2aY
e7V1ezFaWZHeoaOzSyNscRyOBGCQ9QMGVTRkLcRyWb0uGGOgif5DN+720+SrQEraUSJFFcdd9UEz
qFF9zxUA5rdjAFQd89mmufVrz4wbyBq2QwY5+VU4c0dh3daSPixZdUtVmmbKXVTG0/Qostnyzu0J
ZGEbSZLL6ut5m7Wn3bnvmzeUt045BghjxID1WcZS+uVOBJiioZUElu/Wv1nA80cRQr+0ukuUmTOX
t5rejHDhDUhCTAsyaAZrJyz7gVCmz9u0JtBek0jwMSJI5fdyL6NVxqWbvaKWDurKgX7bM/Diy2BN
939eTI9wvyTVWv5/z5PpO2z70JglwoPXiGn0I09YPVL6gRA0eTp9gd2BN6zCVTijJcd5zr9g4JTR
U65B4O0M5HjOAqR7SF2RYQAVmZWlNEOXgz3P4EYqYRegtn7uc1beaP1lPWsQTYDjh+LOgt4BOI08
z4aFDTQLRvmPok1zVCiFYTw3pSjraxk3vJ3C9JEAdmEkHPC9roho4v4LBR2DeneeF/zEAy9D8TUG
1AZ1tntKU3ViwAdUQANqAKV6Cc97sdvXVzEUCurf+T1klH5YbHw/4Euj5fbFol1wzj9kMoRby5U/
XotPuJUMbd5jKQ7fCr2+xzPhAjnBfc2dslHZXt1112E13/BjGEKqKzAkhCqgN9JDfOzsezeiiH4E
6OPpqFZC222IYjo3SKvLZ6TLl/S2Qxy049RYzOkmoYjT3mlY4Nuva9MrGvgHvncjuyZ++ALTxrQk
grnugXlhg2EKvgvOvpcGiRlTM8f5Vl4aHHyMUDYclk4eRRHcK6Z5kfywBvSwIgLKuETZ3vIxS7u5
T14SdSii6f0fR6r7mOiYe7gK/Lq4EMn5t3ushSnRwxpYYzt78TDwzbSnjGlKGxQEbkxvf/rlk0TS
rLBZ4Ex50O433H8JFbftjq6Cyu04U+pbfcVsOkWyHsKKxgvZP7plk7birSO0/tQScKEJp/YDyLgb
QB9j0chlHiu1ZfScVKHTR+KEUs50fMVZyTzDAbvqNT7zi69m8oYI66hxrAsAdf4lVR3btV3GMl7x
fyDXuIaeMKlWgrFXuBILuuysukGx1ficUnfpzLRd6xdBis1MyRZXr7MZ6np8tagdCKFCFRguakyd
ZVtkf1NpSTI9RfPo3SlBfp1k2FT/JUNQLsW7OF2PPCx0q4YMMjcYg/c/Yeg9cHvNlRKIqLdSHBEy
BkCcHABkdYNCUs1z81847Dp0AFJOnou+eSqQCijKiJ2WAGZeT18Nz9urVnSiaIBFTz0+Fq2YmvLA
wwnKtR3HjywG09Fp/lsfAMs8BwrZbz/nzt32jzIOEkAweUCs+5pHT010U6omrpw9rQCoujsv+Cba
epiirsVsPxV0H0O1XS/hrsAu6ReVDRO2AyfDwbgTCPWjmj2MQYFaZnLdKjMYDGhD0/VrA8R2spdS
SW/V9M8xglTdbitqXkMM5BhaC28w+UPn4QbEdeGar/qDWZpxHlk9PzTpAk2fdB8mQ3rmV8tL8yZy
IcPPvj55n6nvbdvsHBI6v6WmOKDidIqcq8nVXWTOOBH9BSLFl45/KtneiVX3/jeAVpHfY1ec94WD
YOhfsLD/qapTSz9Ltk0wVR+AQ8qoCorpPLbJxyveLTM7NpVsFzkbz/OJXCezOrd0Y+sxezn1d2jU
NmYnY8WgSQAogJwu+nBmJEZDjvHZ58Xtx584Ro4ZsWlQlS5Wn28x1Q4KtnXzhZVmvQvIUUDnN678
7vJT9NkG9FK9BWR0gPf+ldHGXjSdpVoxDw7LSdUkNDimdBYpZ3fCV4cFLEuc9gQS1PGGeUW+uOZQ
/c/D3sNcKpHdy6sB41qf0fOQflS8dkK84+CX5/YXr4//NBBDI63XWUPStLsh6uXmOjvnmySTEvLH
xK7RnekYYwM9PZoJeI/dTj063hy1nVtfvlol6bsl1pQzO+KwJeuDmGRrfsBHTh4BZ/JSOk5bm17y
xFRjyqJwsqsY+dDqrBSCp3n9jeA+xHk1tRzvKWXlmYnrEv9nHl8llXX4g9v8LK1s4dh0VDAlK9sN
HF7fM8FaoUKGVCzmjvFZeesUJWYECSmmTU035wQq8kKL1VFblUa/5dDHAc1R/57DAcg06tkPuN/l
1cg9vHcnYwAhpNGp0lhrHzBcSVks0IcRD1IhObHalGkiNhYDRou4VT+TlePvUfNSqlYRMBsLvLoq
OkjyQlNPwvy9UePnM2/AkOqvQJrhP69dKxiUlWEzdi/RCRPBCvGdfu+lxJfpss9Ibs0sTsMMGycf
RAvv3+MNBCcR/QORidlD/UlC5xnNJtm6Oe6Nuo08m2qwQGpqD2nBu/yOZohrsoJ9i7/ZHJcgSogM
MBAxlPMm5pRxP5AnLT0zGOp9OQ7HqKIQhX8N/3xR4fNOLlCKhN+ZD9NJAr5SnHg+fTorOwLzkVky
hpMpFM727iULTUBZxXFbN9EGp7ciVKr3obCcGgKtWlQZGrvNOy0xBevYJprX35MlTip6Gjlj0mNK
L2vxF0xYt5HZS7mxyeeUoz72X2+PV5204nH6WZgEfdIY+f0NEz6wSspLndp7Q+Ic+QQBgBYXj1rn
SaGiGzmJQr6Z3x+yD5aSL6YyBd2/3W7uxvpKYWTNopbHms+i68aoZRrqLmXYkPdGXu9J2mmFMhxa
6mEHvP315GMf9VNfW4eJgXNLGu+P6FrrGR93rRkUasWD4C7TfqB26n1cMm76nI/7MGn8sFT3DgHO
pMK9r8yGePeWRnpqu7ha23Nj85LFOgd6uOjoFtjUjI59FCDr2Oh07xFw1INEGza2xU9YYijcDkpx
U6tUE/NRmQRpJ1w0KeWL7GW9eb12tzxHWLuAgzL+yPJS5fg7h577kqjkE/PPASZ5lO7yvZzeU6ai
N+HktNgsy9VtQmyFOvzxudEnKNPl4lwAibTMVYUym+4JhTqFZMlBINfH+heBDiReTlwps66hD2rp
uSZLIhKnNkINuX5vrTlZWHGt+nLRZeEr/MeH9JlHVF6LvW4RETaQlKA4yUGhL269z+aaWN4a20Al
bJkAZ38X56142kN/ohqDfiqjYPHXhA0ecoWNPPTRMXIyTNv2MT5a8/MjiQoknxIXWC9ndmh0UBdu
FMnFBBdry5gXZfnw67hXOrfOIbwAj0KD3dM4nwtCzhONXgJWj8f0sh8dnY4kk8kkBmJeFdXNMS92
nXFO3l1S7TU12xiRzyuZVD11nTooJQUtombAhTdDqYI9zLynkO1lkwzhQjHYCkWuVpfJiZgM+2tw
44sPa+uOCifNZd5hi6IvDOkDxvLQcpecp6Vy3KTZlSSo8FBfacfiBCrvFaFjaj1d6i42ql6SuTqS
cOSFxF1t/x0g25eA+7ipJYR+LiIxKPOrxm6SQoDz7wPLLl2H6F5rUbh8yV/I6BtIOuBCHpCSt5x2
WUpAO+TDL5QyhK18Qw1JzzHSxZayXzjPxPxkD1abzIorOTAzOi0YvOs2B3+xlOKg09YZZV95bckd
rMSAaYH79jNPA4VbpaIb9Jfaz8VqRVhB9/F6ynFVNTjUqwucDYm8k4p6c9sg9QLZu40GpcIt1yV8
wt2QtEWG95vpjcs3wTqGn7BV8rdBX7PtPwoms7A+g7lwrw6deO7HtIQKvewrqZIAVkvEY6q0gtC0
HFuZfBO5p7EonSOSKI/XQibmMIJ6ECKRWcgYh5l2L6LLMGNqZf9n1EHeFKFek3Zn8LIDAD5td6m+
M8Vt1xaUqvUU/uyT4LKdttwdeZd6pgwKR5GxRvAMAToznjauRWGsSv7lVqSDEBmXol4Etj5hKtDh
KJZobY0Qb4n821WsTHYgvYsEmBB2rkydF6D+oiC1ZLnt4Gs101t0U0s+I1WCnmIztt/2nSSrcEqw
RJWDINN8axCc9HkFqnoPhJQTTjX8wqUxF5BliT9OHJsXOu5qWTEOvMwi/Y2ZQwWYVFeCkJ+a3MEe
kPI3VGCLprbn05Mh+vLMv6lh9iArLt7Ky0WZ+YrGhYxe5MK1x1HpAlWBsPiEVKUZsxPSjgdo147a
rNVIMzqIPKynIoaE+pJMp4MCXo924K9ZLYnlTM/HJEJpvFWEl0MFlYJHCrpQzm9WOl6ANuSnKaB4
hLW+tgeNh82/pRSOUJoM07rN42fJ/XtKii/SQO1/zb9UtanCq+SpVUOKeomb3xLp6uieEa0c7Sib
jiia14ElCM6PBlEI3skzcq1kkXkQSqmUKiCaBtrWKk7lqY9GV37UokTzDnIjU8x0smyKgUM0TDaa
YBhXEHAOTRew14cK1u0cU31p9LkSkgmzhy+m6HY8BLXQ51uaMl5ohijAAhxZKfJIhnNxtOVdPDhd
IC22d91LvrScyBhGRSqk6RsL/l0XbXm5yzz80eTf9bTjQPVEAvWHxqnOlaXqgV1DPRPqlMDQsJvA
1SNkZVnwGfUR0LSaiWcH+uJxUtsApm99767dCxjFqnAz7Mw8hXlJ97VPB7b7lvIEbX4ctVhk6MdR
qinDQAOXOq41ujCRxbOsDN15QDAER7ySc5lv6IKD9yXn1KGDnDZJmZDR4XJA023S5OlHNnNz1L+w
+puDKetLgz6sHoy28YOUMnYhso0ZaAXTt2f6YGLxWStosH+Vhfg62HUgy3XpbgTg3XF+07trWod9
CZceaiwFEKFlfv2P4n7n+ks2s0OVSF9nVrZtbEGvqq3uoxeAZRVtLsvD+gNOipaYRHEEcHHt1ZP8
5DHnRxMRdHcUula/yKDnwT4TseHhYPgSe0wtrei/Jsb8u+W7AH02WSb7dk6fO0TYkxYMcC05bnXG
uRGdoXWCn1WrWMuzfJgxjQaZADOxDt6xM87hAoLuzf1q3PBIXSO83qWYrMZQlKDtluaWax8eghQ5
VuoGtcgYUd31Un3mQcy0695bkAokCbTh7NhhSyHpjp9stxLrfGP015Ke3YkV8xQ3R+UyO++0aaA/
guRbf+8pT3buo5arV1DQaHtVdTVHmJ6en3YH4cXoPnO/pfoMDqFePRcIC78pYlr4GFPjnLBuFCIt
TbypQC31396j1w+SKVex+GsJRtD5xx5jWJKRxuGjeTrMRbziJY1s0gAjNbXIOQ5mRIZsXgkEzQ3s
s51XJg+c1dGSMEpxB354aQObgDvvZQn/AhAgXR9M6r0jtUGmtxyxRya/WXV142yMXeuxwyL5Ah4v
bulcGLOIGT1+1iKGQC17P8/nd/1qCnkFTWiVfXFN8TOFL83kObBqIs2tSDOpCIFcZ0OKtTa0c03r
TED6Pns/Pxtcz273QWMeU65tFOMA7Ous/lGOXbrNqI3N7MZx0qyfajuFz7TZZGswcrPERIb1W2HV
Lc7uye4kcCF2aftfXajPpL6NUEsFIiB/OkTtBYo/RzIBXx2D7BbVP7nCZuRQVd7QVB1Sn1mKTp0p
bYjwWv2sum9QGVRj7IvmOU9wArP/7FL+6jJyFvWcT+pf0u5fjtmTjPR2w5qr0yJPGqBDQD+0ugRD
23ez6M+ZpilRsOIe3lNj5vGV30LJNlJpfswsqTrDR+ENHjq9VCsCztApbstV6mXVCZdF1upaQsNt
g3fM14hvkoWyjTafNZhDqWMo+iWDvmko7QUJHXL2pOduThZxfjKwE36L6B1ZiAMOrOMtvXw746BL
KjHQ2IktYTDDix9NS2nXRYULjCzTGgpFFxk72XC5l8eFBfrcrwq6bArSTgtNPxQ+01XqQKmLxIfb
hadEflAyp9/nDJL2AbfoqRojvvnXYuUdSDaM1DEoRzfnmMl8FtkPByZuOyR6NZzcfKGu5mjf8xtA
40OiAjF9/WQ/ZwxRh1fQbGEPjbeGTsvrDmv4gge74A7up7hc2eEG1idpdwe60MmV8O5MIcrcsIXC
wFsI7sBz9eATjm5EtzgmxCPYghtoXjZrLCy0La+EU/d8EqXA1jmQ4IJwBC3ZjI3jIc42UOZCey4E
5Vh4pQctop/H7OGvzsWGDT0jzsvDnw+QOZghkCdMrsOa+qg/5ZMKHzgXxwksAihRiMrCli/p+eyC
hhih6a2YufqA5+V/nC3gE8PwoPrtdki3wu8ouOw0CsiTg1W75a11SH6wt/YhigdsyOTBaurmGMKg
UN3zZ34q83GL3QP0bwl2AezjYyZujY8vhZtmco3x0JHAaElEt9tXEmReJT8t4y+/C8wGh2BWh6Es
FKF18o8dfPvEAepQN7WprZVJyAKyAA/qnOTbGzBdjeAtBCGRz7O7mCFmoXoK87L/My2z29Mmg9BP
6NWLnrVhwELJJPRNrDHxCSYE03eizaBXOXA5Rvq8Njy2uRNcKDzJkn454H5gr7o43w7d7kT0DV7E
i1RkXC8gdWKtqXwyoDt/V/w10kMHLHr5dcRqdm+8jhMU02QX/AnQGmT2SJY5pwxBDcC+qB4zsklJ
d/XUECL1MN91K3nClE+hwOjjPBrKb8CGhUeEs7sjaizlExLyefIIxpD/BazeDv+rCoc2u95P3GWB
+DyYy1NrnGHGt4eIPFGtKeQUy0LpKXI7QavqK/mUHtrUbmhXN6uPjeWd+uyBT0Ba7Hz9JYRviygR
1DLFadbrPutZ/Q9YJUxeKn0HKNvGnudDtxtLJR0yoonXyN4x1Po3apXxSDDfPzS6161i56yjWKqV
VTmDnix3H3GU+89O2cLiJD8sN4pazsi/GGG+7zUnrTD4stvf+C8Qkofi/iXF5e8OySYzVilfhoMW
KAYDrt6gU2XBMTHKgO7E1nI9vEKdIxawp8Smq5d+QebHcL6CUoYM3t0HQlkFvm/mpoKV0VP+QwM6
2Wxs7qosqMGDSjciREafFdpOHN+C4Ut1EwZlLcpVM5LDd+kVf1FdvtS4VnM9lIsMmZtZEPws3+JJ
R2SrHYE6Nbt7EI7yBC1dOuI9QtDRffA+7/7ez6E7u8F4z+zWAujsXfJePmVMtQWviUDWS42Cuo4g
MhQLzZLcP6uL5IDbxxE/inDthvWmn9OpxK/Mgja9iTDUtcdSUO53q41EP0vYE3xEaVmz71GplCeS
n/nutz7Uw9Kz5PM6OSx604euWkq9bNZ0DlaxfUS8Aivv959tfzTXrbAu7HuNfNGgGQXZHDo5M7rt
sq5EZ7IjFGq5/wBrhLRdeY0haqzRYImo9rLh8wXXLfGhzB8dOwZg7g/ww6y3moso6ICMVG3uhoHe
efwyMHP+214rv6aHdjEWnRaA2IcVVvHz6yoHvPuDZVtrvCyrS3MCZeTlnDVDQmnr+s122FzjcdBi
GhW0RFShVM6jxIeAXfZWaYrNf+Mqme/YooMyOIhajiWcvyVRDp534DbXPUJkaXqAwTFLVp0hy/z9
7lnGremZaPJYiHFC7hUfDE/5PyNPS4ZS/E54gsj5XFbQ17rKwg/ABSzAncCnPIzgvdGENXEq7mWM
1/at2OhennxEg4P5CJ9XEG83z7H5zdX0FQixlwplLWceI9hPm4XD43hb1qRHycw9MoezajpIenLu
vQHH3NHDiJAvCeWpuwZZUWLqa8cBY+YaazO8V3TKr60bAJChrJ2qbhoGefBKUeB7x+QxR3MaRxcq
AV1ujdeD15KgnMxhmxhmBdOkucF86bweUEEIbtbj/bHYs+ebRohqjwsXW5KGyB6PxBNIPiVwigF8
ibWoyyW8VNoDPptLJxbcS9sytcToS6RHel7qUur9eYFsQbQLneHZA7ccYtdXHOhVEEC0fm+2bihc
XeWwu7+Y/0pT3OjUM1BYshEsO6VbXxpkCr6qNYnYdbyaFk8MGyP5ZZFbZW9Dwh1ZuIl+hMB4xIrP
me44TdfZ/tD8aKeHDFrSTRZngbNVpRTN3lKk1PzQYPePaGsG4Uj5pHiKiEDWAhz8P7P6psmfmx0h
D+IKwnSvW2dQQA1tBHeCPo31X4AYRmPygTaMBx144SjD2FVhRYpnjKfGBkwV8qW4OX7WComNCb00
LmMuIkkT+auRfBjiTfT7plXTPtmmE6jj1GBxMKBCtACTtdmdfj0e9Dx0KJd933sAe5xsTaSlDoMU
AKtSqRHPzhrdwsDqZrtH5+bgvL3IQi2m6ODjSTO02iaRpSC4Z82TSoycV+khYrAqKq6hbk8GQR27
320L1kQDvMIKDa8VHHV6t0pDalflibFJtFcJdHPj+ceNBr7yxxtYySRQRmjg/a1KVOGXy7f4ORYq
jPIeVIV1hnJPiJhpAjrP1d/m9zEhGBrPxT+73QypU8AeCRNzetDAqdU2zOVBxfmkgdZXz87N1VgC
yZzaHAU6sjeoDjjc0+BSXMhpOX6aJJPHjKmDYpwPyAus6Sw3VQ9UugM9fKqSPx5qMem+wRqkWV8k
+X4u0aIVMUvw3pW9J5VAYzLaeEYbsJd5h/cEIBYcLUlh+kKZVBEZU7VvDi9gsFjBuQohKr7MxYqF
pD68b8H7sG7EP1JI0516ukc58fTWfHrbNa5F+2by582S6Fa//xV60S1GzsoA3Ndqd9qVKGStemaV
7dzwaz9KaNFMNoRgvc0q90DmP2uPpZ26et0WLCCEoF9kQK57M34VRZ1jft7QKWQ+WZI38Rkh9185
1sh4iWHWi3xLTzCVUpmDwJdCzrQ/Ng276KtQx2CmDc13mB3OtU8n3g0IjXeWr5JVW6g4OjfY3/db
vdvtKNuzLhTC/sWSy8v61O9vbPSpQT/9Y9Ecbn9arF6mYczBI9TndHtJxUyHPcIW/8vij71LOFHk
5S75klhMVs9C5MyV1V173imeR3R3gHJZziog1owZQdYixWLjptguh9eC3ydg1Fj01lhIpcI8nZV7
9s9nBW7ci9Fkdy4LNAJ989CUPiRwQzHM2IfBNsXmANRDZvDZOe/+/iz8lsMdnMb4bTRLJ5akuT/Z
LJmSTukcKHhzU0zHPEZXcR23olbcf7G+VxDc6YIdxMn5g94mbldZsXvMfFhc/95zKjq0KIdffT/z
zcWF+bZoQ/dB4mTsLpHUOSkG/UHao8Yz2jstA4JRq+n4kqQkNZFYx/ndeazcFN1JE6S259Ag0rO9
fndTlbktGrNnLlRScvbDZruAzLO+3d0uh5AEPnTQiOoBxZIHjz4biAK/h4m2iDzBpwD+tG4987xH
7qCHjlc/+n8En95kXJQALiMszhCksOZwc2BC0TWBeZXcfyIrg4v5FfdtfEHoOvNQq9K61ciUWEOG
MGooUcLIWKOfSc5SYhEof8GBcODVywrNMXojOXPXl9mW5DDec4Bj909KwzfcWpSb1GF9Ox5FAti4
mm5pC3t/K4RwVkYFppgS5ODQoGs5tInqU0tyNtO8oJ/JMZVlW2+3aJd68j4Co05a30XoTt6/ofrA
3EQKbIUNo/RjKMZ5gVeIE2XxELMRZMhGBASM0GOnSFHsF5iEF/pZJsGBoNNc5T8oi4O9bpCLk1p6
1InNnWT06lCBHLkHr7ACKjxOhRdvK8wDWJHjJmdz+C29RrdUdPU/dwl958LsoT7YUPXHl80DHvL6
MoaCvSPtcmBxs2T+oI827GgkOR2yU2wgtdod7Mlba7p4Xcqbj+zVyPG51vrklvHB6dtgvwY4NFV+
r9DwBpoEXFQ6c472x1oSf5ejq5xI3cf4YzYawg+hDs+rDwdkkUU4BznRzEvxatQjk4tNYy/BYNNs
cpgN2gdw5JnZZLWnPLSN8IcYHZ0l00wQbzzlqbJYRPNWb4yTTLpvfyORx7fxOhbRBzBmE8tiSvtj
aeqtUuoPfc6Da3n//ElniLryP4ZKBDBDyZVGzSpHNvBht9tCNUpAc/1eSzao+AqOWBZc9mUXif51
LijyMv4omV/FC8k7kDPCWbLvHqKM3fYmw0l6b3Rex+Nav4Qhepj7BeAmyLFQYkUDrLfedQ4BCdjG
MIWZhtHHBUa37t3iMwX1oPNapvBGl3MrUMUbcMN8crrz89pmvjqngmogG6m78MnpM+0VCA+e9/qF
DyY20HKkJeekQv+yi6Q96hK512zFjmsght8fANLXeTWHkVQ0AIrDUBg5Enp/lhA2u03KYxXEFBdE
vdVO/iNSZTygMfSPI6fIXrUgajKAi2yFnfkMuvO5Pc/md3Z61MPBGbYABpvduK4HE0D4XuRSp1UF
u1om/K0Giav7pxxrc8IwtajhBWjKe3SVu7Vtg7Ea/tW8YQaib/FOnWetHuJENVd6R7AjRZLQyUJ1
fJGhQ+42Pyk2Nf1fkUWPDQR8r21VWFXaF0WH9HpVlbD+TBxpuAY+otrzd4kRuHqAbi/wOAfVFyI+
qJpUO2dE6vuzBmbiQl4eBQyJE2NhcaS+ZKKRIAdVq3+Pdrm8ATLueDihZ/bGCLqMAVRCLDUfFHms
MCM7Y3aqDx2i4wP12YPdQTmcr7FEZiWezYMJ3BEFl3OJ61Ro6fW3bwLf0PKswzIqCVBt2Milh+b7
h9pFYI+LOH+n9LjLa/H6j7IJWqoiRcORNR6hYNL2NguvpOgNGTwbEH4qZCeVtp9WrQKH2WS44VEX
WXXXsSo63+rARB26mSYF4uZkflYQM+0/ziXffjMCfrLFAoXvluXnNcKL7hmb0Qp8dDTtP6xd+JCJ
E2U4zqQnfTxlk1kGT+6o222d5pwl6wC3ktK36l+uLx3guPUozudws4wTaCpps+p+O9twqaQw0JNq
OZfNb/jSXED9iB0+C1ypD11vceuE9yQFmeXbwEnV9halCQk0jypKmjvybxiUKMb6+KbEqHucRcLg
diuWqgcDoGo3lEjY3JrqSWwSnU/0+OYwp3ec5EtVj+e/7QXxKVUbad8W4P62IvgRXv5k9bj4G58l
ylcfFAoOqZNK+SU1rtXh6df6zmYiOn0gcrNWsqQ4yZPym6eE45XLOsVlRa3TIsKUsWb3C3LI9NPa
2eYMn4QngMGfDvQ4BuXeWNgu1rZGt+OdyYUHO10WBPf5xXtb3IaEWgUK7hT+iar/L8MyIdvhp0do
tvPD5hD8qQ6tvZ0LEdgyEZlwgshYW3NPoeVHD+zJxUkszx1pDkBH+rUgb9rJIVLqrv5qVtTtJzk9
3PUlNPFvED1gH6WMr3kf6+3XJKqaiIRXsgdcHScSFP3l+VkqWaULTtR1Gs8jJHRHP7GZPg18R5HT
iCBY0/TA+QVZoaUYz5nxZKmiTw3fAJy5mhDD4v0jn1Y6oOyscsN7RAuI8oJQx4ojza1jT6TZXUyB
0BaTVilk+qcs2p6aE/oyPwJ0Y+sWiH2nGAaTfv22RDXFiSvOlHFn6ut7+Gr6Rq+BkMc1oHCDxVyE
2DxvEXzvtV0E6290yWOqQ4JG/gaNlDqErSA5x4r5WwzNrl6YnGx/a6ZE0QK4IqCdf4NNUaX5rfXr
xm3QuzwV71NyHh2LgxF5bJ2JfsoDaTdZcliocLnkcvllyLB6p4ijpIP8COsjAtlW6vtwJmAaCIUm
7N2vuP1Z7pqPok+cZcz/uBIbPR7+e/2/X1/FNzkzd7hZYH2i/QrZjmM+QoNBKIR2+EQRt074VTP0
kDDuesTz26xLegl3G2LDipAoIfRgUUVEPFPBOIPYCcle+CWgrtx8O9vtObUwG80DG38+kyEk8vZt
Y9JUnONKHm1c+Mm7tIpo7SLU7R+iOa0xzJ9TbQCexYKRmlKzJ+wYKQaOnvc/NA5dveV1LrFbTChl
2Xi3Zs+OZBgRiqbTAbAJDlF/DHpcIGD78MW8+yo80dDyrCSqDHXNgFj/wHXddraGkE/Kwio2NADi
MwKdxgxdUxzhnb8/qO0TbL14O8SYbJHM1AxBTQRpsihAjoVnx2OQXIaAbf8CQfZ7dyxoZIYcVJvT
H+lVsY6cjKCjxVpxcnLXdSaIjrmHRDPeMOae6sbfm3kWckF4nP28dSsUO9AhEfg0iY8EOIDlzIVN
ajeDoONTkKOKcQ2Hmj2uKHoDrN4tR6tiiN9NEdtAWYkrtKAYPVVaHN34fbtFAOLSayxyq68hQKVD
XV0AJjHWMYcZRTReqbgnc7rcyk5sH2zTYFvJ3H1H6sl3j5BLFZn5t4SpWYoDS6acG1VtUOKsX+qD
mhP7nCrWc5I6R2xP5fQa2yo3UqdSHWgU6tyID5YGCi3AXKjHT8EheyGib3P0+E9SCE9/rJ8b9GzR
6ceYtZaaS5GIqhdx1E93+zhCUf1gwCr4F07pj2+vKnluIY2Rb5g+6kK3LXNWv6VjYlqWA16Y8Bc9
tBaDT0Jo0+evEOdEyW54BAZ/0mtDpVlRGWsNgPzniwnqU+Jg4maGVQ5c/y65gDUK6pneQlW3eQ8W
Rw6BvCY4r2B43Pezu6fLZdOdwmypZyA8keh5UfD2i3zjiAKoW0T3nAWptlcH08Hia4gOFLbdITIa
yTFYwk0CmTUk9ZIIwch81nQVVOFBZYaimPfNJG83F/RI3hRNEx6gBdBrA/PlYjM2Bj1+cz0QvVt5
Af97EhHEOcwt26PUTZCYUDXSquySZkK/14dUyS6ETN2MSJbjbw6r+VlsfjB1vmYSa7Yw2XSKT1fT
/DFJ7aeUog1Uz1IUeMcqVspcP0RafxH1eQQsAzO7c8NAOxr6tKZnj72RvJF7hbKEXGWJDOWQ00mF
wUzg2jRS0drecYLDbERLg6tnK8MO4RiMWiSSMFaQS7mQ91aCozF1Jcbw4By8zBvMvO+AY/MagvlD
JhEPaRCSXlosLF9p88kpeh8sPg0NZ0GfS3xV6M4AYSGK6A24RZ7zrmcgw6AuELXLcaC20RkYOkAp
GvvBeN9i8gLmtNoBFOG5PgdLl+8nzEWbiFzNtdQeXMrpAqZNu9Acz85MHu6vZCUbh6vJmyTFeYAQ
DWuOhIdk78vNG7/CWGDsdSPJbblRLCXEJroWGGefEaGclzZmtTHbNNJHsTcpjzHlY25lvBEqznmv
gdX4nup9YOIB1rhHNp0QY/RyTQoWpu9jbxklNJp8ox4delFhjzNRC/jy03wwNJxErcK0RSuPCNmh
9BDQOh4qObYmDEdKqroRIx0wumfNrzNNg9ruW9cZqYriy0oFD73NOTMMi+wbDVnbUZaPAIptBQHF
AWR2KlYKlL95dHjo3Cnls90UcNQ9rYM0iQwZ8oxTwmxcqwU4+9rZLk+UsZmw6wwXKOCfV/udWkFI
UedfJ/z3M4Cw1UiwwXGvuUKg8lGBq+sxQwzWRXNwLgGHgNdWjqNxrk4QHA/SO1x7vpZT08BkXd5O
bPX4/95leoIKK551nqilcJH4fIbt4nSHtS4++N4zvxzkh+SdtiIXyEzrNlEtqj6moa/ahLjMkzTC
P4h8C+qxR+t4g4uAaq6MerXbU/Xc6j+3Ijyg9ABEnRvoSQXJqP7RWfhH4Q8DbjdO1oDhntzqrKhc
ikOv0asge5Emg0ewm10RZYOTNeEu5ZZdpVxRITvljGVRbkOYEYU/obmQ8Nb8YYoRhSgy6geON6/p
s8aEYv9gmT/4RVIqhw0fXW9mJ1MB1tP5G5bRySQg3V+tbnUBa+fuaRO5A4kecTCqvtfSMxG4S3fy
bA+wynTkOOP5SNBAkhw4KwcsAjrCk4AwDDN0YMYvn+UTysboK4hWeYfmmU8H4/qwiLOXx0CBJqi4
DXgmfaPv4i6mtXKlhZAZxbRb3pKFCtJxlAEPl7ex4tO+WDckUWCLI0LDxH8Qnf80nqG/dcxx2n0L
AygWyKjw62U//tLdHBIqoXP7ruhgtUdn1hfyvUyHaFUW6fJG1D11axOLtfM5fyP7th3y1HoKJheh
yDtqqzzwPbKLTjCJpjtm8/bMms0+696feaiR2OJOWiB9jgnpML56Gi3dGETQ4hnxjDLGws/mHAeH
QCIVGIQPFN+KHfIZTWl0SXASstctHr8NWV67ChJU5TqXa+h2Y1zDfrGuTqD8zuU93C81qWbM31fN
30Yg1eRTj6/w3Ae7PUfIvfUHkT6auIhnzIEx1ZwLsRkak+vdVtQbqGMFLqvyjjmYNyVa6SbX6K4T
4aqqhuWiGWFdCaWrPu2jXGayv/fR6Q90XyVmbunsxPFrS2esrN1GoA6CLpPUeK5cQ9XkzArZSfR0
QJLUxyNBb24kzMHsVcB+LrHyioMC9CAf+/QiRYRrr3i2dLq2LEHxljWyukc6kRMvlCelss0S42wC
o2U3BEMSAy9RtVraV/6q/1DIRWeR9FB9Lw8r8L68rPQYbP6IGUlFqZ6n/Vx3pQ4BWyUCglxz86tT
kBh4fXzhwURR8xs/dM9xsEOIf1vBX9NPh00scaEO5IJ6KDIG34OG8aRpwxZeMUEWDQhZpD3ggghV
e8aNyXvTsevfVBrN1QsOk0tWKMhITl89CStfpCN+T5HE+OYiVUf98Yx3XJYtXinJsS5SvWPuRxc+
+2ni0Yg+KI9qr48yw1NHsfL3erVYy0PU0vawCrOQj5jHQJjf9oPWLnwqLNn3oi+x0n0JWd0HXEm6
rUY8LDJge1YeCbf/LaGRUrbyO+1/tYjQtcCENOia/iV6B1QGquaNCcaO2C8ciFkLVDldlXjp8Jrw
YPCqS1YfMt08K2bnzXX8urdGPlvHcTKywNzV09AqFhQfykS3eXdXKkKhI6pva6gQnj16eQAerVdU
8TG2og1I9KnIcDL+22Tu/lOT7ybv7iRGgEETUnxucxqP+o+op4TvY3MlzNGGNTNIlSKNAd4x4X0z
OTETNTdyl1AOLKE4f3wGwzPglvLOAaKepX/OngTlACtYLib6d5CIKgN683Pkv11g32rqduLLw07J
pNop/Wju2Pw+eSAZ8bwcd7ifrUyGfVSQtk4OH+eGFtbIxDhmMMTknqGQfSeOMmIk6XDmH17N4aAo
wit6cc+8EjnHgI5AnzQQxXvuWBfDAqY+X5SfK7AHaGFB5ScludG3DDNCuPA0atydXqUbyPy22o2Q
BLltt+ogxnbzk4m6K1+JQfWJO86oCiZG62Z/gAGzFYLmIzULl17W80BvudTrh84sMIovvgAeZ/z+
O9H/2DsG01fj/ma+D8fw6H3Uz1lqUkJ5GVuJDcO0VUWSwjOjw36LRx3j8ASeQTZvyd0U+udm6/44
2CtON0Ak2crJzmyNab9CK/NCgafQ/+EGctTQu3oMp1Pc6ux9YGGFIA8c24D7/8xiVS+s34r64LuO
IppJIayfK7wvEam3L7wmMRJxik3A0y6uI6Nt6C/qUI5rtGoCVF2fUtkh7Ufo2UJycauOIuuoxFdd
GTMCFi3UzJRGyBimfwJI7DC14GOQZj2E51eaM80oYLUEhZLwd9gxrjfq9R7xsSaINPSSO6S3JrmO
Nk4pR5BJjOiHXTIK2/NsUOdowW/3zrpTgXbR6m/lvB4mAbTxRLiq1eaBg9cytuBS7M89bkMSWfP4
QycBXXxyN+MYxKmfGJkW049GBzy7oP6DLtHUvmpg4Kp/lQm+xrJskKA0YAfdso1apGLGghI/VlZG
kYZLAuGh4k8PtB3y5ZKcNYncXAgaqByOv1JqDfbLS+7pR87bLvbMr4RHZySK/X3VjSTRNdC1wzFo
Ze7+b98rxMdYxhSd5mMggw4ottYeKPTfGtvsLQNRBZU+QITMj0Movrhsg2RPVGY4BxFavMixFEgy
WEL/bAWfAVPNCBhjaJR2Ddp6K8NtSIjSxER4716tRsY9iRgfIT+dlj7tYASiph8XyFW26Zz+TBVJ
Wh0GWX7mRmbIeiMKTkJawQjUEl76I3KWsEHb6nmBD728rrDpzlfqi+mPi6GSzUmHNPVt6FuLOHE2
jWeqjWyF5FOoQmTG5vqcfRWcVgfwTZ7EootOAh+E4CIXKX1qJ26p3w/5hGXKOFjjEZfz0ZLMfYha
eQHFzu3SWIHTBIVivCqczBROf8322/V0QAM6IL2GFD/bhG1XLONgir3vtEI80tUs8UqErbhBm595
EwuSUOOc0RWORyzBR7SUtNnkE+ezcLTvwEVSL4gfSHhEx31C82fOhtIqPhPoBLGTGZCVLIXjws13
XVb4rgELLd4CUYrBdU0C+vum9svo4niknkQ6Qn8vZisZy4U8OUoihdghnLFfxijcJ6SvYc1XXDBC
e1ZWRL2/HXAMduAGyWxHv4dbX1FhPlaeNSpRw5yPnioeli3X271l7AGoU5J/nYCQTKJk4pnvT8So
7mOhIjxLHnAmUS691ru8hJbxnpvTo4KnFaF9lXlR9a2TVsYGxyeLq7y8Hii/FjerVWY2Z/Ee0Uzp
MU3t/VDfFxuwRL2u0+pIXTpX1E+cUK3Ttpla75oWKc71XNIr/daniF3KpbWY/GY4vIonBv5cWAvw
7s0bgIsIb5ZBoQNqIsUg1yHhi89Y3VSkHiwsYxkmltFDg5OUxvEQQVKrhaMNDTFGE4H8JHp+TWgd
rAzIozkhpZqoQ9zwAxh4XqvB5n+zWqLPPBKibjq1dCFrrrzBEGhUoeC4E/EPeMtKEr92X+8TABH/
D9igCRsgIvcv37mAoZ7oijui/1yd+LJy1H8Gv1V/kAXmcPBxI6prH/yxVKwh0fS8F425A601GpaU
KRHJO3O/d4TlaRYxYCKCihNRE6rpJmVIM1f4sgQAch9KhurcHSrZRZXdIsQJFZHVTxP7ivkRVpTU
EetxpFQlhUsxH4ImlevQUrOksB/1kx83Dbz1v46yxO0PrxC2plmmgBhGAX/ZYFJ5rjZClHBUaDkB
+CBoK2yxJInS/7kR2vG+ASUMSaE4Tx7ilGNLD1+eOFzugXRUvyXMfmgW2mGOnHLkcMhO+CoMrtt0
dqkxt6lxVJVdAg6Eam3QfAH8cgVNKehWHOIEkXW282nCPOrtQpC+spWU8216kYT6wnv2YvevJMnk
M+jgagIwiBSuzZdCqBQQro9x7JYRB8EzCswwIZ0zqKCus/T90Cn8YXjnw2uVr5rl2PNIAyXSbHor
74KbdsKMlNl7v8n/WSw5/Vr8BOblUECzlb9zPoOki45eYwDESAFBQEurKalsFmamQ48n7gNepkRA
pyIonTrgmdCHPl08cA5AlKmqURLP6Sv1ad2wFSl3swPMv7yT7jqC9w61sVWGYhH4fvLkuB7Ac433
oeEgXtwmj2CMKx9cQ6WY8oMfjM+eCZDoOxKe5Q+6hm72dpZp0OWPKhnwFKWzjputaLoqM1X0WTpi
iOY5t/0zWt8iO+wb8NnfCIH7tLtjBbkLIy6H5S7wXVvMfM9Lda7DREPy3d05R0jZ8BLktdOIzWEI
OivKA21xPs7+NvPp1ytSSp1lpZXftywvxzk2EvHl+l+vVvBdZ4Z3rTVCyYb8B5BxL5mF1tzFW9IA
BkcWi4AHk6G4z/INJHMSP1f5Kjc5uQ7lFDjer6KQ/EbvaqTN0jPldFTCcZRLyud3szQXtIphbuaH
1dyu3SFxfg/2gsfn8JBpvYYLk186FI2dnDObg7plpmAMhUCWMyXPUnqBPONSPqUwlq9UuD6YlcyK
5FRIaX/j/Q+PdPZh48JP2P+92XlaK5zXd1IOtouN1Darxb9vP/Cl9VRYLptkKj5nGSQLbM2mPfPb
yVoJhQR4PhIaxIKfwrGpK2luaXDSkNcAI1vlfSWbl4+2iAWIZZeTsAd8T2brrMslGYU5JmRsnbpW
JCzX258dMBvBZf258wL92S6yCZk4a6Qz6M+V/dxvMyssNh6MdtZdQL66BSjoYpH7I0h1q9eld7a2
N02CNURzUL1P88WR1z+E1aZlWCK2wENMiaRDixvRLmdSxSKJIVNREcnOtSTsQ6kxSjj6fWpdV1D1
loUAoQyg6+EV3X/bBhzKC6HBwBWfuLqsE480U/5B0yCn1Rn2JSXpoao1fcBUbLE2M5A4n9al1qje
4Vm4k+NwWFWZ7vCeq8JUhelfXivbUskWT+5fYNnp2Kv4UuFxhfxGcFR7t/dhdxfQxGYN6SNWP+Sa
IWWR5d7yV6NgoqvntDQtnGKoHVhCBWCRIHTA32/RT1q1CydCwjHAaE5Gi89NfSWBEeAArnJAuGfB
KY3pEAGRDkNyu4u50HlFSar3KJ9KyCvl3EjEoKP6Y8+y0sMRrLQwSgstm6J1PcNwLf5EH6tJA8Zu
1//myfNeZt4x4nobZTmSB9OXskFWJg0VfhpgwFyRz4OOgTkjdP7RSp8NXF1tpoTEBXMrHzXqND/j
roLG5o1qTwJBHcKpQJDfyJJ4at7ETakPAI10b3fek9pP4IEXcIHmEQVJybMGDjglODNqaS1xkho+
UE5rmRkf3if+N5K/eVqIW9vwkZgVkjIQ+o9palJbnj8FjOPwDjiPBoCaaNRfqZ+wBSxdI+3ZOH2A
jX0DNPb3zIx4k93SO4Kti7h8jUcjXrDZT/rmJmOMPSabRHsz6MIuLhLyT0hUayE/yYab/LcwEQTI
srm8YMHHmvcsBYN73z7YmAHYlnQRiJfOIDEDsbXw+crLKCpj/HjOcQtwDld+UXfG4Z/QQFhrg69w
0/63pqpHpgGyAfqtbVUIj6f5vl+AoPCFIag2/G3Z4x3wfYzOhJAoKKAHzF6y2rI+lbUmxQftVA8U
V7wHjZHS2ycOzl/hu1fACnK3TR0o51ppYZqVB8/6yiAZcY7qrA0JpRtB2h3DIW9z0c8WFRpKbcBz
M8NO/grZjAwIX3HFJ9e897OXlXYrHGz52+9Qm1QaFVuj2BYT3kM8xAPZ62GtIXmNa0Gfy5KRh0Gu
pRJlulFZX1HIUluwZ9BsrUOdJ/FECYDSWpGIlun0rsd6Jopgs8Ti33YD+pc91qPoszFGcjRYZoUZ
P0dJLNPAGaGXhV5RbUkDM9RNJKy6bTfeh4RV1MU3W0BGM0JDjDFN7rhTmnCUJmflBdsGnC5teiLz
cVpYJjcPnPerLDIzH7bX/zSzVYlpjMrE7+I+qAVI3UNGSn4P1PfdKgxVO1wO0XL8Wye8n5yexLzq
I0A/tAquzbcbojhURcgFiIVgwaKX06EoIfeQDnCjLJw9UTH/XN89T4FstSB04Iv2iaKRUqe00aBi
KAUG77NLA+vN3CHSomr7MISUvxI7h6Xz3eiW9BKdTbx2EPun4xqui8sL5xzSeodzyHVsrtd06/Jq
StBT+VUrRBiRO4SPlpa55B3TB9tkN1JvixttWYARhTXdkk5pQ8e37qKNI8lUkBeZZ1XkN7+xZNoO
AUSevG8R6ZuCzRux0ty05c3DCXvD0MkBS45Ezqe8YtcVKbWbE+WM7xtorARGYzELXhbavZS04wso
MtOccL9rmPwUoWpmuLdC73xn6jsRal9xFmDNTl2jdTa76C0ngUQUm2dsds9jq80zl9ot38gNpGsg
4nHy7FgZNOHOq5i94oo8VnROT1Yjp9/o89R34YM8uWRoUGcJESFJUMSSxmjR+58EfNQPON1M3bDz
3vg9GhUeUho60L1XaTYU4aU1lPXgu/Tl06El1XwnGOObnRx6LalFoKkEdKOTTGvri9TMD9KIi6rR
mIx2SOHsS+6mJEcBLc9O47zEu1VEWkLAn5Ccy1fruaDLt0UkopNLRfuIwMtZ82HGWybDsoius3O9
mOWZzBPKl/zZMUXTBZvvkOBOaZGpbh189IldZ6vbk3sShdZ+s6JJ3M89J1lhljFfmwCo3jcQw7RE
rndse7LYovx91WrxdczOeL3QhXwek0Wq6W1bXWvH4nfuELBZfkgV1LeuBRJjDTg5fF5x6QLxJXK3
Z3MjpSAnHuQPRi53tpR8b8Jqt8ILJGnep8KQHOFF2trqegGw/PjzBkJzXxaj2KxiAMXY52UYizZQ
dqX+2Y6MfxJTr+xIi2hZ9P6MIgwAQ1xEpH72Qhemej6B0Yx2bAo7+PamX7rnhUGE/4zbWoMu1oj4
gIVAKgQRclDJlJQFCHENHZmusjDuJfcgu59u1HP/wWkLY8nUcCekXTt+bEa6WDv104nQoP7sgjx5
q1pH9BP5Cpbzfw7QYXaHBs2vD9xA5+lsHZhPL+D6g+A3VJkfewvVNE0WDP0uHhMrUFAEtZNgo+s/
uQrDXHI3X+sPYsEFCtkYbAdbKb90H6tUjmFlMv4KnruR5l/xDeXdl8K+7TWpnSa766XmSJrI5vrL
csPSAZTmxdYCvRIyWVWGxny/Sgp4K0nvyzTRc2YGyT2AtdpsAgUuYCA48rs8WGZfHVWl1J0EN7J3
P0UlHMXvRyPSyhbNzceCOg99Gaf/oUFjOqU2hEn0OkM2m698p/wlr4F6IeGUL3yFmBoVVBa1Cphr
RfsHlFIywI18jKEHb0UsH2LWkIcMfdvna4KhMIL4vrD7g/6Ijpcb+5rC+3UqL+bEt7da9nN8YGZ5
ViOk9a9D6jk6h+MWVejlNeqdwDc8yCAP0tgcwPOllOU1tkjc1sBA2RXHkmLfh4bm4oRhhoMgSyyP
SD2Q+gA7/BZTxNPNRj3AzqbAEdSckVDm/Us3MXnNAmXAhaKNwx7cUy39urilmNQ22lo1lSDfgAbK
6SbImy6KpvY418QBZ3E7mR4CSYnhkAgJgdA9zw5g17zOuA0hoHA/oziIiNe0XSzKpTi281Q3drYI
J1ylpP0lhfwxccuxUDekZPIrOo6nf4Nkml92mXj/q25OKQnOeQOpC8L/dJBlnBfDx6FWSMMz5I4b
Wg/VY1eFHthNNL0oaD9Y4lTW8i5FordqQEn2EgZyiaGliwKJCPTgutYUK2DASKNEJN8StdEki5rK
JP7o8oqcLP3bx8bmIVl7cg2ZgMMMprV3wS039CVy53/wnN8TfnEpWLV/1aQDE5N4Za8fpOR5Lb5E
3RrPtyNoxma2Cb6bKgNh5gcyYzmo0hDIzw1w/CaPl3QVNgXqN+JIRSCGfKWAib8Amf7jX/2TIMAF
MQpAyH4xeAiXpX3nwGKFUnxTS/Foy2mC+TO+7io4tNnEI0YzrwgB9jDFxjGufGy9AJXrjIq67vdD
EMR0mWEkUusw3APl4/o2h8q8HsitY69JRV0+AOB8ggJvK2M+X4C2Dae/wFyLweyVWX1ejz2ZFp2/
qdGwfqly1Yea7SQqBjUEmTJoGQrep4TJT3qmXZVl65ZzhxsnbVHUALOQ86YQhFI2u0428F/JwE8H
6JqhHJ+3GmZEAydnEp4VCPuIltVdLHuBF728h9bsyA2Xuirwzw0unSjyji2WpKwPfpy87SuanjCE
UVDCtfmIiKzYHLVS2wGuQYVKoVhPePjBgQT4+rC0yDK0Mq87bqRTCOATrEVdXrhYzwZgeD1t1y+P
ldXay4eVwKYdRQ44VpxMfKRR/ZPHBWUA274Tx/T68Qf2crI6FTUKGWCdQ1Jsw+1YluxmFcV3BAQz
5tepjgjCEAB+jNFQFHUAOT6x3lv1t+8rQZhsVUzkdLp8xV3Zef6WkpvO9Oe+FxD4OXzdUQZeOx1K
rPTU3fHhVtEVxmk5Mzw71ckSJXf0tIvBaAqybfxNa6ZjgQy+u2n45HyCzJZcrDGCG1jpEH/I+5rO
CNgs6RyQeQ1Vk8aaqFz+9MnVCqEyVEIiw2PQ1+9kkb5BzrBewd5qFXymI33mn3FRKdfXyI1pMhLb
8VX51UcUVEZG+T+rUN/o8FO1DSYUnXpjPOx8VE2eG5h/0zyKuWujrtS0Zs4e703b0gnGMLOGDB32
0cFwHzYkgHKZUDR7AXMM5ez+22MyXetFC2CHMpxHZjxJdKddm7unxdlOQ2zKWv174uz6gZx/2mnC
bOxXkIM10jzAvnFww5Q8xgkiCCiFtcc6HuVoS5/W3xSXV/rwCSkFsEHryqM15KdovrDqvX91kwwa
UBgGUdFHty6oMgxDZ06B0T/DmNmUFSfROI9aZx2e/4uhGCtTsESHQNv0jgQ+/QlKMfNVmwBaqT5s
dPba4v0Kku0fLEyGzyG3lTCS3I+WWs+xB0ucJabXb0a+Goa64JGrlovxqx0FodwXQTKRAvaZ1UjL
2pPoNQP7MjilnvazMLs5geqxg7JBfEKKM1OtIm0pmP5sHi2RH1f9PxhB22PRZ4YkMao33VAxdOca
c6YuifTY0Hm5ON92DP0A2R2a+DcihoDTGq6vkx9uJJYdJmjnc6T+gF0N4ubCrcGw8P1F5N+JRSU1
SrC2UM3pInRXsULcI2M8R4Rt4cANUkbF/P2o+Yj0Ou8R/apPNZSH5gW95krCZ5KhzW9tHMIGQXaV
d5wOabKuKKLUPpSAChf5e39vo9Q1qUHe6yr8643mPQisScCiClv8kZvq//TZ+uf/KA2WZHqMh3Sj
dKA/0TUfjii1EFXnDCbU1eNfVwOyW//Ai79uQYkeYCo24+yCnPD2/Jgv6tbbwFA0cGC8MYaxirUj
pAEMs1ikxTobe15CvDpOcEUT77bhdaW5r5rmet2aZnM8ND0rIh6uc93ng19b9nBcN48Qe5pRFibZ
qFkvkRxK6rXuZ496AFBiB/A7H0UMQYdTEGWcxnwweWl9lxpJxdSQIObiOeHJR+TjZPi0LbO9nlEp
VlbUBWSO+H0eWure1Qiv2yO+VefV0Haw1zeuUBukDSsFB4N+C1+kgx8frXmVDlnyo7HNMvR3BnrI
9LOHK+9MID+sZYTW+W4l96oRaTbWHGzsvMi24yfsU9uKqeZTX4PLDu+04BOfSUe3D/1wdGqa1Lc+
iXcTTV77ewHmJzQe8MsTns4qWkYU2Vi0RiriyvAhSB5zkYlzih6+pL8PfzV2PLcDLiK8fLYNwgLR
VkuJY0za/zFForMKgrl9tE2AC8qg03kaTnWh0Vu+A6hDSkl9pDsRaEG7YJY6KaCtWh+tFyBmUy0E
xfMc3DvO1nf/jxtYn7cxZYGp+mkpdxfJTPwP06XUdF3iBt1fmipcUT5xBj8mpsIsD8fW8DcA301c
HO7uIvPgdZSo/KUtcsqEPllc1BI1EOCJp/95In51Iild0X3Tp+kxMrTxoPgpijpe/pMmdxikLIvu
7XTTKcy7NmUjB83MldPbeJ93+zaZK1qMgB0f13ZpoY9aJPr29R3xspmgwt8iWeHnZTGFu0FLvLNd
P+whdyQy36MANZUKs2PR8QOSqyBVvjK0pDquD4ODF+AFnPUenXVdjhxpLgFBVF5A3WXMC2JSILX7
1ka+ARvwBfz68JBEjUkbtfFVd3FuFXmuXKhCx0NrVsSf3aflo1vDEOTxcy8EhDbq3uhT3Pvy1joc
36yBrpNSYT3kxGd489amwte9X1SRGZtwmyg9DnevnyqjPqm03lVvew+Q2d+KxhQ1jBvBLBCVz+Qr
b71rUEfZQ7gkzaTT249jb9mEWNYE5OyJ+txuKJlWsqkPi0J4MqHu/dAvTwJp8NVPo8VshZWpKupt
53gUbDgWzVnjGRKGFrlw/joEYCAnQ0/fN6C6FhaLoc2lxAtqTsBp36Th9Q+9RENEM3ohxuzM3oHM
FBpLa7equEQJ2re2ZOLhGg5eOHFDHDwinui343ZTNBQsLVVEi1sVTCKu0YgSHYiCZhk+IubihhSu
2Er+KQF/7DwAGCzbPNDLCnmDlWXtq5f8laeYsdnSyCKz1M/WruT8a1Gmw0wdXamp/HhRvm93VwdZ
ernDyWY6Hn7/3vXCnh/8/tiFaWah7/NjSvSagRH0z9O8c/eu/uumnvZqP/Ob97d4cfEWUntCUjov
Vf+iGOelvIqtbT0T0ACbnxgkmvp7oGlUOmcB7yLaAkXzwtoYPU4Rp1kmgRTsVJ+9/bu8QLPWCpwg
Yt8cxCuqIIpc05XbZyoZaT3lsbEuRJpOZEh7g85/cM1yd48h+D+jTppVZKe7A3NDnSWf0x7zxQDV
QVMLbPIIxz9ZI6gCKJ7lf8uCafq+oN3dshoIlJT4y9Y4LhxUILYW4abzGSnyx40yI0y3tqGqYS9q
iptiU16M0eJcToohxQmt0IdweMcgZGKHxPGVm6eaj3sV8c/e7NDS9a7bbSOYwalYov+t2oQJtxSg
qtEXIrK6Nr60N7LxVbsK2LpdEUioCbpl/ojge/j+IQmaM2yfIeqGgfQvgkkuG0HdNSxDzbMYXRjX
0XkK4CV6hT9EsMHEPcm9A1s/r9vLasbvCdORqQVcOZFfKo4tVO09vUaKQp8mmBai0fdbDMNQwEBK
uELj9RTlQ4jtayaJgORGkGtGYihV/qSilfAK2WwiQGTrr+O5gQunjwdtoatlkfIFUrnxE0y04wJH
3qgB3c11J3f0N3TrTE0+oLWfMYsPYxXbOFyOgISzkfZpJ4+iOqVbTzeAI6gMtNbzaB5DraYvIo2n
XMxyCYjKD784xOn2nW3U6ouDf1KidtdT7wf+uqYYgi0ab8OOcRSDjAEFZ0RAC6cqt+5GXWJ6mma9
k4tcqb7is8hMd1ouoGvMbipSd0qcy/EiN9i3lXt+EwedcUWnDxgKSTrM99UaqkvGIX8JnqBJuJsJ
z8eZOlbtnfmmdSd5Ud1zIUJKg05VJGqWSM91rVCp+G+c8gCV3gPFX4wv1/GJO6iC4Wzm+QTUiAM9
pj1n8Jh1lLrGkorR1lskspo+NjmMoO0xVOoqmJmolDB1OVCekn6PytoRv5jxIm69nTCjtJzokCXl
C6Z17v7atosYpEecPllpw7oO4qGEma3i/Qmxxjc3I+66OA7oW73YYTWzJhEvIom0j0UfJan8AfQ3
8cCmCuFr3URRod1OZLIZhm7zkI8iXXu053SSrNfiQVOfkIW5F7hK7O0SO7FAZ6d2A9V0z5WXRpxX
8t3jfuy6YHlYq6So3X0jS1lQOz1xCD7NaeaGyaQ1CVTnEmX+HRNFklWavlk/6qi9KdQ3+gQFFotR
RCQR39O5tUfj9hn6InS3KU3x5vR4wz3vUymk5FrELf6CM9hMEKl9QuLCvFGOySGut19Sgo8jDiJ1
Xb6eAYxuzb4dFZwnkj38ipsT5fNBsrr9kBVXKXyHoZB55nhInh0kRvJCaqEUyd7+uWp20ZK1V7h9
rbAoZwebig3rwjrrPjgteMTOm3MxKdawJMJF5dthx5Q79/aB/u0Nt622sB2lMgmi21/UAA7HGopO
nzJLHSZw2GDc1gNCnpsufw2V7rQ039/qHb0mgzLGN03QHMr5Xt+8V4SI0c6+Lern9Zsy+cjA3cD3
CJRZ4AkQhA7laAAwwHQppbeoHOeHVo3sTFzUbLOmt0KR8XYON8a//ZXkMNVF3aw1RqOmVbLiOH2t
uK7HpLMNcP48z0fWfYTHhfcqbEFnHmqcnRXmNk4Ia4imcT5s5TzQcrxRwRoGgjGqHFB9m4vR7ADp
LIs8RBW7faukkabhn0mJsSQf+SiO2Vt4igurNo4vvSK8+qIFeFzSj8v2LMK2XhKMux8m7N2l6+IW
6Hl8t7uMnz3teL/agcJMERab+j7/WYTNUPdIf1MdIW0oMH7gqWa39uEs/5jNefn/Ukl/VAPJ4SaA
kDy65vGlEacYKY4WcQkaEHs4pM/5cZwtrtQFQ06wMe7uv03EPuGOVLppdyhMdgJvv0MgLKUJO5Na
iXy1LP7EId6x2TnhLDWvvsquG/EOcBbwDPxCK+r6xhDxB7W/v7l5FLRFNemkaC2QttFzyeBO4+GL
4lkt1F72MOnw5qCEKXg7C/HSiSKG/3CmolBJM/WPpBX1r8QnKI0LD/pljKG4et9wJpOp6QShSVkb
Gk+/qetw0OIB16nB8CnBG/39kSATLzEOusdNq4UjZh4EmER9gkc/epQNM286n5R8MPNDcuWPo2co
V2O5KthRtt/K+fnh7hJP18Mr5FmvH9dYfoHaVEXx3I3IlKXItVS/grvJndVBOHXLnn26MJ7orXlM
UNjiukFYhu3vtUweZbDJRdxs41AuB2TrQbCimrbpzMQ4DOxp3EIvLyR9OSgSAIk01A2viIBY0+1E
eUJdOEnMam+8m2Dk9j2z+kPekRJKU6t0HSCT9uakhw5CwXdKobRysm5tweD5sPaPXRxVP6Y0rtPX
3IqsY40pRJyWRhvwCwGlg2pS990rFR/g2MMJxUatavW17tRbRX6b2oEtb4ifcsYFKPJyjC3n9khZ
SDpdMb5yscyEqhA7totnaI5ObAj59G2tA3opo3+6G+LDjevX5XLcz5/N7OWYmMRoA5mdbY8ODIhQ
NSkd/xvGa3HXBJL8uwkhMkQq1xHuQpCuJ/HxO/rUYSBHfvuB4qCd+OEkRkeeyBDj7ncBZvcL/aKa
6VzE87DUO8vnkWkOD4UOMV9QSqtDfBPQSKgasBu0IuPcX93Whxz8/QPoti5xxj2yq8jKzkM5b6pZ
zmkLpmmWk/UWwJIqILg0ZVCBYXRRSBHYXTE6BofuXCEAEONBNXzH0yJ1vdSjPEyEkIfToaKuBx6M
+T/ND4XZWiRX9ml0+SX0Ef38caS6fsSp6jWsq29+/0n4oTVZoybYfkdPhEmFo+8r1m1mg1LUgV+r
cq3KH9c+Hjaxl/Z6zZ1iiovyZuh6zreqY4IdD7j+xu7+jNGrvwxS7eaK2uVAl+L8erOrk5TMta6v
9IBNP166puPY3NxR/RWPQRgkPiP/EcF+pEjBmzSR6z52kl4hKFpIN6kvDlyXK8TBcyY3xQh9duev
dguHysquZGBy3NWwh1calIvfTNX+RQUJeV6MaBzJrf6Oy3ott5MSt/83WekcKE/z8NC/kDPqD9l6
S2AH5jzN5xYE1Vvd6MCztaRMMPMugtgBe2MtNyyEbaPd/dmcPMJUoXo7Q9+9VPLJc814Krx/lN5B
06rh+8mjCZ2wzbCIP39UyBpRv7NUtqygX4Q7sO8uVhxU6x/q5b0QZT/vUJZvtLLg6TdY2cGf4BGn
L3e5i3RnViwzdG21ZakOvZ5bkil3PWnOVn1I2ZZsceqYbamVi64NweeLkfB5eYvN+CoqirSzZcY+
I4zZ7CG/JkDVXEuQy5HKyrEUPvQmVSy4F8q3MxrpN4TBFPIKl+4+ImEq4p9EVUWBfIiABRQAgznf
bDL9EJucX0tFWIyOJqxcuJRoUkCoThx4O6X0HZUQRYqHZOA9BTLNF0JoPlwpr9t4EHOzxQ3zVfZQ
z0+AVJdsWueVCVEBdl9tVLhajyKTM5+sbxlkHMlW4l+5lrnkX/C9T+c8qFndo24iomCM2wPukc6v
u5CG9OFsbCN31JKbbsQ0WkxmNJVhUMXTFjtaxhAlYFrqQfUCI4lBIjg06f3XfwzO4xfPvyn5oH11
ESHrYV9t0T94O27VSQRHfIIRySAL2uvm8RV73CmcvHl0nnbT3Awg/aZbFO5rhj5jP3+FlKJEd6s8
L6UufM+toPua9MK48PMM7G0uC6QLq8fNf3QPF3IOupAEYHAEW8AWeHIE+dHVJkUSPbH2x4dsl79A
utedLkEcGXGeioOmKTIIIAlaQq0mJt8yVlUpoh5QM1PPGAfeZQW5DScOFpXkF5vwg46t+KxrcswQ
Y8qU8/PVvLPQijCB+DWUEXPiyljcD3WZq1+2YNjTEZbfStTms5oX+1hb13IjFZSaRzikWi14owrd
DAOJFI/5gqle9X8YB9kmL732T235768/jD9InNfsNuLjuISijYIS3JlY8hqJdJHn+TKSPgGI6K55
E+jFwbw54gADmyOoPG9wm7dtRmlod6n2erTG77q4gfaoFTnaBIBvOi9GyIFrLK4BbChNKTPWye8k
YFrCyPTsgLqZ+7f5ZG1HXuXXe93kvm/uR8dbFL8A7yhGUnQbO5ZO75Sl6DrCnm51eDcUEeTkkAgF
KVjbdZ1K9LVoTZ5ao+xlTt6GlB45r+5v644VjIRoCRGTpjS5xIt2QEtXBxLN2HyJOFjwEdGE9TZD
gmX0vAkUsyegPn2LeQopl1InFF/YmseWitpm8hgG0vcPLpYqfRasy1Gp3mUFu4/ErEnZDsb+BI3T
7MLGL2eUtxrMdvs5i1fIf6h1fStiAo2NGB5mlI7sMJ7rN5K8HmVE4Td4Yp6t4ACvPF6QBzIqJvDO
9P4tUICL6i92hxeYHNR4k5ey0lndfBJ3REDMm8Bx9+Ej1XuGS29YWMKgSUuTaJytPhvSgTh5f+no
xe85PKSYSfHjQplZ8/R2U5q+2yB8i6XcbGxolE582NcId8oVywc1U/L40JCzvouw1v43v8l4/AZn
6c9cWQbuJLSvLSaPRX7mU8StCQeMbDUpJMFuStp9UOwzFMD1s6WJ54XpFB738uSkBi/CcZQXkuGI
SP5PqOLa2P/SspL5Np+aKd/slnx6saVIjFvb0vWWp0zj7LhGMqi+QcXqJgxZqcshvVazhI4zTUdD
yvcx4KSlvebKwmjWWVtr8afaroCDaslfh5/ivEhYGFAOS42uJnHagxherCXJ3XHuW6B6nmTF6W5T
o7eS2JfRenEmYYjiSByPCkbQLS1I8nDeFQlwQq/lIVuVzmvZ5VdpZx7L10m5C8VjffQgisIC4crQ
ZQfHeImYClkZiUfJBxeZeInhOaFFZBMSBemAuE8QwSkk7SX0m5kLjzVPrk9D+FHSjOgjDBAEPGGr
gvb0aA5SnkLppvdHEwPMcotb24wGnI30VElSBkddtUsn5xG7vvCYn/vyHnliQ66Ghm7thsEnFTun
newC0P32x8XdIdN4d/IqEj17+VAxQmQiJSsk1UVw+w+9Q+cJ5jz1O/z6hryoR4g03x9++Ne0a71+
FvTgVC2+ls5WDxhUToz+zzF8qqTO22Tg0sGsI0MLeD/GZsGv/GnqLyojzbZszokvA9ooS7zvvgDq
PLcqQRN607c1G1VWws6AzLGwkA1tJR6+4QC5Fm+6KyDerjUSse+6geEzM0muUjzzFHdXxUSbCfJ/
NjZX3N2sBVcYQAwuBVCjWBnlnDS0K42MuMN0T6nOeCetV0gEGh90m/dWA0vv5B2BjP58CSgchdv7
ADobflBor/1PcdqsMaTRNvp+AXfKq3l6gvF79njuzru0O0hu4kC8PWeP4S9jh8sm38rb5jjIcHwc
oLGEglRQ12hJWGYUbzyGWHVpiW/Hke6uXdNjWc0/xaHG1fACERv44fUXxDcDbw5paYVQCXuFOFtI
KsCzs0IXIFTkWUnQw2swUBRWAaC/LOgnZEl01CnxZtBTF9yFgaaM/Q6EZsQ1PM6Lu6CPosRE2SAx
JMdFSv4zZqk7z9AKQtH1hSpuLcWxCt4+GhaafsICgVpKBuSceFPWpJpki38sCwfqskXnfjtAtxoy
av4KFtYsppSMGm9zbjug2j89MyVqwMrMuEEuSTian2zuwIU98GEoxgjKM/NMasupvaKrNS4Ei77d
n9a29eCLvRVN1Sa7LjbOXsXwPFE1xadbCY5g/MmhGttQqlQdcC8IOfY4WKrxm819elmFMHPfGmv6
4xZXXufNavuoWQUMVb3hJnx7DDOZHk3Da4H1pjt7VE+2n/xExg8hQQdKgh+cGNKb33p3uUukJoY9
iumEj2jr2BOf+N7QEo1LqxwHODy2s6bqBxfib4JQVWBQjxnTgixJHWcz0L7ZOomGrEuGzdI86KMA
Bac7caZZPbFEFWcjBedKR0R33qI8TsdASpNhkyeeITP7UrEfRej7fnziuHUSAeObrO60/YRJ0BM1
tjUZ1z56/ZVnwX6vavwphJquPBsBIyY9czUaUfLSvRszVUgakP6hhq/JY9ibGQZaAOeONPdtqUlQ
JDqCCdNk+XiJCIBueG79K/oNROtH9HHoyU3HZGDUk6mB2mtdeHPRY4mOHnZfyhPwCkJ+04OXqUqJ
0uFpgh5mAwYNQw+l8fZMTT6h+ipHNGWsMSVFWaNJ8jv9CQZF8MVMducJO0ga3dWvCeCKOLKy0yC1
KnJ0YyIPWoYgMBGwfXH55Spp17LhT2zde6Mrz8VIwNazfIRyn7GW95iDLpZ/uq+DunxpIravW2xI
BDoCeo1uPr9Ez6XXz8R6uHZBO7evq2uQE7TPuDHTsGjrVARyMaK9P0N1aiFVzkHfS7i315qq428e
3MZUgs1ry/oaR4CY84uXsKRNiFUagM6V7f4TpqHQFmum8ho4I3i9bpi6lspBcIPKfhaIs4K3i/ge
uBw1pRITjlrzeqd2O5Gvs8047hlYCaqKRQkANJluam3kff6CDG2CFJs2k0ll80MWd2YijUOa9EgK
23sQ2QCdQNkrHEZK0B5U1NlhTKqlTWgHnjENBu3/8NccZWmpv0mYSHV3Omu7YeS+iD7yTawlbJuu
fzozxgsO09K3MAarmdD/lCC3Za7MV4mIHoFQdSN0TJd/jp2WsLOvtNGTIc73kPfaufaILLPIsq/j
FNgTzGL9cUZeJ2p9Ad1ZkECc8+D3i4jwOSwNwjYgoEqdPgQgkhiqlrYZ6mOGchnZjhmUEhHzuokh
3aXtuTzKnm3YfGedTF0elq6FNN9k5yYHLhv+zn/evInHqGiQeXmE5lotGXqWGOJhN2jPWVxmJu3E
gkmPtKKts2NK5JhxXBI7TbU6Z/cY5rHMvRcFjFjgbdWEq35h9W1IZFUJH4qy82sVlcR1ux1+tYSV
iqwYwno6jOQsXILdD8KrIOSr9sFxDcDmW+21zzdUzn0s/cvTX3ghuyW+EJNniptxD8JLYapFWDSI
Vm8j6f6L24n7xqR998MPzTkWda0WTx04j/oZXs5buk1eTge//farI4QpLCPMdxp8uhaBvnN409PB
orlPXKjacuFXXifeNDZwNGO7N6LuD2zq83Myxe1I2BQpuamJMA36PGbXfejpgg/YStzbsVTz+sDA
ecibeZ+5wBa4VH5oV+ePDq8YhzLpnoNRpV+r+txZsq4xYIaEgjK/uKq7BxHDFHwvTJplIIZO4mMD
UDb5XomxICkUdsHcnc03A7NQNruHnPgyxFU2FuizsJni2G0ZEDV2LGjFQBtjapR8On+B+BmynV2w
Bq9QS4IGvqHkIZoKEVM/IHd/+8LuzznDbEjwkjXPb9xJAWWAQXbZRElfi0yIa2PZQYDkGtDvd9B0
s+KD5b3zzQd3q+pfIhf/oBqRlD2U6kpGpyq+DoU9ApBFUly55GIxBfzwKuyC0wa76aKf10RTUn/d
cT8TyaP1cSo0pYtO2vGQTgaAhRoZpGgaJAyCxXfrH2fi0Zz0p7Tsf2UpPNznNB9ORJopwsaUKlEi
X+5hPWPR1eOdTz1Q4Scxdc0N9jL5nFY87zaOTq7tSqKXw/HqQi72RU+mXmyd0qhvgz0PLAQeMDko
al2O7zvCwP1rNw7FgAiPVgaGpc/+s9ZC2wAduy6E0FKez37wo0hC5O2gOeOeYCFvoSHA6fS/Zzvr
fX2iS/4DsD2I8K84EGGsp6blnnDj3nLaYEgriy+Pb7nwDuh52NivssO5XAw/HWf9CvF0pHzq8UQ6
0el28hxsrz1cls5VZPT7wxri0PhFLdDJroKkYGG7D7GfFYxeHGAwY8xiqQdxoFcGwvk8bmAFnhO3
6dY8AN8BP8FwOh7Wg99auxDcit3nf3Y7pdXCi65wh7bBNA5Pd+OrdL5Fb0ytD0W2TERgdGES141X
41aLYu0mvTYgtzL/y086jEkF6LdFohV+UyF5XauJ8BFJumtmeKGF74kjqJsz2LR8ugVwLhUh5nE2
eybgwgoAOQmFwlAMrHAzbbjOzPtpH5AYTgqlwdK4sqSlQNhUxr0EUE0X1JJVhZST3gGKIA4GTNAc
+mwSk8tRxRP7CjUqAYG0PqalsZ8f3myX6Ds6dujklbDd6rLevxlLctBJ4dDBea9yXDXhpqIwm5dJ
m2yJ4Ln7zV9NZWE8n7j61j2wuyrHG02Z3oia6TlUevA7Wg9rl1O8m3LWrxTVZ62OxXK0bcApdHHB
sF2Oh14lwFgdlhiYj4cYqjnXmW6G4VeXkigWTwR3BQ6WKkX1lq2hEXf/i/j4hCmkHJ2EdBQyDV/+
tObjIACw6nnQXGGSOyaE9oZckx2DKZBBslOFnfWzoFqqIkLhofQ1rb1x5UEw7XcTqkLCqhjvKZJq
oZLNkXi9ZrYJkTOwnM47bSHFlQMvWM/vpwB41YmH13m8cOKqHFpjxuSMWHP3aT30JyjS6z784WMJ
PncVImHfwZDDwmvMI3HrdBn1S86USSw5eacV/nbx+772e2yG2OevUFqT0L0pO04q4DDr10vds1gL
n6YZu5+3inawIUqzhuo+iQIvelfzUzHerlFneBFG48Hgm9udl1nDINw/BbzFE/6grUmUX6SJDEGF
ri0j+Ra310rb2pmTdCqehyzLWfZIl5ZtWajH18ehTvIiINJfrJE+TMLMN6OEPUv7xK6C7QLJGN53
IqEu3rmTacbp2n4As8rnOdsF5y6gTjgVgy/XswDWwxoMyy0h15Y7de7ZFW17hXazS37NgW5aSCPN
ydbzlPpkoFRLnTqcj5RGHZA8UMlMuqbgaoaKprfoMbrqC3gGjaTdLd/BvMN7W8E57l8vTeKwWKOP
ZyHIVuQfRsdQtqUDYuXxYOf+7h8Q1M6NKUBt8v2FbuUrtkspqbgE60Vr1DqQZKLtC+qOR2sqAVxK
TIevUFQiiARmNtgih1je5VnaM2TiYzqSMPFB8DXK5D8hTQlGjTDZYXc36D4U9kB+ssyrS7e0l3jq
006L2dsDdb1RdPFGwKE5qK01oXVyr4v3y6PX4K+Oikmy9VK0ICKEIHr148UEVbIogQou1R+ICiqe
YqGmMmkCxQru2W4m+Y8/mJiJ3IU2suLjVanKILX16Kc20OepvS/P0ZxML/d0Uqo0aVodVFEgOE89
IDIfJTAPrgNkh0Gf+y7WSjNmKpHuQbxZEye5Qo7P9ws9PzZJLhtWelYbyI8ZLpSv7uM6MTxbr71Y
q0rvmJeArJ7Ox6vGtsFI7DXA/ts3XpzcHdH/yHJnKcWIqzCremxu+/DY+lQShUlDHfhuWRqt/wJJ
xvBhwMR/mYDRS83mZwqSCfjgMNmb0Wedu3F+r2Agt2OAlIp8A+re64Rg1XEFqZeTB+LJfQLVeESo
uidTBH15COctvM6+l0mOzvfvqCv6JjxUpZTOCVImObfAksYySWFiF4jcKibafco3jT9YqoTPCxAu
+jCuzQTsd1jzcJAyfNat3Lv5M37R0PYbkO3TsedMS/AbCSzvZcI/jG3DN5gAgc0DY9u1hNgcP+jY
QLPneD+7grzwBgItmaPX7NOsV5XbVc9e4bh5SJ4QZOgN3kFmpTJU01L7HFTFOoBh9j7DZfSRwmyy
6Gr3ZKDal8vl5KcKTrLmZBvMjbiqQLJbUv4jbzE+7Vy4bgyxrafq66vylGyatsmgptjSRWVNVV+I
tVzpgDeXmNhM6PSArznhVed7dWLjM2j9aaf/uo16Q3R5V62nfTZFFL78ixqe1/MVSFos0tyme9Ni
9FU2R0rnVq2dwZdPmYvw0dEdtsRvTd//YxqeIgYf2q7hLWSKJZ97WnF5vTN0e+y4Gmh04WqEq58B
POuOv6tEZGxvp5hq+/DAu1HemOvUGsmjWTU9F/SbU0riKjGaHyzBnuVTF9HHzeRegSbp8pQBwAxS
B1KSQf4xcM9RiX328i+UFS8IeyuoIxkHtTEmfPGoT3yCwIE/63ZfS4KE8aa4LUWksF50R+OUzS2Y
3B6Pi3BxOI7PPmA7MuKKjoFg3OWE8SOIGs08+oE0g6arr9yHlHRV+LJIr0cfMylSCK14VvchuVpp
7TWen3DALwkFbXJGhnaUST8N9Rp+N0cEqFo/QkWAsRTR47j+wIhQaz50xDC+38GCnelJDb37nIE7
FB7BtXMYqDPv+OjCD7EnNkdnmDazFBp4iNPWD/VA9ewxcF3X6RbfPX2N0rv2ZAV91LNrkowRtakQ
VCrcFh24U8sB2s3rkQIt9Fg2X6urIplleG5ORwWkjQiunvorMojgEpr76VyAfLBMoE2ecnKwQezc
l2idLuiSiQQ0mHO3Rw3KoiRm3lWEALL36wOFZGY/YJPnJgxRhZFH129cisT1zCmVkYlMoaJpyQgp
99Uic/Oio1iJhO1GkdIJBWoitD8el3stfGzMbt+wiYM8vXq1WSadioZq7gEAuqldUN9UhLAgi7Uf
49mLYwUENR4gWICZsCy5m1LVDzgKAX7EUWrGvsBQYuAVLsZ4CbzitHQmxis0WVaZ/w/Tph15CJYi
dmIQ8mdfwwjIlP+m/Cqv7mYpm8g3X0re0oZN9HooMoNlgHYSe+IWn+pCUMhbFh9/gyeIvQ81Vj0W
xid1eSQgt4iaweT9ZTgItoMJuFppgRQ/WPo5FCcNWXqplzE0BHychIcY/ZEk1yE4h7DHw+IUFO8L
pcOR9R20h8WCdxrh5C5BzOtbmg1YeqbteaTFMaa076TALXmWJoaNUV+PTzI49YyJgNk9aaCvNrSQ
HETG3DXppOT4WlSl3wnLhUU8gINQk+QSY40Zk45LDNwtVuEitiM63zlSnD85KOH7j0weN8jdEmy6
qhxAWEiu0OXvYin/0o6mIHWFj2xjdpiEYp44tR9dUMuAymmfSCxjeFhHZDrp4fMYIzETXrHZEXFB
bRay3pJHlFTp8b/HRPVuHEEaoSCnvDjDkco8Z7dsrOxDYHeaFutA6cDT1xRzRgyMKkkoNEXWDCeE
te5QQDWePzqmmF4VQUYkG/P7W/MtQgdqa7i6wF+NZo8vgkz5wb9QZoRZVFwyvyCLCb2jKjJJSqJd
XRvPtcho2Hw/DCNRayE7HqHDhEDQdqbbpu3uz+34J87z4dWqigAmdxVqwR6vCu4QLLXF71YfRzgv
nMPiIY6jyFIGfXv20tTwtlbOvaKHWSQGvbYU+7Q2fGN0yZBgXBooMLhYMeSfTIN8E7cg+5cvBngC
RM+f0rd44BgncXfcqz+OVSFGe0G1tLP6pxt4PoRBXSVM2zvDQdf5vAZBYdAOs0JDy00pMUn5Nnif
ZQaxulsVb5jgWuJ3EgCw1mlOB2ak8MQ2LskhDzaH5yk6tQ+C4EIvefTrjc/Z1aCpSOqXNu827KDg
uiinaZ3PzW8jJavE9A+9DtZIKI+XaOZiwjvIZoccDOjukIuIF9H57VKLymf40R2myTHFDVAvCIHF
u+n1YL8GoFivTlmYcvgOFi0hnb4fW0PtwOn2Hf8uGgmnF1c2Tdi1EZBjiR1k8uW47UvhPe7bdw6d
3MR2ulzkr8LxPqiiGd3rnkaMjuGGgkxHEV6DzDmUCgHgMAkp8IhhC/9L1H8+4kB9NYMLi4ckOYcS
COEbGjzsOp3lbaphtH0brE6ORs7rpboRsf/7CNvhwy1zplrPrW3W0hqdWT90q5TWzBejg+iHBltQ
c2NM51wgA0RSQJYk839DHpmeKeJfOo7Kk8OVfx3V6IN7861kZ/OpQbqCHO2jdgVY4/wYpjhG9prq
glM46U9Sp6UejIoACJPcWpV0RLrI8gAIxGgLQChu/FC+/u/vufcrLeRvUlNhvVzFPchi60SL89y9
En6Hn+Y7oVCtQt1uJo74eigJBYpDjwE0M059f6aVXhwFJ1Hxy9C1bvF03nL8yKuzqu5GobBFENPc
FN4qzCQDYGzwB2OjTPG25qSdqh0JrQraicXl4XYHK/ncnRSYhbh3V1YjhhO9jTHF6nMCI8dg2DXd
GyX8obFTnMkznR9g23RekK8TnhLnXyvT36BRQWSU7KYQBod1dIHeI6Z8lZq+V3jHV05lKiRBWZUC
rieIm9Tei30bTHhstzmxNi3zN1v/NB7LQgTTIBTaTDSB0/eiZRiMTfBLoHQQEyeOWKVl3MXdrQZ7
mNYLtU93J07CQUJxg2QLc/wPW9lk/cmmNN8rah0GqsZSEWtlvEI6cPbV1lsPH/mQjlYLpmdRwjuq
Wi6exkSI03nQ2eLZj3jx787DRwafpeIkFNMgCcoVvGXgecY2OKNabTRlnbOgfcy0hrvgNEYCigtK
Q84EXCx8rut2GEsLdhK2K1GeO8JhO5e5XGtPLd5a5VRVrr0jGuP+vf4LjPwAicf+1ZkpLJ3Zw6UH
GELB3jl93KS9Cfa/T+jjZua+De9HDeRwYLyCIIz+yGK8HB25sMImOl+hf4Q3wk8rj/htvVzLemc1
MecO6xTl4vKVQQKgPKdjRByO20ikAtdZNzpruTve53oHy+gNr7yr34ltBVz48iDAfQv8yTFeyiJ1
QUzRUJBeQVyHA5ifVgQQN74TIrsbQTdTDU+NqRyND2WwF4i9Fx30zo3AmTF0NppBJ/Yr+Uu/eKiq
3saH9oOttt3Z4Mp63DDowkdwtAgxo8kknRCpvZ8YPQBzZNeGXBQ38/NhLLUiekcBORHL7UsJj1ft
QwwH1/fEYffVLLBfDl1dReVa0KYTqCZo79u6GqB57Yp/pHGBCULJ1XW9TgbAHL2OChRepAx4y/Wn
5zYWS2H18TzZLH4ANuboZ4TzGlNz4I8+pT96GEVjAiTGa5yCPfsNfmqwVZAklq6+sG6qmybfv0E0
2MzXUntTTcT6BB8eZcMS1B4fX8noczo1iR5iZrNRc2XENfyG96/n05A7UXSmN8VsMaj1yq/IVL+c
5eMpfDuzgiEcMLC4zs1H1arEkbxtb5R6MJPVzFtIudPQ61BzJ+bAi/eUCEqXcYDIioJQU4HPId/7
o0qPnlplhEbSUC0YND+OO9lmbTZdbKttaZ2Pop3TKBeqbkJGon7GthMujflFE85r9+02y5cg2aF4
fZg8oGSnMDz25gQvWIQHRkOC3vjJK8qrGYjMRAVDUi5y8lhr8VmS6Vd8M5vk7Cr7FskxZNQpjJi+
sQcTHgPbevtBC8IcfDEzsWcuFl3tyhRtMmi4G458u0S5Mmg8fI9/EYOMvHCq+5MMcaY192EH23em
uhVeqjMqeMRsavGkJCAlcvsJKF9KoLE3nqu/xCg0fi0NSUTdeQfuQXd+Uy3OvDg+lq8b+tgrX3gp
ae6f9UYxb2gs+a8S6R83V659LrtBXAeslijxli/MHaWYlDUr6nTcOcBF8RnZ04xfPurKdIk3/Bhx
i20jkl/Vwmsn3/BRrrBj0QatyedjCnTqwOodOZzRrW27Jrubg4iltE+wMnHR9etxSE+BHwjzltr1
TZ3io0SBuakVhtf8p3NEKLb/NoR3Bl3TfYsoD4oyTzPO0yNDAxS+wz89VBV+CJclXRzwmBiAVLdI
Lt/KCaXjK0VydMmBt68O1YrsI5u2v+NO0lq0AF5cRvXjzfMRJ7v65dB2OVJYXPvnQAzus5MMx2cj
PWkqxH7IXZtKejzn50QjaR/GcbhcRBP6y2S3Ms05nRhzCCEqlClGjgVAeBzl5fmHtY+nq97wbiV7
zTk0Z1nrojonIRP5zic7sSYsgiFncfvNkUaUaTGc9Il7S2BaJ75OBDypacvibOorrpb8B9lQpVJC
QfSa+l50ihHn3QOW5ZihJobCF2KgdQW1QdSzhoG2KzWGJy1816xOlqHqeu+DTFREan445H+G6MyX
4hTjlJIGhtLpMyIF/UEzA/CCdCfPZYhjRntdaaePNnG5T3NDFchs8+iyE98M8nTS/gq2y6g7pqKd
J1nevuFhovS6A18Bqzxt1Me4m5ytLoA59b/O25CYEb1cysWqtlVaFxOMdifJC01Z9RzQ3FAE8q3h
QigVMX6oG9cKyh+pg7jyWRubut7CuRbhP1Aey6GyD5vDd7/9Fi7xbDq9uJc3nHl4zDhZPUZvoT2R
ze7z7uvhV45HJ0vALdndPdakz1x+Dt0hZx+PtLWUdyRDFYsc2RuXwiDmY/H3REOdjo4clztNvq5q
xGsWbWDPGFBshs6GOHKs1PeJMMDqwybyC07WBY9K9S5Y2aAU3qjt3VgYwg6+CC2+PAzoPsEG5utA
jaoJU7Tod8/jFMTnVGUAnSWVwLvt0xOV0aOSEVlS15k36oU4WxRyg+KK5YU4Tqw3bGyJVz6zy+tJ
ccQxCr6XDcnolWworDTFboWZGJ9X70UWvzDOhFePS+dqtMXG8cA33CQRoAugHPteRlibzAB23N4U
zY4JPttukKwL6MtkHSKJb2GTAROuCbLYghC0cZy8QwguoaqQI+ZoanyIRoUbI6tNdZaRPwgw10BD
5yZdPzmgF4azUMCCMwwiD+ONsZCmRYmBfoCZKTNwhuSNd6SC7JhBNIlKVh+secJZ+y4HlqP12k1L
7gwGr2JmGEHXjAVQLCGHVPazHzVQ2FkZyceRnHJJaU3Wpgq4KW6suhUv0TxmStwlWAvmUlngxHBe
otoQANsXQS6HjljeKFYH92yS+vd2w52aeW+S6YM25sRXi90WfWRtikDf7JPu2rbFAJnpKg6hjRwg
n5TehZOf2gSgdRvIYBK4XKyVU3MmOWTrIF/b0SKx2eM/DL9KHYRG/2ZmhJOq/kNU6lafAhpYLYbX
Jx0vdfUSwozSEdTuJjpwAzPQzNAiFtcfLlUQVZP58YQwON4MGgonnaOfRzGkrPAiLXM5Us2PW2Uy
elefzg+yUDGdEhaMPFS6i2I2JXEc2pgncfOyVJ7cP7HDUBRIee/O/D7Fi7byYApegyXJ+3kZqYnc
RCgqiR/wiCg9RudfCqBJ2O5Dx7XDVPgS9nO/ExImfVBiujR6njo+e4U7XBUnFOrQaJFlxrp8ZBGJ
PiK8LzEGURjDJgbROp9If6PO4ISb1/wQI20kZ41BR5HNOYYCWgO/3NA6adznfOIvWScMxMbRhuyd
Dgkup/vmbxd+LkXCnNimM9M+uEN2TYC3uP5AFt8Fs0rTSRwoYV19VRvHAQkEbf2nAW4z30XlSwgE
Ch+QDQSVheIMqHCHk/40AwqAZzqI6Z+Ufsdmg0fiOIJEt330VTBttG6T98gYzPvNVRIWIo8EZImF
4g7k0UrosbQ/z0sLhOZaThO3c3SECY6REiZj7WOkXQ67wGQDFtCmXgM/+Mxky0ghf2Wp5rEEhjvZ
NlPZ4nmY02d2RQogvuoXLbgs/XzlICJX7pliencAqXzWACUIl+XOGCbt+hxvO5MPpkbGXtqqFkva
6EM560GRRY5QkWXtQMjRU2ddQjUwRiisBfN1vkHEQB1uaLzhHbzRGTOyjD+iY+6pLeyjY5HqzXE3
A/rIplRoRgADG/auLDVd434kPN7eNRwlus+QxVC7usZbdr4Jc8Aqn0/FmwAzOmodF02AEyZr6Scq
ySXpptT0p7A4RIAqDBt7g4dP3vXqCvg0pQ3wcTYugEuGbhYkfcJpaK6OIqt49negADl73YB3fLEL
fgkEuuNHnbrjZMnpZnkFbx9ai4tqhDo6Ue5zjsWkLvHSZR3VwJfeHD+G7taHn2uPBD06N2QU80jY
v81nnfDsh1KWpqdfg67Zu1RL7H33JdggPs5RfCKJITrGpeMyhWxtkiTaJaeM891t88Fjo0sor/Jm
5rGHvw8Skk1gnXjhJU8NUNuJLAygqz6TjjeVYpQFdGnu0uFEeEP0jcY3ove94WFI5PIXMhvEpGUp
1PT76XqhA4Kq/G9kQYZ0v9pHbhuRACBdBqkwq01C0bTlH68mctJpQNYwxtw3gTUmoYQ0xYHeXZR8
nrQhXmxIeMOWBQfqzXYYvbRtU+6Jlko/2vVS/2Wozr0ahdgw4hHVx6zWbeBIRae3b3JtqSR6Yo4i
N/ht8pXHwIvPMchRHU15CkVMy5dvu8jjDQTK3TfMAizjyHRlRjPxRLYVRXTIE1pLaAMrS3wiT8q0
UMuhhAnNN52XAAjUZi2CSIa8QFIjGDSP4zOK4WbRq5xaLeIkW5eB+Yx35eh6YaX6qGP8ji1BppEk
ju5GB+zlkazPRa19JzsWhsyLGu9Te9poRSULqkXvr0Yh+q0hysje8Vfq3KpZ22+N72CpVDFZm/2W
BXWHmaVUmp+Fe09xEidFcM3YH1HlLf0t0luaTXGoCARHgKA60nPKFhoRgHPUR1N81viySybbygWR
B+CqdIvXKvISlAX5G9rJ++cyvXLT586t4K+q7w4AuV/b5sICcXmBlNErcQT5FNUGBp6/VUCTrvCx
bUihfZ/4vVwitkW2RZxBgvPVlWbJRbiVrP9ROINOcIxA7gr5tSzzV+9j31qfS59TJxoRlGmyuKaz
0PQ5mLZujrSmvZnaoyx7H2T2JMaVK2s5UezbRswtF/AAE1pCVEzosLxtXWDWqa4ZQxu+Oy7VI0Wq
QuCp+DnzcvCcEfQ2+/xrU4KW6XH80hRh01QrIZTNwlidh48ATnTBsaJJxe1n4ZaKw6hDjtEKSK8u
JuIHuXC1bCHQUvoCIeJ/3tiOXYlXlWq2DR1EZboMwopyIdewkZZbb5brjmZy4HCQbjXfBhFRN3Yh
p2/u64tlIXfzM+KjqfLq3e+E9HV5XByLLYwPcFvHgX8ICbf3j+z0KoaY3l2yJvagVNZ9sx8YQPnf
hbOhDS8m1dJ1Zyv8qIQ+gB099GWnn2DUpDF2S8Bo4gpRNadEIhtkkpz9rLkDGKqZ+1lBfFEtXn2R
VyyN4teIepydxHinTRjv/7ql3vZv0BBdUV5tFQecreogqjyoQpIBITTwDzKXMq/HfR5jcRnWjdWZ
Hlq5r0biHtTLmWlij4+Dk/E2hhxDvBdq3cWDy1UAf5/u7fYkeD7740VPVl/sD+3RY6SEbextnOOg
+NhOJ5jFmGh1fAHCGCvS432/06hQPPJuHi7tVmZK3SK3uykIUVkEOM2WgX9GJP81xokWgrTdraQG
q9JTBgedUONo6p9T7isAom9YZMi/81aUts1Twva5UzHrfyPb202MuTn3rwjEUEPrrh5MbDCC+/PA
KicBTKD2b5gzml/oBXVajYKclCQc59cIYS5oe9fpu2l+x7ZUoBDRLhJlO3Q1NbbdvCX7XXGa9hXd
Gpa6SYbEbOgv4ghkRGicyriKoriL4gjtPnvGhp1Yk68ol8aHQouwOC6SeTDLCIkC+aQG96upEs8X
fJbz/dhnozGD3eDzlskt05k4F5NHjcpv1rrgBunrR0KA6ZmBJyUMylYy/MToHjNLMq0tyLrs0bxk
UMnKgQG7f9ihihLuEE7OzTLJUDEneKITEFw93B90WtOtIYSevV6gcE26DF1Grk+H8X6SOpijS0X1
xQfAbSD2DrUK+ezA5dmm1+vAwzkdJKLMVimF3VL7b0E+2GsZy3N+qIlqSKbeZejBXO2FW94FwV5S
hAMUxgZxYSG4f+t3INniJPWYdHXdggxkHNDYyuE6Kt2qlr5yr2KBZVDp0wmClSEBO/NchdEb3lTp
2cDmEnsypqu27J+MGQSHySUM5vg/9gM2yFgsFjMZCeiVqEKY6onjjou0ix9jsHHGe9/5ugiWJReQ
RNfaNtrJAIbXZJIVIO46mMT7N8RMgSzGZ8owpiQ5S739YKUNssIiz1kEfLCLpv8a0tqeOHxek1/9
/Zez1JOze0ixjW9N6wNjaEI8WrWfxI9nEgE8B06B5+7qMTzpCBNdlJZqGOr0Wh8fF8Pu3T/G21MS
J3je29BKzbXf7pVfW8xJa1Ixrd9SHkYb+/36xCBSe0pQhbgtvno892U7PN9wc1COK2apf/dHrCtH
axpJNutYx+u8l1F/th7RuCHj5Q51ibiraAbWXbjVIl0eRzYS75sr4QFTGEH1vWlp4ZfALQb3Wy+y
MXvrUTzxKJnkVMuYrksiBGOT9AU+tP2ZL7YVuIppdnqKsSDlI0KkR1goCa55OkwDE1p5aJkSxkyd
w3de2U4+a32kSVdYW8e5Fd6tvbiEOiADj18BGPReq0zgvKozVk3GeWPYmyLwsjvJO/ChAe4nG49d
nYpnpzYN4mfpduNMGCDW2dJRsKOCA9K6rff4o/TvK9tbdwGvQnpLxOaYVYeCjKoSFUPF5aZOKpsK
bLMRpmNAInMCWivR/Cfpp34h5/sADDcFqraABCaIyw7oa8Nr6flxfYUgF/A+2uLWRtvSne0LqxTJ
T0f5zQ9Au/mQLWEiYz/h9OKIypy3Z1SNCm2YycsOQIMMeuq1mI6oDRoG1bl88sr50INITzme7xkn
bSM9ujwFFd/Qr+4G85nvnhDQn3MNqxLRm7K2hT3zj4mgF6vgeP8OJ8OqoInC8Xq6MDZdoyBzsfZ/
tMVEgUDNV2fBico/9yec4EDjOlPr3SLKv0nbcWQnW+VWRUF9HUg50JstFRz24bf1+Z/u25MIlg38
egYhA0WICNF1+tglapkTgSjs6gQCvA0SLNH+UwD8XB/ZeEiaJmGk3R7tAagKSOfAb5aJL9EyQPq9
2kfoBIdlNbNscsmu30YnOraqgqMLZ8UyVWPG6gETSZPewV9Kr8CO5k/TdPspD3pqnW35sxvGnKGq
0QD6HBslUveCWzUSUbUxZtv6rxoWbe2GDIgoWFeFhvDclLBaTtRuCaXhhY7amrwpHkb+5PzC9res
cfRhGNhbTThCW3Yi8tW+MtqHZQI15uUwrgK6tIr8z2In4rNMfJo81O9U4Qix+h/ZDffJ2Dni6Aiw
HCJZ9KiI8DImEej8zId469yY0SZReLd+bFXKBSgivmTWw8nMg985EwV+ejmtWoAz7/JLvTwTv9bP
hcnaUebRaEo3vS5YDVyZLtASscaEHrM/huM5YvHcyWkgY5OYeoyfqPzUdM6OTsfeJS/3UE9I7uWg
7UFEf5TCtyc61XqFjOxu4HYBgpAplInVoqVgF0nZ/bZcK+B2DfhWiH01QxUdzEHVpIBqnX7onH9X
tzGU0+w5Mr/AizrCEes7EMvqCsFb0lqw990t1Gt+92lhSIQhJrnjDOpftlbekxH00sFnzU7yVoJp
dORotsc922oCkSkdSPxQTjvoxJR052rGVKAD5rGJveV/RiIBr09VYDHbSAMzJ1ICYg5So7RSml0t
LhAzOdcylokrwP12gsjS04R1QOHkTXcabq3VrHizUMLv9JNBnNTnaWyRiyH3iyNPRl5W8yY1eeDF
glTt1lZUbTtfD6cEf/BHOlrPsGrkkcj0MBQV5VkMYGNNcMgW3My7na7uEbnRLQn8PKJ/kAU/Zipc
cg7aYXSkuwACFM2Zir2/uNHB2gtlkVhL6brTuUm5kC1g0+OnnI3xY4aWcfOcnE+IyJTMCoswajor
LNTmji/uLC7iT/tAR6Nk2cv9FrHHeGD1frDg947PfbHAJZeoKwg7Goov63Eu0/+N1baKYgJPWlHN
q1T6a6GkAgJkU61McNyv8hu6aRh6tzb4bfrAx2cARdcMYZm8mHHltXvVrCGiVzq60kD9QKGPLkbL
WGB2nIWHh94KvStsDdplt6VeNHRHOcmwCPF+zvwexso8Z+NvHdYA4dwyzjhUpMslKDB0HqrUECFc
913rMtgl1m9XhhYD/aDNX6sqNWEiYLvmHgDInYoUARyXZjWqPenwrbVectGW7WeP1jItE6pKdd71
w6Q2Ys3uNXpYLjYjaxzG3YX86HcdWMUBDPshyGIPAuAgbUo4tSHvllWFzHxoVRYzCurU9cUimHf/
0FED4QP2ToV1dngZMgBgbMAVP19SPfrWOGw0oSibcAoaSMJnVjMWuMU0zmg5PtKd6o0XKVAFzUp6
LULQFbM8WjcWpSUgtLpsF0jpIUGXJIMRcA9DLKL+k3TJb6U0GKjLmEsOfjGCs8UgX4Sg18JVIkkv
VkquifdAGynjPt1bxBtIsCxctpf9kBqnewW+3l7sTJ9H2BZ8IITT4ekH/nCExJ9A63rvCPv+7m3T
XC1Wx/8lfIdFH06C23uPRoSBJL4QoD/5mlGAsfVWR+Ez29473VHI475BuYXYjHTbm1GjhAVNk3Hc
bNo8zLYU9CamRCL8VKWbnv/ox7Z46GtG4dJE86quzlwmWWVAQ6cI7yFAxCo9/XKKBSLFDxgcKX1d
OF+ESan6GNdK+i1kWr5MAFPOGp0R76XHiABajw4KoQZtRV8Ex/Qw3qmVqsVe9b4ejHPpKQ1DbOE5
edwgY70iM1574fSXhCrXCvuG+XYBFamC/U0jJ/QObk6FD6C97Y1yJrNdAvZ8CILblMo33H927Gsm
5pIj3csZn1LrCj2FlYhL49xFt+muNP6Vss+OVvBRdPhZzz+SCvdnPCKDPf9Zse2O1hKoPJSuc2Qz
6L3Hq1TQaYkKUAq2y7AQVoDqU7xeFAXVrBiCNrO6DPv/yznFsFdQzzvFJ544e2z1cA22ZZybKUTn
tLu3CiMV3r1qpmkzgiDtpVlzTMCZr6GJWxA47ECXXccX9BHWXKxLvttOks6eEpJw6XCuOI6ALoyU
ut/IBByMyABruzxZFScl46bbXNvPDo966ax4+Xtj8GglgpSUAFeHqHiBM1Op3eQbYSpg+Aghva8k
FDoVsmNbGAWHS0dzdzmPHYrXGgokpBk+a7uhFbkoY55FL5TK0B44yiSbxb6lf/Err37b7tp1BhqX
wPCnP+tGXL9Vd9wtIoBQ5KnQ0gcddwdf95Bw7uHzY5t0SzOflnfyNDnCtZ37hWOyOv7SX02Qv86g
VL13Vlaax+XYZ79HD/7Dw0+j+sidyOAutf1jfBBEocdeP8iv4U7urMemnyk9HNDc3412oJNkqmfh
hNss3oFFIASCPFPDJ+Qt/9DeWacRXeR8VnMzUfikRfFTjMFZa8uC8DG6j7WEDY+wnKxLH5vfgbce
FfLx6IsBIZq/K3aR+EncZHzq9oMKAk5bwzDRuHTw6Fv2YmuqeznsuP8WACOQTY1WPSVsuJ+NJsBB
GRLqtDDpfUyz2TsX1/FxC4DXp/my/lfQeSrr656wVWRsFqBf5bIWTR6H4UP8e6BgFpDsn9nfW9Hb
oEMXmRB8C1LnbKTKWdSTMEVjY9hgSDorBtsejhqOrnidOnD8PE3Y4tLUzNU/fK/uDKH7TpWMk5An
ojg5H3ZxxtXbZgF1gBRQWnbarEEmIOTJ7kaFbFS2wJ6QAAeihBKmRbaZeXCUOJEqtSSBVGCsiECS
/4Q1yGZRGGQ+G67B2z3lnLLy8Wn5A063xzZKCAh3hulYosJ3PVU2m2oIGh77I8uv7Sgmy8Zb8WyC
YdRE7THxLVpxekQJ+6q5IoEYOMTSCo6kZnQB+27CMP3vC6z6G1hTruy/DGgE82ZmWqcNmjXDOr69
b+c4QVRBEDw4SWzn7pSqyTcgmxB6qnxBoP0aPXPADlnAGgk0iOwbSX9wkDhrpbXjvZfTG4O0kThu
1THOeXfb2z/9nd1YTgXpV79HWOs64PpB/4fJQo8PaiHr8sCYycxKqV02wIrJs3lbZcQlTTrGQrzG
8nfUvSaXBS8PQTJuEWjN90Nj0IUbBQ/O32BZQUs7wazen3D7jNOCrwSRGft/TB77qCjAbJ76Cs/R
bLI1KtNmyf5+djeoyQilECD+1/3eBSt9F8Tqm7Eqegt/9HNf1i/NHTNtzZQK1fG+7hsE/y5EGW8n
1vhut0cQUZ+An1eQvjuYAhFZeuXlI7F/c4XmeGSS9ONli/IALp5eeu2Vv0ZjK4WihXiUzYeeVQdv
zyxjc4oVjw2voX1Is2OZZ+s5oUrF4qO7RCcpEwN8ox4mtCeo6L9pYkhtV7xzLU5O7ArYRGGDv3zf
G2p9anLfqfC8HlukgmAM74r5ExJ0Tf8T9tsjOCzbJPU0TWiWJsDclZKSs6VcQdFHNd7AZ28unQ+K
bRx1xZA//VdTgoH0zaAkAKqbaE9g3XpoKociTZMWRjW7v04P5UiJVKL/PvzR26iGMNqFuBah29K0
9uZdzAs+nNIF1jF7IRlggaJUlhSpN2vzBAEXxMeNVLV58T1DK4Nq7GGFscvTO9+lJbYV8Fvo6hER
wuF9SBMkcKns0NOKqSVqOezGZJ6rj1gPjSei4/EHyAlBhz3N6Zd+CAdDiP7WLH2LmGeUQB4YQuQc
JK6tN/NEct0Zs+v6jU6dCK8CO3CyhzOLYAFPOMHADr3aHGV+xfuaZ/php4lUqWLok70Ueg9+8ATG
Ow0oQF40zZFieG1dbvHgSYX4AUQLx4t4o43xQLbS2l+ujX0lpnuml6+Le6h5r6r/0C96ZhkrZEvE
JfCct4LY0RkTlMmJPpaDe89miLTUhXPjSpadH7TfEdVLVISM4JvLzYsEYOMJDu85jtJqT/VXP7mb
6NFRwwfC7H9Cv2zFdh0Oy1I+GIfHuzqRAnlTPjz0ZbJ16R72YNhqaSMn08xQmnqfkK1UdlSxirpt
XxTePpTREsTGz0kFp6GZonKD7Qyb3nx7wF4/AeQBEnE9liVHWLvmk/YA8Vt/OIgzNXL1n84tLrR+
a1Z/0LTourw9nfC1VGB2girxaNFfHFuQgVy4lUZxLAbIuZI/UlhH5EFIWJp+8/CHSlDryJvyvr9M
m/2fXECkuHgARMdiUuSYU+dZkrbOtBZlJ6dAUlOBLqlD3q/vwi8KxMwIO4UMXvn3+ZqM4lnCjYd6
5UGboH1dZNUald4Y7j0NpcJAN38BFLENCuq6CLLmNsf0CoHjtsLA0S+kf+a1mdkWnWUGL9dL7TU1
VMo6XOnEDnCGTnB0WeG1wehoDg9gMXIoC9L6cMx2u5vScQRfemyvD51o2Lh/MqoQlGxOQWgFVIJw
1Fhh0gP+iGXHDxrbUGfq6PHYJyBVnmsyzvG4oZUbwZZnPC6x8ddJGwuoA0Qle1AByAU6XiIz65R8
CfGbBWRaVqvu53FcXPhqBaYd8Z25QuDKLL9vZwcYXXfO9IZ5ARR9gq7ACBnGDClK8i4E7jFuoAil
sGIV0Gq4NRd1UkvQsZ3zs45vtAV76gnThmng+cTC6ZyfrTBu/hhwsiT1vXnpgasbrQWcbZZ6gRRy
YdJOFaxjGp7KruOU2gWNw3PC4fAlQ7QJDwuXd2p7P9ctmzl1x12I54bp89uFySfuzokMBQQtepSV
vyVjC1CDQOMfv0mEh28usY2jYsOp4kDvwFKXcSeh+j4wdyWiChaMXhxlSzscJ76IN9aTSVeleL6Y
IIqx151+ZAJyt6YWJMhj1aVanGAdBt8p/lxvG6oXmPgw5YA4kCAXFoDs75/flDMQYiBfc63CxRrj
8lSv04aQPlE1yj73NLwpeTcQ29hMFwQ0/SKKH6KASf7dDf0Ugb8/ep/C91eKbNAjxlL1RBM1nbvq
thxjyU3QgbfqHjGKO0fVdUSOhuVB2ZOWG2GMiPfLYB5T7yVXAAUXVSj4ESfPpdx+MGAtuRr7+ZHo
WtwDD88PMYi+TzoSjaufe/TJhLWcA4mURwehKnXNsvHRCwubQW6arMKjIiF4fXEQn9EpVuBYS1Hs
iVcO/lWBXcUiESlUYS1HQfZdXbZ1DTRN3Sa49HCuzjW75zwRiMEZJyKgJpQqE4XCp2Zx8wQ+BR3o
TD+Xd/jxmbGtmGu43HLECiay3r1zrZbXQYrJGMfu/YvmIM3syGP7sJCrKmXls+Dg0UEqVaWP9NRd
LwpODVQCMKkzkCyx0LiF+7nmw7u3N+Al95pvLh1vutwoWIO+9rX0yE/m0wTG1wC5PpJh4q+nhM7X
O57jj1datUs0RQe5y83J8EcqEoU/gjkJGmHM+pL0+Lv73rO0H72/5UfD7Ch2/t30/5duOiqsS4Jh
S1cBJT0fcbhCd7uWyfG5ZvYIJ8dZfSvG1QocKYaqaD9TBfOX/mxJPJrk8c3NCvCSMVBo9+S0Sl39
VuqLBLcHFWipmatvKJDmJQ/TmOXZ1/98C24RTaHBE0fjjwqKe3zYLLGXQm3d6WzHniX+uGY7D0J/
tzug1nAJThzYFxztGOefdfBWgUI77y5VZ0NTBWUAOIOyVA555koHIg/Aa66Zu4UFqFVJi+OgLi/R
35VsGvTYndIA1ZKl1bfeRDfiER0dNmDzRXkIju9KGMtQaX1TCjBZ0thU5XJk9GfS/pu+JVMUpEM6
C2NYv7Fxh+H46C69X5auicsPaQxzqKa0gpKLy/IKMYKQnyVWgssC7ETyKyr14v8RklemzoWYHYwl
G8Hy2Rmw5n1u050BTLJWAj+JE+9HtxK1SGhan7HBCP7BLnP56uWOZ8sp1fNuaz4tkYF3Oxx9hgN+
qqgrpuVGFWys/cbWI50tvXLsqa2Ik/NN6tVZHgtCjGTlSqYWS757Hc3qvIKCQII9ppFH9E7LXJsT
NkDw5N2OHROlXebnj+62flsRnEbn98i7SwEshvhGHshbrcOEs2INh/gYEOsXPw5GAly1gkgT3ZT7
0AqRVnPul6s81VsW/GAktiI6oW1pTpLJ7LMp9J94h+iJhT2UyUoO4z8oEQsgBtOvc+eZfQT3v/1M
vrxLWsYcMeVcolrtb/cGBUVBIyinmi6jam5edPH6FC6aITHbkK5HvygwCmQQb6RF9QjyrWpsDFMs
kLDUQK3Wswr4jrzWYMYkt6oItmiqyI+Y0ckjzu4WTM2S6RXiswSUZUHjrXQV8ktMXbYD0FVxDEGf
hpfvHjcj7wvDv7tvf9+B5Vd2v5lQANn3MrgNOWx1GiwsSDykVTaXuvtHSvSVoaW7G6UQOjwIX5j/
uc+kX0l4tRUwfFk1x7Ru4mHV61C6F6RqbC6/KvgE2NjFDZUFbXoehgc7ZwOCLEuJbJJ9fzPqzFpY
UsvARtRnQFM3X1Oe9Jy8AarWrtwy9XQ1eSdbnUPsHBMrPo9nS0mlNuex6EJ65ZaCz/H2YwDXwFQu
+GfMNPFRE7MgQuUuQmFkymjRK5mUm9wwFQiaTs0gc6r4eKeihxui4oXQgVaGdEUt1leR8HewBNOH
z8lQ90XCX5d9jMLmE2IJZOVOC5JRK/JCJw2WvTmIXpHEeOrKEp7cvsilTVVqSGvW1qgOnmCZzQJB
F3f1lPqKxfUgfLKAOxHNURmZZ4FBD4uG0wJma/k0XR+nrmUxn+MtJNpm4N02EOPXOEP65+Ztsrac
zGQU/lI1EM3Nl17O0Ey+g3bvBD/NGywlJnhyl0bGb+FkQUJXIcE3LjsHxqXhVuN/sSN0dicRtfVK
PdFprMCF1gzOI1IjeamkEoYGCR7eKfz4ZDieOD9Yxw4a7ELZvDadOKBavBS4sLCrqmhFykL7zMuJ
eQ7/voJuq0KrAGlmX5wRbohFe1cCONUplyLwa/EapIySNnqUVQNb/EJ238jaN7A4At0kChbaNatN
sgfL4diSsE7LKKHeuTI/gEp6w89Cd5WnFKq46rKovGOn2P/uW0luToj/6ABVqzN1eGJCjrvDhpZL
6ZFM1dS9wZG9fx87s3cmOnzZT5QxQsZbpGrzVaIzuMsZ4EIF6cfjOJ2mg12FaFfEtSFYqaHmmAd+
NOmuNNVKxh9WHHgxdxx6KS6wXb1QKCTpr2GeeAH8QOrWZUPZX22yx3RVa+OndZpR8Z4H6OnqarSN
FHUHOlJpvL+t3JAfNeK4HPeKBeXkoZHXVl75Xri2QB5O1jmCP0RYyVF5QjRoZojI1pNJz7+zVrKn
p9PLkSCRdFaMQLJ8A61qDMfJ3yxPfAHDnccKOJQVY6JSVcwduA9OxrmSwfpkyAkG38KwJN4WFlv/
dLSJUxcLETt/sR64Zkp4TZVosKM1p1Aw0No3MUvUemsvL+4OBPYi4N7pQgAmlKxySyOdeSs0yg0s
SvdgPVgKdxoS8fxAk/C2jzzveRAx/cDpcRc8JaLAP1SO2AFt5u/Ld7OyRmGDn6KEyujUaD/JXUAW
HFvkonKjmxJwAmYiiG8F830cMH7Kuu95xya1/Eentll8/4oWNOre04PVLph78JFdSmohEElVdPuI
HF7lezzDQzkVidbXG2Z/JacrfLw5Szti7OnZCmffFsojUcSSLT+XP7hW1NlRSVHW6yekdGnNE6p3
Z+2LkcScB38rC7C+ArElxYcRBCxL1zmsNhah3eK/eZoEdRx15FltM1TtxuRQkggtHxpfPNs1fSoz
7ZO94nxlk92pSrhqqbDPGcRlAsO/oHaTf/6XUlSC0gBsHC0gMmJ5qYYh5hOk5AHm6Fv7xJ89vrw5
OEc7EYft1FbDYMZ9s4WlPgR2ahquW5Q/PHJhCNoJUszUGQUPSipLIf8m0HlQbOtStGkoMo7MVU2l
mZce8EMfbVuUUwNMvSi6dx8NTLjAQdhu196RFwuxC3dU4WCG/cUZCUAokvJX2blykog3WmNpzgtY
KcgboE7/rSbGREUeJoikN04jgiJVO9srBizu7+s4cr1/CHliDstAzD5i1GDpYytML3SzawPsAYwM
TfCY8lQeg0RuULYTkG5o/8xxQiKzov3zUoy/LTGNy7nVIVEm1eZzQfGy6mPnH/Dsin1AArQUUYbs
kkfzJz44ZVXQ5bBHp6SboCUUsh44dFXv3BL2WdqhmC6Kz8eUV0fgh7vcIGJmRrQjf7DgDJ0UDH/2
etKtKUc2gKpOWIpyRtyY7yqbZp5TdmlNqsUYLfKUyAKyzdHXSUFEySnKqgm/cl7T1vnapcxAQ7vW
tiUIKDRmmUPqEV+k0Q/ZbL0keIs68rF4Lhm0x29xB8JAp/vg3L8Uua8v8sLrBEm6IsvL2dj9dMxV
E8YroLQuie186QojVUGtuKkRCEHA203O05a7B8w7YzsaDJ5jZWTKGW+yp0JVhev2kHR4gcilv3Ha
4oxEhRyCKqonXpG3XLTig4oiXh4IBppfjvTymff+m7a2poy+1Kz6eBbKJP8Rc/JsyVCOgfSpbBmY
pjYHM0Du5v21lWCroebciarsLo9MwE/56Iyfv9y2AE+5QFcoiCetVYMz6DeFFUd1Z8Dj2YhQM23e
qNBxE4/r7/yF0KUSdXMsAGVzWt8kE1S9eALSV0Us3BdVsIKHx4sG4zDIsZBD2n7VgB9KFpAmNG0v
MNmjAWwMIIKoKyLuj7m3cYzHIe4w7zYljwPMlZ/u2vgN0tCPa6UK6HzHuqCfPXA1/LytuxI/mcJs
sPHvJY+1MZAg8v1wOgT7PBj6fBxdRDXiBf9LKkB+UcH+L3q4CMGr2uZv/+0RStw4D2Mxpe3z0fdA
fc3HPDKZetPZQ56SVwS7qTA3ByOjTQW95Byd4OSOQZQZvwnmOEEQdgH9+qt1yVtBaYdtvCIBUiNh
DmdZcYPwGL4VmMZOikD0PQl2j7Bv6tOKoEJHp7xFUNmPcec1fZR7Qgl8ImG7fTY8i5zm6Ic1XRab
8Pg8wM/BP9F9lxJ5MSWSgA7cats0eoorF4FjHlfecYxlfui2xtfonP4Eb66mggFVYRek8bGu7mi3
9vhosukX/8uUNZhyGWB94qpUKKtMpolP/rS43t8hdgl9YTBQjb00JzHx2skVnHnXRA4+UymBovOL
vM+aq/LYoGVHAClQUKuWEd/SxXZwlF3aNP8oA0QjUwZJk1Mgj3B0RpTqRflTkroHekclngBIBR6d
DJPeImyh3C5Y6iLiUCCtrPlhVxiQ6YnmSmRT1PxKvNuP0eefQAKWfdZT/Xr8gWJRm3oS/vz6NIka
jyT5H1zXBwbToFWhETXbXR38NxuXDDUr/uV9RVMd21UPXwU3ugpGeRfDl8JZdYRFIdrGqRN4zdBC
wWz1R1x71MK/knFstiJBlP3BxaZEmZzXzgWKR52da1ykQfChmmMw3u0V2e+cyT0XF6WVBOmqGXs/
PcHNeuve78zvrGQZsO74IWTjtlf1yPLF2/G6F518bPYmWEbjEKPdb3oJHW6Qwcadyl+T0ni6shu2
xkvjGjCx3J90D7G0Fk4M+VDoS5VM00Tpn9NgeFEVfha2nMcf36cngokpXf0mhgXeohm6NQmNvs5E
zoauyGUPpOIcG1P7gRWTdCWTTwHHMwDQ7aYEgLJv6TgB0tpE8idNg0i/TeImdfq2EmB9RO8xzGC7
ovJc+dQ+H7QlffpcNrmSDvZfby1x4Ic+iPSnSuVE4dNyYiqsICLP/HubtfXgbh7Ov4+/oMBwviKj
CN3jqq6BXoBLzhdVdsdEGv/2s9cYtBcfRxR4mIRimqgSjg7olP/PCGSuwihiEDR3VN6SM+9MWMzx
ZeVhIsg+adadXNG2IZniXbDXmRx46vMK47fx4tvyMGEA9H4IepanMckmxBUoz5cWdtkS5d7f84Ir
b13Wop+O6NpJIn6wGuGFx86REBxZ7/1rpx7oGiUIk8Mn1MAmOxZMH8NnwTqpfMZvOUVuRt84+r62
cyBsdhvhQ9kQ2XTdGWYoVVkwyaPByWS9pZX1o0vOA0lTyU3Gwiz7lCkO7dcRul/39za0MWmMODBD
CVBsM0ywGAn65FpM9NW//c5R2yis5pNkNDDt76LggQT/6mk39EidnG1LdT/FQT8fn5+khI1cgGkp
OOVst79Tum2ftLxMtFFU4CSRSP7Ifu9+FUtUYXwGerZEWFieeYPSyAw9WJ72Cw9U4h9LkAOn++6k
k8RWMa8mD42l/IFJineNUDkp4vtlVC3+ffBEvChXzS2XBtcBCmo8uuK8wIG8a4BdoBGnLjZlwjob
S993tLeHETWzz/QiJYCfXy8MKFvp0qb3r3TaaYz2rjwc6ccCxLVRn8saZ7Fil3Ne0f8Xq9xtxF9j
90buk3mTZq/DcAUEH66rvCP/eBQvlAC6mHWBTU9IxUdZrteQ0eujCyzPgWR2yQwrIydzHrI3mU+k
l1nilLPlhaAJfliHrtDEm60Mhw+ZTSty96jLyHgY3njazakGrJjtTHv0T6s4bvtRkHYJxQMsjNS8
Hi1uCt0gomc+OP8dIKW5zV1c1xy9PmxCdNvStk80+DXEmbz2xbovfiGrmZPisTK9yIxUXe6OODEl
zDb9t5fKBCSs5TqZAiq7BB3LPDo0r9OFGFEyKYO78uq2qeT96EpJAy/Ka3exLxcBLmR7MdgdPrVK
QobI93UkULeOqXfrsub07joU6Whbw8+ARaZQwDVyG0sIHdjz5ULYhfUfubms6tkbwrCJ31DTA6bE
jfMvn/LE7DtFW46ex9wGjTblhuLFLymiCOLrfzHzGRtYCqpkw0dp5Ioxq2bzq3A6r5chTDNT08+z
QYsrGwnzxqgPz76JpQ9wk+X5y8R/whsH3kH0zs5Bo+dtW37dXMXa6THupgqLy517u55OkfNJINFT
USSc2uNqhtssKiXBa4y3k3AFSc0j9Gl4pnFnCyItc6bTcNh67EdRQ14PoZzvfn1+6ank9m9jgrRc
cm+zYxa8XpTqPyAOk/j5qj5r7JU4M8mbATErdYHFrJWg48pMIKyF6KfUIL69nCgBdVDagx4Eg3LA
rzmAXYfGIoa3hFermhIT46XDYHU4bGE1Jyh3/cetdBHYJ2vmcoLSWMWVdv5zp2eYBKSuQfuW8SwQ
hAdiQ2fryI6JypsdM0WFrldqTEQ+S8ziuA7qGN2NH9Xv0xh1QWJx7RkdSLjOtBpWkyeDXezAB8ak
cl2RDHaa27osHrL33U4emGifbcpcMNZ5EF56ftiKsJHktBjSt5PyGAoHrftxhbbSLoVOmZVEWu2G
7FiAV7B8IMDqjrKs9o4tn0G4JxggxfEr8ewv1OQgaqMrHtHm91JUXIc2IDD1COFOiieL1V7eHULi
EqmNPPO0GCWVYwFiQ4Ji9HWhrG3pDPM3tc6Q6hiCcmCHtJdWDYjWmtGa6NQfo6+UYltO9iCncVsC
xYM8eLatPj2CTwLOgDSRhwDQ4eAG90RP+6+/c2Q93LS+xrFV9UXLzzyAMksDEQfgUtpi7AikQsqc
S2drsb6+oA70WDT1yxTcbgCJFpXXweoEyKRFG553QLI99/sdGsHywqJ7k7aplnXFVm6DeYxP46vz
0EifWtS4FHXB+xtodh83VhsLh3f3FxLzjiU5UkUk1GPX6PS/lRt4WBgFrTI3kYqM2krypxHxbLPX
B3ZbgjhqYvBk01n7L/+T+LnfmMdBlHuAZ+/kGOdQLVpELAE2UCT0yzQzoh4THv1oVbL86DYaDQle
JJ6UGbv2Rn+67dvlSltT7IikFzshP0gInvuaY02snJyw1QSQAfr82BstEe0iPjZ3GJVMbKsUv6cx
BJZU7U2KJHfTgqLj1jv+oX3FM6Q8vgDgC5eryHCtrTbWFqZLag7NchR7KJ0petDop7K4bSMnTg9X
GFc56R3ztanZqb9f2TujWIkRrgYkSFUxbfz9idmbl1wjEWuJUCaLtG4ioFwx11eh6SQ9DQCNNQQM
qwcDK/5h9ZB+LeAH45exy/ojniHZp5L6KuBurNCsunDKvh2hodzO2adfvoXRibQCFsOJkqgdiZTB
hniqGawI0nFHSiFTRgwOe6sT+bGKE2aOV2Q8E/EwBJ/vrgs/NYTuOTolshGeiVpPADCQo3v3E1sw
2ST/ZUBGtVfv6FTFpMcL+ym4Yw04O8DPbQdNZM1IuqDlNCoxkbH0D7RP/+xl9E/9pvEXfIhw6jH1
9gHi8qOBSgXLR+lPHX47JJJVpYHgYMtcTf8Gq6ODk0fZk1J+U7Nj/9UK8FPCnFHnxOW0c6hmbLX+
SAPLrXdJJwDobYFKIWs26pFx+IEZfLreo4lonURCZETk/6X3KdoHEQdBjGajNPPOj6uWxTxCy9EM
Ms0Xx0scvC+n0JGdEarOhxe9yC4CBLm1vCroscL05OcxhuYJaQ5V+fkEaCsJXoZ4vvOyRP+jX1qN
zBihXee0VkQk9MK6JuohmVK38ERZ7r11LeAIlY02cXg5YwRlfzZ1r91oRvxqMFzcQByq8jSbzra/
lZn/GBFf3WSixePpUPUpl5zxxt1PxCwQnoVezoxv2zR7SekkKXQEIBgCWcBAHL4bxKsVacM6N3kD
Hga5OboaOjvrlRWDwz81jChogJ28gbiE5bgKMo6sq0NnFRkyxuINOfdCEHAiYskwyCKY8hOwlZoQ
SJzgNsuOuVPrqyJQD0g3lpR+TuZeih1WikmhqWy1OkxApGQsIQPhJlOuKf34OUzsBHZOiT1FYFFj
YSIjNHteMEEiHkpKBsS8KpC+yDoQa5h8Zy2hYyyfrAqA6nssPVy7owBFiU6EMIRelDuDStIkuHys
tWqN8yt3tphrZruleWVzl3sKM1D/b0+SZprJuINRzu0QvcSoq2IeBN1rsqEu+bxYEz0h1xvrTxzF
xA7WlJYfVpJM/muWkXhqMfMuAwnxwypdxDlY+M6/fcbgesLl4pMe8+loOuHKBIrpKjD/F8sc9Sb4
16nO/j7K4wajM4g3xqSpGkgI/+d/PUxgMMCCngQX5mu1C3DAnh/TNlit4fb3nZihx8IVYSRpbX3E
ZEKWP2CMLDEP04KYytMK5bV1oDO/woiHr5PF4bCS0yQkTonSoJY5ooNoh32v1LPJQDDBaOuwcGWJ
bYXOIbr519Qp9q5U/e4k4bzEt3pFOscNL71OxdmR6eJ0Pn0PDFQlEJQVpCILQ+SicSNyteW0/mOX
x0DJ1h3myB+DFbAijw7AfwiC1V2I/U9j2m4iC3RNEoCPcsRO/dP77QGetz8eenrRrPKCfhtOnIKr
uE3t7/7qZOptZk1ZOh46iRkzg0UfxQvli4eQKY/Dg3PUQXytUow7kURfeZbptfA0s+URNz0t5b86
jZu9YCjwHkDSUGhybCuJq39tRB6mdEW80zC6/hkkEdMNZqJmUf8p4LKR+Mxn0wRyuJmL3qKedMUy
Q38FU1goBIhGPOFRkD9wirjkcvo94Pgts9GNDDtznZTEM9rojLif+gY0AI1Z5KlxsiVwR25KV9pT
NvrMUBaiiIv+Djs9mYnKkgjBVoq/d8GhhajabPwn1k0GwwfzviOUPHfepS1aVJPZ315ncGSopNoW
U3w5Wzgz9b4xv+ZgZZJ/lJnfvR1H4KaAeqdOeU5QIiB9U4z2r7vmoverwy2Lc21sR6N1JPXqMo7m
JsT4+DnaVVf35B9keFYkAgXVb/VkJGUQAmITrLGZ4YnZXyv6uOTkroxwVqWPkTJpoRxT7rsS0qq7
ZryKCF/Ky9kD/euK6MJMZ1mrwvQTgbrgWeciGhJKEC+TCuNI5gr8eaChohE1FiNVWW+YNRad6ZKk
aBS9lZIMfrW0YLchSjJUqzFDEWHEDjPNy9D8PXWBL0bd3E7qKkb01BeEachV0foBnjEPl7lKR0ro
airfJYYO4o1njdE/MEdyCvSgsDL9wOlhuYXWz3nqnfw2DoW6CwD6FEb7g3LJUMVxRN2bvlJEj6yQ
xNANwBLwgWE1nqd+PTBcE6RM48ENU2OSgceV2rNp0+Quj0I12kRu/TkOqUuoukUhijAhUMNwCNrQ
/yEsbrSOUZ5mG7LVi2PMalcAX3iEODwd4mtVI4a8P90Ni3Xx0dytEd75t9sVmY7PSf4VgMBNmaV1
ufTcIXwJqZNjqK0ymjVwHXpS+E6hoF7oQLbsciuJavFcquJ8APjg9AZmpwlO8SBSJIEBYno6XQRO
EtyoBPe5OwQNPNGw0ckPSxAZ43HRi7zlV+7VLlyeauPyO1e66Du+gawMoTJSqI9ivBcuO3h/JWWe
WvLRM4hdrZHmFEWwRqi+D7Vl67CSl1M0ISpmk1tujXT6KMXBsHlCozYqtvT5Y2mk3h/WuIL3noSu
aFDGk4fmGBMzaEzPjJQYBzoBI+u7hkU9ici14CM4/3mcYHPl4fS0L15dYzFxAIFSXN6Z9yDjCu2Y
SoT/yt2U/fXIxd+CNnyO4eYGiBEMgmOiVKYtPkx+nZQifLlgqk/PYTs5oOTq7fTiuMoK7g0yO8V5
eQBisXQG9dJFgdL3ydvj1vHZiLWyyKGacm5XHh94xpESzXnWVh/Fvx7FJwzJZEbgivRQDrHfgpbV
ymmqzwDeICGzwaeOUqB04MCpfFniDfsHB7powCchf60E1d2NSOFAbV1AUwbF7UjeH2LonVSe0mcK
wF4bglNZm2gtUQYVpCen56KcrgCKiKGXOZp7/TBla19CX1ki7Pa8+KgyffSMYgic78RtOGzMKGGa
LOCRayIW7Vglpt2V9EyvKeWQzxxPT9b2KDgu/NrIhzjY5x7zuogBhbsxozPRvQuMXJZ0Zs2Lp726
rZMm04dUPwEoJRPMdlyLS5d9Ts3h3MnFBJS+B8wIMEQIwrmMMLcXGgMMqAF4t279VjgIjCyWS0zg
MWV70lP/yrUIOtmATpyaecPHtY8RBGg2aTUnxLp3Igq21pJAPYCMsU4Rm1qukY4L82BRZAu/dPqg
zbbHNjPMSd3Fnx+6AEQP3NGok6DZlSs5WUZ/J8W2nEM0CnpEEQSYBBD6TKW0EMh5O/vfa5tFr5vy
7LhDo9eR4S2YN61ByvLJ/yS1MvO/4dv3lLYDDDGIwkaeGGOOO4nrf9hLCdcASHgCEC8SCkYl9J/9
oY95qUkNzTnvnJ5dTOSVNLwepbYRk9OpxBVThwQKf4gzAreg3Wwytyi0p2OmUUXryGUnu3Y+aEWG
Azl/DSJ0Ot3ATk0KN6EUNFoI1ZhTTDRniNpsoh/XtcqMH1FTC1SJhplZMWnm7W1p2E2fVF1Kf6lo
lB/bM66gg4lUbPY4ztK9sPDz2pHEpoY9lgnk7SZ5ACZl0vodY9aH2rej9QvTBz04Dp9LH/nf4KNs
xgEBqWzftAgEemFrBQWZpMlMJ2WKkgKteiiIu3ffYILEaw4sZYIaK8pa0XPLC1xoFAQwBGbjUpMn
ffzxTDX+DuN+bofCj3jFyyuESot0HuxelhffZLn48OJYHnKKWQsoNZzx0dDmz07bJy2dB2aFkL27
7wuu9CXL3ZHIE6N7shbwuefEXHRUmXba3ZTjGy7ta0MuBRCLQKt7yWEk8CmwYXbnDB9wQInDNVc6
qpetRICndvhD4qDju6oLMMpLFdhnmpSutOPZwsbsjlD5lntee+qNxkVGftbO5skTK4h2rccjvBLQ
SYL3YdRwjehEhjkr4kYstPYLrPSFdZN6TECBhD/prjbPwNwzG0uPsfYfh2D5y3r9YnMXOZK2pxHc
xxPkmZcoy4/s4LclZqi5o2UB1KWX/H2MOUumaLxDjUrjEBpgm7NtFLJpApsZA7/+t0nNxAQi/Pco
8pIRl1Ts4GlE3kHf0TI/vhJNKoakHOar6yTpBvaqzhYIfM9qKRz41OIW6uP5cIApmFGg6UvPGrPf
aboIFh13RlH+hBd3LnafCGcvNd8gctjgNKlegk+qftBsrvKrPKmJJW62GOp+xvHe91HA/5uMSDjT
8/cOcTOPNVEf2NrArr3F4NXSzHazqX1/zZEavzCdLi23GHm05Wxl1PiHhyTn84puQGl1z+WrOKlZ
GsVeLN69mJ3WBHQHiMORo3vkQFX4wAS8iMwfQ/9shdbr3vtnTsM8F9YAgVAhghLENhsz6AqUZIlI
iVQM0QaJBiZnvvYE1wDnMnY/ui0DSoo3i6YJ+9oVEGcPMRg2h2N60IFQ1/L2aq54uS+6atYKeAzM
4M0mo2flX9DpF9BdH6s4HTRxOOKJk/CaRY0s0f8mhzh6GVEqj/gvysPO4hmGJFdOoESdO+AqKtJw
pRIDeJgwuNtnjI9JGYCKyfSGrz2c/ErdkCNN94rJ69cPbulzT8suQ7GV8cNcr9xAnbNT0eSItVje
YQPKUUeZdmRK8gYwqhCqF9J/YxexyzC+Fx3sZZlfIr2AY6ESuB2ix9y83i0n2/0d+KSBtPlhKqYc
aqa6BSWYKOo7qBFTwJ16YrM1nd7bsPONtTt+kzG0TalQQ1j3dIWF5W3XncPx/lDAychm7TrEXY2H
GYAL+0RQyASOqZj6ZI4Djmzp+FxoSUTUDfST6Gs6plhybafVTlb85InyWc6OGj0gD+4l8a/QCJAn
+muyQizOmMHmfNLyp2CCvLN7BN8xDH3mTmeKG4j9v/teUS1BNYBm6d/3ZPnDMQth1y+Bat7Vr4SU
uZU9uU+DZsPBh79qqOv99Wg//1UhX8f6OtZWyHhB0k63IGcrvhDpnGB1qn8i1LqpVQXTs+1/cdXJ
GOuaedATNKeY6GOztaipLtX+qDsGZLgt80Mdco6AaSvEn6GOBqcryspsQIHJ0P/tYNk10zxSi3zt
D5m8cmKXTAQitm1kGdPrF6f9fcrr8Rb9uox9QxMSWGKIDkhRCAXSUz0NJo+rL6W6R9cyg92cyBri
BfXOk7zC6NgcEq9DnwgWY++hUCEByzMRoA4wHkIZf/Iej7f9AoA1lxZKDQQyYq1JJAm09AeyiFpq
hKlY3KNv1/oSv3hO7rqVL2m2HSCpvKjjZLECX72runhT4aZnH6pBEW5/Ro6NaKP0MKUuucmmifmA
gRilu3hrwVJEzFNAKHSyDlAXCGtR8X16vjOI0VMYg9PhFL3l8FzabynVP3ygRn3ILmL93f/D64Dq
FF1pf8kJYYAc89tmFgTVUCclD0k5fszvG34xzfkeeGF5Ohdz1J6F0E/CgIGNkezIYxOR8ZTzAMRY
NPn7b678U0ZCHxx35j0ktRk5wxbNQZeLL5Pach91nTUwzJBp13mw6QS5E3Ud/ngqfYM3AhTRlwnz
ABQGCcsJaf0aclmG+u3jkDTcsHrBp8wSz4jn7euPlCqIpX+2HATF8Z+jFoSlDT99AE0zHsOBaj0x
Gr+JmoroE0PYyG6SuCBBQNDEcAJ7keR5e6lxEpIHPDOp9y2mHmkwlRARaDgWq7olO8FCW9+++7M6
NQhzevNsNVWf5u5kTQ9U7/0EAoG+JBHktEHHX0T66MQRjwcxYeer9x94yVZrStu9R4goyDIgrcZ5
rijicixILI4Q2mdiGEZ2abNRy6LiPSZMFiMTfziTKcnC+vLJJjhdstW9Zd0E8fR7FJk+PPYWeFve
kNEfKaVQiNkavvUMdtvys/K20mg92L0AVi0MduimVmLr084PlSNUyi+NLi8Qw4JVQ6pIAe32l+e3
TVvnb4qFTLjfPAKpuXAUtYssl5nm4ZFwJJztTgaHf/I19s9KIWujpNVNfP6mRx95ahJs9VEv/+9w
WwyPWKDCr52w1T3tguTjdGah6+Rv8SfrXv2QqRLQqjdMiKvPjX43lRXvaRRahxPprulDjRUhsQO0
h/YRu/SUOFUVLjihotsTmo/SGuqqynE0PobcPIzZrKPZP1FtdgXw2DpwzHdGerl+6peYx2XPUv7z
AH/UFI/IulQRzpplK+GHZXifu30yANLNWSpP3CntddVM09mR4Pb/ornvS2kV05AEvQo+oojClffe
ryzK2XvYP1/g4X7LdOhjc5ADTdThdhWv+hhHonehSY7AOanaaFJ907geerHqxwP5MaQPZwfAqaxE
CumYV2b9prk++YCk4aMclWx78TP7QW0BsuW/Ht+CDzly6UUObl9rydkRctfYH7BYQmydqPiAHuvw
3pKDPoctzTDNKNiWEVnXz43UswhgaxSBN/S2pDgj0HYg7dfCNIrltHlVUA6t/j/jD6r9YHbx1HSM
ZMQHA/OWws9UHjfIdDKwewmtv8HUyVDYjvXcvych8PrkadaNLo74oHYhPJ1+nGP0SRDw0/LbuUlg
DnCpwAA2AswbX+Efeqp6B4oixAjXekqovixTD5/asux6CyQdjB0YM0IZs5d5U5rNAxTLlug3AQ3l
KbIeIkmpwrKKTbAc0de0TZtio6D2ZBxrwjuurraZZmXXHViXEQyDYrM06HXG+4yVpnFIyKyqeTTs
c0j3lSC1qVHxM7zs3A9qaFsLPkOpOMZMF0FpYligRDT7KpPfo0wzVYsNQ/oaqDvZJJEBBCPVQCL0
zy1f57NHFHJqzBfnz/Q8Oma3NK2BRdhKVACYjPp9hQz6OWo7NSKJsfJ1xqLrcck8Oi0JWxzbO20P
MxKOo1HMiuQjkn66cM+KC2ZtEK/IU8kkx04O2C/WOcGbOgsHYRXex/IrNkId8px0rnQybg5OwTS1
i4Hwc2pN3MjAJEzFQ+9coHmtvdfFs4XuYuawwLeUNvHcfXX+zFL/uhJplSSlvFUV04D/UZabdfur
mwkf+GgOGWSyUnB3EadfODqOOq732lJMv7RCmh+2bgSXwv0QES6p15EH994q6mJzUbi7GyyrWb9m
bH13JdD1YNIN4bJQTz8Hgfy2mwa9NL9IBNGpDYx3oRS+j2h2WwfNXQVHqX8Ypfeidl0kKyDhwHmh
dO1X5Wp7XUKmQUrPvptQFbq6SDLS02Ff2btvD3bco9BZy4iQfkxZYB3lSU3r4hXWGIsSMY7grSjn
SRq7Aoqt9dCLT6tQrm2aIKHOFVcPoPb1FHMn13KWSGtha1Bgu5Su66ToOWei9+R6tsSLHGcXz+Js
pBPrSGWIrqnGWKEF3WX3rqiLPkhXq3PN2GRDx6xIxPHklzyc1L/pNM35zW+uXhayeoa3AY+BZSB/
jSHwhi2yeaSMdqx1ppiZWTssBs+OaVSueJd2A0Ml8VgUU4AiEYpYhE/mkuXqyhd8VgTYm5udGSCF
6249rtKYhcOWXrER/8N77DeZNnDNJcEu0amYPv1eBZ4al78/S7aqx9bdJXS01pqII1G+ZTWRPhly
3xdlVvwB+Vked9l0mX9ejn17sxpBuKqgGAGRnxvSMntVNSFVy4pc4fySMSsc6MWh7i/NfyP5QPRu
XBX2uT/XsrXjtiK2DXloOYtXiMI09xJYndD2gGA88SghfgOapYO0VZrH+nSAfLDz/Mr92wNgkvZS
2KMnoOtT9Iaa8NKHxtMYCyzGGfavbFidpMLfkzLoeuZ6NOIdwhbBXm9SILYSM4ei1pactc+KzT1w
6W8z+BRmnKb6eaSM2gb3RbpT9Qbvui5eUzNFWkJCpd0Dr0008QPT4qV4ZNMPyyLSJYvQUo5E7aic
3FhVup05U/kSAf+smHbpZ9F7KPAL+majCpEg3haKWBj+zsbVknkhf7Wp2xOUWYHlfZg2yU3jSHGP
5nhUpLfcmAF9QtvYXSx2JvWWcVnmNCcLaNAYrBCIbJZMQUbAb9eXD9jW//kPwWVzgRu3PFnRXal1
+bcfY7zvEzhgGfuXQ4ohnBr64aJyz0bHzTwDhK20+NcLAzVLgRtbS2Z9YLeZ4uiApk+wEnAbPA0f
gZ3hFtwWbeVmRLXLU5dHiZQ4KdsLRedFThaHC+47kyHNAOL1IGBDWXowc54jsDxuplMH26aTTKrD
nhykfi3j3jfd11YdLPftm3WqjK7BHeemThmzZ4clLdRiL+f6r+y08azKWC856N6/FzXQq06K4iaB
cAwEgMrc1VnNMdUmw9XPHJ5J18UYKH4ofvfCThsdY4M2GYtFpkJ1cCU8cK24FaqF5j886eIR+W5g
ipxtRG9wclY3ixqGHAfv3omF6bHs8g42NoSClp3lmSuiGaWwHGZtSnEPIox5BB8RcrQSh37n1tPQ
VwbY1NKgJXW/h8+33CivIhw9qNncjnXyK9ZKt9pwb4/vWJ4h6fBDD95Y70X+PfCWwdYYpzTqOQh1
B24k9eTPZdChAYSd3ATAnmcbd23t/IYLxUMs8GIzr9NrzisWXHsh2wfteD2gxzcKjqDN2EdWAd9o
sv8s0Ob7AL0yeJKw/G5Gn7LP2XodpDmeK+zPEYGai6ZvP6nxsaN2VvNpQZZsaYqR9POZKjttb7uu
6Pk24CptyeNXVuK0Wic9Oztx37m8QY0DZrYax98FwexX4+sFLJ150XzIep1xz4RdY+sCkx52b5xY
PankMLjYhjIYTwfF3Sl0l0F8ZkF2PZ0SCbk9vbLxPNCbfTXkgRaAFQc3hHrM/5CTDQD05NL1mFPw
0WHtQIX3As9rVrQYMJlqibjKddUl/X94kCz5jxtK245Y7Cxp0Wx/kehYkAmW3CO0t8yPI+V1iv5n
lLkwJys7sIIzf/haL7fSg2P9YVar9Gxwgqzi/GytprsiDX/8hlECAMmdQEwpbR2aOLofA7Xbfh+S
nqUFuc05QQzEeyMKfdOPAQYPqec44F6olMoEt/B+AEXRAO5Quqfzi2VOUE7vv2aDvZK1Mu8PsOu4
SKovfSNSkg8TN0j8QfALIXN1hUlkhlnXBEgzdN/FPCJxGNOXhqHd2kG7f2+uNty32n7FMace3Zpj
Ot5chk13lb2sGF6xXLrNGq7v++k/+chuiCt9BqpZwoSMtCF05XvLUH2zO1/O3UdkSGBPg5u5o3GM
z0Os5rA+4zjaT91bG7DcA9DIS45xzH99SehCN91JYjxcT5e6lGK2DwUnrFx3Ql6yhYlC49z1qX1G
Qn01TlFvo8Qm8VNcIN8hUvOotKXyTwzAaxCLFZpbFDPu4IO1TBlt8v/1ex0BBA51S0RCW3/2jrhs
JJ6lXeYyIFRtM08QekRE74mp90TbVo65A4mxxhKBZodXHIHCOnWBuu2/RZt6guzaWpI6VJVYsYXx
LKUkCLqQxUxYriMWVq8Sq9fGCq4hsEGeIAqUFjjo1h5ysLu1dtlADRuGCIL0KAu8dcbSC+PnXdLC
HfB9Ye8UqNUxiH+N1lP13AVJ03loPoQiibleBbQv0wothh7A/z1FowSTDSyJQjuCc0h0hto7ANkK
GMkJ+eenUIDHc+ZKOArNwkbUMojhYLdBLmuZZVFA2crDLbd3xe5WMROT8TQMBzI5X5kKx6femLyx
thyYt0g6qkH3Ri8v/bDX7xBD94+DEID2hqXP+pzD6GG/0OuMPT/qi/TBWxxBiK0+6xjPnUgkVO/b
Sccjb4bZuQMiwJ6US2T4thUnpHuDbmGDpFU/a+X+1j5bY4GzAQ3e5Zk1JT5b6pGwMTVcZKnY3aO6
ZWhpOMWovi2SX9rY8z9S+pdUvaXheFArgo1jvSXwwCtbmBkz/aASZdZCyduBBVnIyWTbzYpKILPl
2/fwJUK4+3M5aLOwO9hVTp8o7C0aI/gZKNeOJMpLGZmPldnwPZmBA6tH2cUhouK9FZ76pfFEeXZN
/KigGHbv+pF/YhUxGQrbaWOeKaGm2a1yBU90mjwNC+R7q5OHuq8ax7My8Jvy5loZcxsdQ5e5pBQ8
5C7q6+zAWzdOz26T7x98cAyAYd8QSd4nmCGuf57NA1btRlsNN4WEoUNchzKVLfokxs12kVgWAs8q
W8zJ/D9bkhBTH7HjqJ/mVLxv57y8Bt2wPp/ETSz7SpCSik9UQQzDeMELCuxqQcowdV5zkQM9FVNs
lunFASvMvCCCy6qXJ8Pkd+TOcHfONwfzSZslUZZg5QIA363SeInydeyfKNtNxO3LVe4GakA7rqR5
gXwphZc1l3TsNWvVcuvLf30FdTvVMiJopscuM1Mv4vCyZvfDduda3+TR8Juos3eUCG4odthq4E+z
zYpuKZYYEBd8slBts7siebMTScQ3hw0UrriOhT5IXr3RJSHOY1tkU+3/Nccm/qPVaGmc30Hq2Vt9
8oI9ZmPPKgiFZGaJ+X4eEDh8p0TvKV62kXVPlddYHtdRLsd9MtRJbh9oldyteCy4BD5ywrHAb2v6
q068i/R/Ffx/ecIybMHk3L3RPuMtJQ51ScxwNZ+8Ho+4GQl6BdZ7LFy+HsmOohwng+9LFCQCeaDg
LusSqWJSUhu7Or+ChtmIvb9t+WxWxQx6PkhqGmZrH1koh9WCVqOq55IwnO0QBJk3mOu1jJ8L7tXK
XegzVP/8S7demP+L1i4XuHAssEjYcQBFovNAUOfEfwJYWGZh9Z9azfU+2Ddy6tGEqmOMO+h8d/YX
jhAj4BAY4JhdPG4aFqfpTwfRmfTFPW/UgETG8WYjLRBIHAYQusoZ817e1s0/vphduKJMfQ8T/b98
E/fENyk0c2VaJKs7DDVBRducjtcGwn7STDMQzvolwuJRm82qVh+t1PnUR3oSwDAOcnXiZyhD/e0h
114v2yfHh6HEL35WDbf7uhctyX0K5MBHPaSH5fitsRIzDd0EjcgSUojeK7tJQ1BiQmP7zlOpVHmE
E7ZXActkbHJ+VnFVqUJqyo0FA+NTvA/j2w2XnxF/qjuG8qAehONshwS6U+HTR1mAUQYFoSWmtcpm
9lmgHqy14yHbmd54cyQU1dv6+OpT8H3qBN7xEG/p0Ig8k5IED9uGk+H5WXmPyBFjBmDnHKxuzSRV
hoqJQIoaFMn1FQq8UizJ9hL9xoFaJg7sH+Eh8o1LguS1jYDGxy3mVi9yeURx0SbAgb5hQlwKk+Wo
okV4OZtKjMcSC/rA5CDrOTSGenQxnGU4nMBriW8s8AGbx/2OyBhX4o2Jj204LO3lWL4EPJz/UaKh
3rptbcFy8FeQlu+TWqBQ9NAEGW+txH05XI5aM230YNogFP7nioBRDzA+Mk2e/umBejZzgkrlRNBo
jfMzDOZUkLZKC98J2ocP40z7EWVnlWmLtriRLBgDLt6PkRzsOxk1wh5bW92F2aViH7/qi4dfwE66
ldE1UMdfow0QkCmyo6REY6GhGuyHL8P9Z4yms8AkomaN1s8XHg+z4P5C+mor2CaHfbTlMnRn4/pp
uO3HhPyTntiGooMpIUIUJQufJLEVNNKBPtBbpsk0h/94j2JgwoBOqE1flU757SAgtye1DxBagnrg
BoPJsEEwXkzl6kf+8Xlm1zM8vyQfM6Gy7J20Z+5vVJV9K9mbICmctxSyWV7z39YIuWmRZOM8HI/I
nTHPAuefCsStNSxLsUKF8632bhw/rHgREt9QkgiH/+CJV8FOFYrYDHuJq6nGkwA/70Litb7Iitgv
6t0N9Q9tZufGWJt8VhyYTLYYErLWmuYbJBeH10gO40q4A9A23q1P1cQqrnST+sFhYW5kirbTT9Pi
J48mEAmgP+Yt9GxbGaDd0KUTe051Enu3bqEd4IkcFn5pyj7foOolqCb1teSNg4UhcOVmExiDmk5I
qxZB5LX4g3fiMBkXq9tNNGEXaD2jWaUzOA+RwbUWptN4I8J+tuel96ts1XJF0oj2xUKpr63++62+
iSLAQBCAM/+IsqSF7vpIw7NY5Ljs8Sqtr7r+p2rQ1SBimX5hz6418yLARSBe9hAbMzz9Nz0qdYX+
GlJ8hoi13IHFRAPmCtxfHJDoOE2ktyMIIt02kxF6hNFpeTHOmQ7pRMbFT7fFKGtsQm1hh9uWZuKS
ASqvF9CI3/Pkthqt9M6D52VHS93gdgoJSec519qqjtrfsBq5N1IE1k9A+t/mgCoEEi8mqxjwTzir
rc2/25tWyZtikUpb71MiBY6aYsKGw2onhSiiO2LojAmCJPmJhlmVA9uNOwU+gj/KWzhJkw8TZ50o
WJd0IZ8/lTtCjMzB2gla53RYVtmEVdXwjPdeC/kHPx+NPPCRB+A7jVGwpjP1Q2w1GYQO4yBH4Q4X
Hth8qaXYRzLzEeHVCJVLv/gWLW7NkUcM+B2gon7ZH9dZeF16kS+1749p4h01BCkqTNy9xBsDr1Lr
HxkjmgqaM1T+jTzumoD7QzWmANlw39/taoXlxAyWdT5SFInP5yZJ7MiZMBIY4QFy2nu3W+3akQQV
OjDTK+B6p+ZYHh7fvs+GdZuBRTd12TseJ0DJ7HcsWIKEIQJRhfQ0GaqtXA63eNdjnm0vVwzaGPNl
sb6E4n1vbckw0kkkhvX/HTEl/H4TSYqQS/Ys15I6uf7ZcMDcUbTBY8kW3gtIENZDp4rQi+dhIZLR
IoykV4J/mjkYt5lynHAkFhYN7B7DonKNEXIB76PA7EoZuFAv6NSW4p53SIYgHdJoPVmiVcRN2bwj
5RCD3n6Tjoo4q9l8c8QeQtgAmJO/67lLA/LO+8ac2xdIVvjxYowhU5rOJ/7mxNQ4r68zz47xEck+
pkZAmwIhlHsY4P7T1FY5JUJBftzCSgLclh/rIa5dwMM4aA78q3fM5u1gIlP/uARpygmCjrTXwjeZ
+pccqnUQJK9RO3cdnqsbWL2TNF9COfYSIjDHfNlp3j9uCcS314TDLthD3BtooFIOGx+cp84uLpv8
q6q7BQBs+BwHtD6ysAh+CR2gINVGqeeVhkvgHf8pWaDNxfGMOxBv1+VPOxRlEmXc6sPsSXB7rgIs
MV0MyzbequDgIMvOVafdaK5Ia6CnAbzPKbSQqFwEZ6q3+74DI5pvkGEfIh4F7h7GjoWuUdbt/AT4
3hL/vyymXpBk3ZKYXpsWWCcf2SWOH2IqWXdw7NHOR9u3in1ZjjfQNBVJYn3qwRtg+CpZa3zu8h9T
FsjTy++2rWDheyGlNFQLFxWvf4qt96cKtjGLZc2b7DTvwo3UQ5YygiLNXixzrnLANk8qK2+fjqKs
/oGa+62dZNrGceor2BAjdtG4wm+utpr/6Jf07dBPZOMa2CBADFk8BRQL367wQP8SpPlw9tB6bKZ3
P3KzDP3bMePK9tZc2Ip3SO+gVrq7nkVbFuF7vn0o7mMV9xU8MwMldo2tG3j0hJaXJtb+u2CTL0t+
Rhr5ccvOUf/XeV025HX91Emc9rNSelCjRDpRnLnf5kCP8vPqUI7t7dJAAzfYp8hjrrhUFd/qFC4a
QlKtaAIHcVFEwu9euSY6Mo/1Z1v+8fL/qDiXC8xRVuxqrqqb4eejLnXY1mOtlI27Wg0va3cKd934
pvSlLLl4kX7vAWnHbnSyzdDlLp7l9mGSNws/E3u8xefL4bXOZRqZQCad2oXfgQQuOO2zhT/4lfZI
xYgxsDFW9S1p3qJoDcJnCA+IpnT80RTjKC7zs22ij4ri8IJxs5GgNV7BaGBFXxEV5tDGzjffQEk3
CMC8FG5SmtyADyWGBAwGVIhKvl14+qwzb/QPvvCx9TrlI6e9Xndtk3iGp1b5CagQkDam0Vo8XWD5
qz5Pw/GgB4nSqK1CVYuUFlBwjXn0Mr6AksSIMtR3xltU0dEbscj4GX0Fn9ZRS4HfiGMpcYfnLJEz
G8BDZmFXCePGc05KYVDYZAyeUlxxJ+CZ+JFtMGOjE1VN4Fw7wPvk9Z8qMH6W3Y9OjNnyMRzIeLko
wZe9U/9NKhFrjXhqfsV+5/xBltBdxJ2WiNF9OBUMZ0dPsxntzYjLOr1dF16TsIIC2IHrMW4Z1cUY
fKVzzGG4OLuE0no2UfFJrbHia4KzU+lqMnVPjJmoWJLn0Jd9Sf2ZQs9pl3EscmgYJ6fut4/P9iHi
h6lkn1YOi9jOxNj95N6UtTyc6qw7mCengWGx9b6jN9vCAYhk4ytdTVe81+XehFQpP2xzuGmVXsJw
5OQEiKJ9RceOe/uZqLwkypvx6vJwtNofMHBs3BrIJWRbsuZ1mv3TbPrAJYdU0oHCsTTGObqfyog4
6nbHhXXNBlj8Tm117ZuKFLfUaGk1Yv1S8fkyPUr6w6ZIOL7lOjx9rkhxlbX+SHFHGmdJU+qata91
OJnR/umX2s7MYxHtmvZ/b4gspz4jipPpoWMJwN5QYlwPBC+nEB3DDbkSrXg0QmBoX0wwGwj9/94R
SQErBpZaOeyQoDpP6ZFPdWON9kAzTXMuexgF/pu83a3tyFTbyqofnOg6xjfJKUBnen+XZSN2qtYZ
dcX6kluMBXUlu4icVL4ReahZmOEwrXAxjK5utcQ4UiSXHatnfigA7TEH7Y6ogzdAQ7JyWUQ5S6zA
Km3QOce4OXnZ5lN6ewmgr5HPUaAwFjSoloikXxl1ChJcojVy5Ufyvdgv6zrpVukVm9rWlDtaMJQu
OrTanzJ7InOiAmJW+kxRSGB4j7p1QtJsZ7Sa64x2RNCdMoyoqeQawHAfeN24uRaJ6Xc9ANnHnKYN
jayCKqqWU+eEHYyWlFWtaRxeQGasZ53iwZoTPrSb95uovm1xVAwFfNJTN1WttptF07dHDpNsvcqR
ZN8mxYPufHFHPlVCqaMbiWiNLqEfXmVW4FUD7/Y0dt7Cph0yvg2PbwI5V7rdsVNrnGsEUQ584NNL
VKgDsZdOU4k51YaRs8Zn+fwKq6TjViCLgAhRxPiiFCYvO4Nj2YXTFeC8qQyG1ChgUfnIl571pRYK
1kwQy76UkCd5CWyMZyL0kEHnX5uUM5DzJZu8mcUqN/Cdy1nCBhKELpcOXhz8LoxSeNkjRfNcQaHh
JbaK5IeJWxlaMAWYXWWYtUhXEMlzqZgmTCWL50yTLd8iwidgzoKFaR0SdeCI4sRHVcR+oXY+upO1
J69uvipuCpMHL27kStHVpRu+E2D/ednq2/854zxw50Vq83L1mUMO+eN210bhs3Ps0N7D1TyO5DLt
7AbLnz5ULeGxHvXlYbfPzAT18/YmzqLCTIFtc6iOv5uo8WQTPNNY+QtUYKjcpruC3OLKTW6Sb26h
id0QEtv/uUCtPg7Qc2Lyf42lmy7qFzzsUWX+guFZjmfv0mtZvlOtDGmktFetYmGtcQmV3vJCpz6X
gTXedlxhmu78aYHHKiccC4yFMmhq0y1IUDMLbZKfR8cJq0MkyU+DrpYIjlLfYmJpDjHINQ2Wgkfz
AVC0mIE/EOpno/K5ygXxvqMsFVRRw+ghZA4wTH/bxlrNJZvCyCmFEcjh95bd0VZSDSLJ3z9ArwYl
DBsmzIQW7LVTIxvdW7omORrGHgyucAXNeH9GhGd/rPlDKfEKzX9DFTh43ECJlQGbyhtRJJgHXU1M
T5KANjkGLZubllCXhE22QYJGpX1eC6pv2QopTOZitvdChwsb+nwtsHqWxztxaElu6l6uhZWJVpQM
NPBYT98QfjQeNvO6tYyTVa5ltccBfDGr7LGIS6XQWIARlxBl86Wth0ctq1t0o6/Vpvr9gr/2Zlcq
Gwkafl+MResEHQ2t3TpOZbJhj1IwjJ9nvFPNX4W4uBiKrO86FuBK8af4WQqrWy3n6Rm4/f2IgQ/x
CCJH7ugE5LcxZiJ2nmDUWNX5HnjCs5UFCS88kR+Omv4dX/pQ4YoBdmNAAJUgoZYemNklGbqlHRle
61feGacctFqhkGFEEMKJtXBwaJCQ3pHGeJvnGUy9XeQykCwaVvlp3tYPJYToybzGv26/Vp1FV66x
UpS5UL5LQvRopq1DuagzvroW2Szb+01l3OfgzR+hNFRl5EiiLpZraVZwMPCcFXp4onphvwfpG7BJ
cAbdO+ChAXIKvIzo6kcksBXvXfuaKsQh6BmWhUMDTRLbqyBC4YEROr0aNM3Iyf0iLAjWM66baiMx
gggypNpKDzs94QzN00LbzBbKke1PnclDTvtlT7phOKMWikvl0Ba1M7BSdU5FMLflkKUvIMY44ovm
rhXHc+d1ga/1pRGfYSIbLpFl9FnedZ5nmrI4EdIRsXAiNU+r1iJ980sbX63aWRYdQe7/fj50ucgH
RhksEVYGZC/gpmQT3N0AV/+6eMbvGRCV18hjco4T/61C8IKHqY1JNesInBhPJE0xRY4YH4neNI7X
HRCwU/BLEnpi1a9LevJNQ7q5vHx9kp+PrPqFJuClRywW7XN306weXoqqAQKD+ifHNsEhlkntBKxG
8VueDQNGeNlBj025p0m016REmEX6VxDuwd1Z3QdQ3Zs0OffAaj9D1yjudyB6xdHB39ti8p6ACLas
xkVmgAcjfyJJJE3kdl/lrmN6mR2knPCgJAfoIAXtMYGeqf5+AmubAUNqJc8XdCViQaYKyPGQ8gvK
EYZdc3hxbpzIzOOuVWBIDjqzeEG0W+GsrSypRRcAwvXAY3Zxxnk9XW3xZj9IuHQwSUWHg9cq9Q6B
r4v4s3zWrVkfG7zY77r3KZ+eVZ5CCIStLixLn3gqmB1IC1Kk1DUMbqQYXQxgM4gyv8fTbkZU7vgP
9HLRLrnFVfvliGxK2CpX3/pEy0qY9AK5Rtz68TgJBWy455qzqQrxFgwj9hdyHJMuSLbORvctWw4B
t0UulKt/gFyvYksCWZRPGe+3SeF2NJhFMjIlUfvmEb7Q4eiEgYjEcar584/PiTQ7B3J8l8Sr1ny+
3bEJ5RzihnzpjlTED6LDwu0+2xQ8vn2JJqsXN0xekk/JEtYBL7sK5hZ7kDPtRo7+M4U4XRpwc+cI
ziUE7JD1j6pNYxHxpqFaHAZ2WUTL6FzMrFcerCjkRLDbEK8nE10G2ayqZAw9wtGfMXpj4D5y2Mir
wVJJiPr6NarFJV8AgqNR7XzCMZFaCrDRjxCXnOtloo49nW7f/FN7+Jb/BQny9BJ/e6QLypFqmO2l
baURUGKx/z2HAt9ccZvk8ne2HkUxPYg7kWZlKtIFARF+2Xly9R+k5LKHg/iY+WXHHH7s3xqnMTew
PqWxc6ZhjTCYJ99LuOJuiUxMfqzMd6QtoMYhSDmzCCn1OORKcUfRw88DQSAxTuAB9dC9yQkUdmtd
rK3gksiQCJdN73zhjKAWtrCFLjPAQPQf4LL+Zh2B2xeIeV50o3TktnYLTJ5vO6qIGvyGZxXZJoZN
l50xmU6ASBwOKLgZuQRFOfjXNYrkiYv09BZff1SP/luTvfpcHztLxC7tVXGc0DNSeA2mL9oxxMl/
jkhnCigSA8w58iwPMD2nYE8oHAslfxh8eTtqS7dEt6yqMYyOopxIoW4c3dMBb41ivvtpkKy5qXV/
igwqd3Xt5By1j3MYtstGHYXWVg6gii/fKb5pPrwyqQJJfMbjvKVoeuoDJ+i6ZlQaS+dkdb/ZdrrG
OiXgSKCf/Ox8vYqUYx/ZnS/X8Pvh1ZEWhj8wlM84Sp+weia9jMIup5DKo/wfeLfOp/uMzSR6Y6gw
WTNbx5e0TKS1CLDV0gKOl6Dyk8KISBDP9ln7KGn+NwjUryQiybM/K/KT2vZSgjm+JkMywaqojAaZ
FFStaJ7lIzO3omSq1x5m3OKlk1lgrFRCbAQtYLpyAa1H9LCA9kX43V2GcjFyEw1KOuzUVyzPdyRt
aS/krdW+PDff07OyZtRZML6U+PSm93THpNOtVsiUk/U8h0x4SWnc0Wim8npLCkdcUmx5Jo3lQ+DY
JMP76wIke52wlZdc2nbccgdE/nJL3ef65gxVaTQWqs+kSFfqOIfsSbldY3+b4cvFXy0Jqe4aj5AO
vE7laA+BqCcf9uPjRPrQvEH01P5CWOacBNZGXjchrewXJC0fzcyUD7EAVHYsW5d16fHJG7VIO6as
V9wRlHXZ+4dWcVlm6/qTq3Fi4jT2KQNJOEhR0OnvqUFQJgIlFAWzLIWgF658N7bRD6XiLDBhBu87
4jB6yPI9DgWC355UAmbtYvTU6nFEDNOm5dUT4YERXeqfNDNvknO0skCVW6hoYE9Agu3Fk1ILPdZj
jjR6OBE0U3IId3H72kiG+3wsS/659+hZd70pN7PV1upKCVH/ixLS4r5Ov1QoQui+C73SELuq5QUA
MFNXVt0hCR7Jgu3bxCrxL1pFT54EuAyIuAFPQubCzhExI15cfXFo2oONlGGLPgI42AHD4AL/iEOx
jAu0Fce2lMQ9cBRxSAeL9DmQl5cai0zHH4ojBBIn9RwQrkO1ZaHqe0aASdHIG/mYI2g1pUJuE77/
2cd6KwzpyCnv9yMx+1cr953YJoyf91lZ2a8IvFr8vLA8HhJSFm3A7wWO5vSocZOK3gr5KuVgERUx
arEGlEXl0oRVzlcGEkLxexI9qlcWNWU1FrG4V/bsHlvcD5Bo4wrT7f9E91b1YrIikT/1lK2pJOMg
Po8eqaEMGS7p05H2n7ElGLsEXVnGGyub/D5KZ0zv3j9z/yaeef8Ks5KXVp1TTYiQ1yL1VlzrUxKT
MvuCAPJJb9szyhB46lfKaVWLVUkMaeFteD9j6/0MZaGmKHrb2pUaGcp8OKf9CXh4nqvH6XVKMbsk
fvCNwwsHo0qVvEVMl+OeZXRzeTsU1tDn+iPmNijJqYmiHTqj8NHeosiXdST33nitHyU3BUAxUfS4
bj8E060jROxcej9a5LiiCGcVa7ijF7gsfFIC+NYGXfFsCPRRu6wQW7zyiq4tclQ3WXVHSzUEGy6+
sT/VWRvantUyu2FQI2fhA/zdTMcGHUbcx2eyfOG9eQj+lfgWLKrmV1eBfQkOVFCggcZ/N3luRsvP
tDqqhrB9eZet4ldn1Q5LGcHdkJ34QJr2/WiwhXX8C9dUEHVaBox/MM6PMViERi2s0NHVAwNgiC3B
x/WudFaCOrQOw37Ycpdg3Z0yYrYe7oeQtA7fl9Omf89oyDDvcknENd/2Hpajx8AyvoZLXMvS+jaq
NylLq0Gs2DXNXNrSdi/k6E80GrFHoDpzjZHazyFmhDL/NqMxD6U6EW1mItZM31XW+XBVHQdngocY
GBd9/V+PXoOJHGg6Tu7uSC/nuZcFm2RcLQxO9Pc1R6mZI+91Q7GFOyFbN0ngNqkdAm/baws64YBb
NmsJfyZMGepoQ27eYm0aOpB9jSdevF9QfK84HIPJWJxsIyESrkHPTMM98INfXFSHCre0RXlqNBA4
99O5h/h5eA8EzC/JPpUgJEoVkpITmbrxi4qgImTYqW995cIRruTQRx4ypWFwKJmkQlul2RULnxwF
JnNBGMuDtECLwAUheQPpCwhIxzc6i+rOHBrHTJ4vsHBlbTRlqD2fT63F/7atjQExxCLAWPb03Jyg
BEcyNg02b3YiWw+vppsx4A/XiOHar38WuVH6blns/Qrz+kMp6i91XiMKAbjh84djP4oaxLGwFpMp
o0SEW6ERRFnJbhfgbEUTwdgVQiszjx5X9dhJvcNk/5JK69pGRro9xEYNbfcIt6aQMCibYR+Luw7l
SLfv9hMciA/dpD/6JChTpZDJ19Ge8llcVS8PPfYObHrT+iL9lDySM7p7Lop/J6M86DtMVecfJ3wW
iAN3+jpTjngzOxkiiqhomSYbXUJ64I2G9GxvITlt9qAFZulBxT7H7wcEM82coZpAm3pgOgc0h0Zg
uktqsGGZvc6kPT8II2qDID7MO6uraTFRr8m0RwH0+6gNDogYT0QtLvghrJLWyGsFMCJvoILGFQrw
3Nd5OHjxNXRJurnnOwBBm2SfuikW5+Kn34sg2EypxHiG8N5YS2iB0kwZES7H21tq8g/GUVwNfr9L
yAT2rGVMuAQvmrcaDvLmaVmzKL3OGn0Ysgy8au6ZUM3kZjmk1HeEODi3fRkxYCXmNRDlfsM/ccoX
WjYuHPYTCLl//GDCr/m22rnso01NPGu+tEGhsU5cg31+gc27cncwFyibdkOhLwK7DgHl682me9P7
3jg/Pb2KA+tAbSVqdRlwascn1s35MQ4HIy5xUuibDTdzJRKwT8YecswnM7TX6W6a2L8lk8HaqG38
QR3EcORBT7BN3j1eSspdO+mxRBpDcKQqS4RuQBvROSwxZsKB7ffsUa9kPFgWdyR7sm1VFdgz0pBz
4HPjsqR/wlu8o4NCvv40a7cm7JEMlmfzV93DKusIa+mppFZz5+luaDnnXqaUykkS9nQZldOZGsZ8
GnCPRMXuRQP48wRuimxWb34XrqCdSv/npraUKfC8dHW2OLxpeLvumpL4H/8a30nksVYz3BfTihzy
9ezUVEZ1UedpkggrSh3OzQ/bvdlMkFHVIT6PpVSX7ZklslQzbjsoZ3jdTwMx0qFPgk6PdhQx7WzF
rD3fFfyXztPZ8dKHGfEPiOFFr2O01gAe07y291zj5yjbm87E7fkIyr0s9Xta4vkxMLu46svGLKtP
tislDy6ChBjlSinZiqT5/sp919CEuPfsD2JghuEqFkAt4bHIGNP7VYrsYuFt4z1mje4SkSmwgnr9
56lP1QpiLibvmmciu9sgiXe4dIBisoz7fcZlRhNKOrzTVwu/y0CicT86piXR1TtARjyZuxY6k3JJ
1OZnv5b/bo04wbaq1gpnRRJCqB8aMSfrKQRYe/DO3tbfbViZ0319+xzW7AaTiObzmR4MNmOTjhUV
ujKHKNQeNkccsKfiHqUosJYffXDRneL9nwiiXKsJQXAzHxZKZQEgNucLmlo3osgpHORPsNTzobDg
T8EhelRMb9vvGraPL8TWkswuaYqA0eAzV7aHYBgjT/mw/ZjRCq2fCAddCo73wMPuCqvcIP12KL6J
23jT738puYfUoUacRyDM+HtFsRSO+T6AKku/Kjh3JPwwsJw7SqRF/pDAtOD6Qx/7bvP+9PBsQshx
OCvLW72SVrCigqR6cYMY5c3SgIm4L+eX5MlbjhvbRIHnRcDwPDPPdJ34IlVJszTVhxrg+DAbrQaK
JHGlNypeWGPjMSigWAI8WIM0XH9XfJVEOANnr0TJSsYUNJTLcVJ3JrnxztoKVtHRIdGrLQJ7Tg6r
o7O7w4q0RB1K0/mrv4WdkB97gBrkfldjUQKEjhfq61eyAPjIm01NWyAnwnB6jdoNzhiqEp/1ePQh
RwmHi3iKI0GbASe1KM+KWKKWaLKISJkQ4soHbCLli0bpQvtLD6w9q5rETMVxV7z0s+eh7QNQFAPY
PdpXaVLfyYf3DZEk/xHtfVT7C2HRiBvGl9/3YUCD5FqmF7sO+wwPD5Z/nnG/hQnao6NzKWW3oiJz
Hh9BWk3pW/1gQJoKiCWIsHg8nTtKL53a1RZtx7n6fKMg8uq2h1dUI1hMH+gdWLX1WFubF2Oqzx6l
7/g9ZuABIIDS9aSklLbT1pntqB6IIgmZbmpx4z938+gvPFDfH7u2MgcqR+x3Qvp4KskhnHnujINz
jjB0qRhqkrqKnIe9lEMlfBEB8BK3R8yOk8xNLAa0MhFGvRq3vPGg9W1eT6kGBmShAYCmMhBpnYUE
7W6PEsGSGA2IMtkmV47VGnWirHXVb8jSdJGsv29HAgmS9NxdZl+2m6YCb98s6/vjISAoCachaXAR
3rKgyshLVFO7NfYOLYbJaON4KuZg/LS/8zRuSShFtmE4W/UaE6ZkhK3fKkY5kvlcosCB27J55fI4
CVhFyARS6ZBq7SbsCRbAjkpfoPUSdU+yGrNlsZ0fl15vNtlfYeLlkrwdBo+BOQXelEPJ5Me2HOvB
H2RPw3UACI28/Y3ZK/e85P5xJzF9rV9uGR9t1Z/zAjogb3/1y+BJGUEr5oNbUysAj2PxpXCdFI6w
mUgC6uBoS7YyxJvO/GO84HhFImZc9oteC3/iXrCssNBpIiBQW8OTwL0y70nE6qHisbsW2LuVbEpx
KlX6Vcs/C3kM+xWCa+k/6bk/kr8EgxOWi9E9MOQVPAMZgtK3Ig1Gl7slwaMAftFddjMMAeQ5bbiI
JjHSjIKy92NLhIlczIk+b1cSJSGcWreuoIW2gGuK8lDk+8tPoyoCm9UO8rhlSUhTe4ofI+C5Q3Pi
Ts38vPDubAVkvMIHEB2RqNciPR3zDyY3cUsuODlG1i27IN7DYIBnlNDWaJvFwMcDmflpxt2VWkAT
nxZHYNjZM9DOKgsUJwWY+S1BN+cCMYhEIZMVdywHYKyxKkUFMzZIpQ+su+ON6Z9btA98YS8REzvc
9rTvQr0MIBPKOkvLeRyqjb8xLBzIz+0oJIqXHBGfx3oC9sPketV70RMaa+OCtacupHaFVZr2BBGo
ByJt5QgIA+kX/k3Ab8GiI362zAN+OqCMomWU8Fa3yoZHbb4TsIBrls/QJUbF+fRMK250qn6V40Hz
OE/MMcceIIBag/tnGwYfE3JIJR327rjFNmUguWMEyRzRkMBYUIht41wpIbUmmpupmLCmfGFxPiWi
LWxMlsEFyqzNYLRhR1u5MprkKpja52mctTazVTXlE3G0VklJ4UJ+wpnbkCkPC7lOW6qIDZNYsPn+
FC7qnCeV+Odqazyt/0rz9LTWDTSdnVd8KvoYHWRutCc3u1II3zTpwqkQJ6ha/lc64X43hprUbI0/
pMMZuoEM4qYu6zbk+eAbwnuT1Huve8uLNe7bbiXAMpm4xU7yOZU2xjO031QIz6i5F6SGJD87kmS9
2X4tazWtLhtaOrUfYxZ/Ee77kXJ70BC9Zs+GfamQhCh85fuNoddhUZ71l8uD13Z2vSiTvL7s/WfF
zIDLl7kZHzlS6uPioJHd5U0md1vnrnvHMCQBsCGrkaI45jq6Ov57nYCvt02BFdulDUud+l3CB+D8
cfItMqx0twDRgg2KxeEOsFxlYyvpUYxTtffVYyuPI4LC2qJ1lQhW5VybsYZ15MfRC3SJAgrjPXNm
IAP5RKMDrtawysZpoYmiZUeeA+SYtmy8dhkey4NjYj9Q9hyQJTFJuwA9cabFO/paRCpvOZgrB35J
ybfue1DcEGTOoGeDtaQqIMRjMwO31TLiAwB643VJoryPQ8W2Eb45pyD3Mh+lpFp82maEZKFijLER
cyIBBndGFLSmXizHl2QpYJoeo/dQ2/0J0hQf0PBQLMzjK5IexDWixnje53igEM0Xtst/6asY0BVT
dwd1UEOyOmYlx/HnJhNviUju3Tfk7lhL6TKmul2g3Servsb/JKOm/vtDmQrNwPcd1DWqP1B2TTIh
8fSsvqww/le86p4xbtQz19IofhcvLHttN/eAcjMWoZ3uINICAaDmb/cN6xIU3oYF0ImQXRCCmW1F
GCfRHO4MZLgOUg0KiOsu9sRd0jSYYVbEIBg/UN1C/56UetD6MHl0hs/IM29Hf9d8MMV+v4iw6gDG
a8bGzttLMuHLo46D3whhQKGmUkyyzZvY2KJQfKLgewmuSELO3l4Shp2f6xa8Vn19CG8vqe32kih+
ufyKzc2f5k/h2+Yhj1NsLbChNTTfIJXZ4CTK5L9Jp7iUlf5eOMIIBnYHLpBuAjhcq4tmGRjeIPwe
XDHEwR+JcGVXBpEWAg/KKBycLkvA50CToKNoeNuUsE6UrBKsX0dakr//J42I8rU6a/YwFWGPHTqE
E5+uKKEZqAUNdq/xP5QVMyL4DgRv7WTD3lsKXIWFMIx8Cz0aH4EzGGb/hZkAgqDekChllkqAt4b0
Q260LUbWVg2j8t4pjWuJMqiO/2RLQYMmqvttjEQFNHcNqgH6h21s+B9HElfdY7hgv226BKIL+ncI
NXDKfMl333rt9wi/Rmg6aBDegS/gPqru9slZnl61EGVLD8QMuRlJ260VOgshURRe55d0Cbn0JAY1
aR23K83bIzj1AAi5BqYGdutzRlLwvuPtTaMtRHBhKbNLPA23PH1+a6leUg33nVq6I0MKPpMCyxur
dfkEMEv8qIrSAdyOKP5P5BchjB6dSa/Q1p1sw9S8kRvvKmTFPTYkh+dTccIaNvQ+Wx68Nagdptpp
ZHrlVFDZ781KTotkP1oF8657aP2OokNZ08SM9yjsCZSkCoLfBbdfWm4BvyUSAw0uc2bsn4+PRASx
gEoGESMuguNfP/nyPQUmFJcwiSSlrVHbjS8/Eeh4nQfIs7NRGAHKVg+eyd1Vz8LfCiV4iSWPKGI3
nBRU+AhNZi6ZmKuI19MDe6GYGYphUzYafH+UnpbCWiB5WBUyenSAyK3xkgiw7OrPJa85cMo58/t+
F0tN+SUNqPPaQWk0ds0txOYLMCrbBYx3MuO94MXaVB202bK6lwxMVqCYbTAN11Zb0lT9aEpQ24en
Yqyxvbt4dWUCanit9JWrYpXeNAXzQsrs5CnoPcRXbbWHq7PiEtrashAlxHC3G8Wi2B8rALFlDvBq
D9snuglo254iKQjFDFg4kH3NNHlf4bxr1gM0x5dqwysFhXiOTCB1ydF2TGZDL8v2wDZfPsDzD5RK
b1sv14EnHQfrLqJQ+wikWvBPfcTPkshj+ORfP0arvybOYdCxMbeA9DCVjfXkGLHL5H5qr+GJRgDp
WMaRI7AYUtuEowbsHkQz3ur8JXaNynVXFmsZipgoEEpxM3wFO9A3nN80S/4pBpr09+rx3P3BT1w1
sYmygMUBPWLFSbZ7Ma8UG1p4G1B/JoKxmQc4EewRy90MNJmlzqHHV1WykiKS/VJZ5ClbBCFg+z2U
BhYZ7CGmAmhofmztkrZFstcOawRQuz3fAMzdQRjXqyqChSMwJtkz7Ohz2nYFoEkYhgjsFU5DrBFY
PQcJQo8a63k6DjaPh0oYA+OqCIPkCZbHhZcgtLVrUsyYJvRfxFJJG4BMv5xpZYmK8RUIIXpOvJKZ
zmCZcDBzXwrYXWGYxiSFVY+H8kXKKyisF6mgBeqpPFi0sRJUdxQDXynBC9jZ42FC0k5mrNDCurZe
rnJeNNZ/iuqEK210yCGaK19P6eezAwsNQaSby9b2HrZ5RCibkewGcawLvwUmVVcEaqJFTNLn/Ziq
5cIhqH+terXCFpjWjsjBgxSpHf/WjXtuOLl5/PVriJ5YvYArcJRC5OqofNCXOgNXiuhDfC7NvC4N
x4433LAG3vJ+IL6Gqq9Hv5PRlqJbe34SQpwKZ2RxjsL2s+eAtHA5GCKajC+vzhi9VZGj9GwTzAgG
Bb6pMbgxfZnOuHaHdj5vQC89iheU0tlQD0FM6tU7BrO1kSvIUJ3GYnZzoONE/HU+nbT97Kw8o4P/
9vS1JxGtV7OZtTYPYJ9IvR7l7L5WnT7ouG2kuT2C2mU5OK8NiaMJ88P6A9Iu5Bc5z5NlNlh3uRSX
Z9somS+8xFmv6ulalGGSPJ15FyWFVtTDKLP1oqYSaKagFvx7aQFM3vnjQlCqVnBdyNxLOD2fEhGR
SSfUkyvYj0i9BPsGlzpDR2iLGPhtNiCRxt9bcEOM0Cb/tDLYCuo5fWNl/6zR1v9P6qlxlA1MKiiQ
JGk8GmuaCj/IWf8wOhpMWoCbVID9dqiN2B3d465qvMclzsHXBpfSox4xSWAHkOiiWc31q4xYX+XS
Vlq6m6gEuPvIZXiWty6v3e4x1DgQZ2U9XoPAMvsYRzPcozzr5XfrrkcTd8oTZAco6vPBY/BAh3y9
kdq/oTYnscKUHiVlwQppQ5OMPbe1Xf+CWsIod6hyhWgZjQTjvJ1cfr31zS7gs8vgWiezg6pOPK0k
mcSHsEK9HqLOkSTBjrrvCxLIaf3Niz1LSFilIxF7utJdoLSe1zpqLYoHbJeuSjWSqsTctRHMhBVK
czXtgaywUCySZLO/9nfXp9qfT8akg7lpBEAnovcaFAd8mlOwsFQpnVOh6pGUADWbWUMd8+IJiK9F
4ziOZ0IFl9ajdNPXuh3iYCfmYDvqgYC2gk4nsd/5R2amcGBiC7fSp68gmK7NkLR+tR/dj2p8jSy5
sc3+GSeY+K9dBlG0kEUkkl5I0cl+YmDALNq/9pT5srkyA2s58D01jadnhY4td3U9wz+YkdXwuW12
5YMNjvT8PCwHp+LQplf51+W9X2GyIE7VdwDx3PdY4p40IujXDIzGs3jBHZ9CjRUpFpx6BP0Ug434
IH5mzID3vMc1h++BSCPTzRWjk0HRbgkcOINX6myXHBr4om3xNkzozreHGKZYMLsN4RcXlaPXy3zm
1ZE6lg0wUYSwUqpFNOqrF0Ez04kzaL6M2BoE2twJPrU83Rw22l9/ZT4sDVyVsINW7QCwkH/Z2T/1
sVuwgOyrraZ3w73MSQSpK+sPkZqQPQC4YFFxqi/olCH4cD818HozpvtiUAqpehE9MeRhXCywXHQr
3bNSkFI3mPfl/V/hN9ohb5oaS786iSkOKpUa6E89uyJjbx0zJY18vhR7s0TpcdDCsfUVd0K7+ZKP
CmjqT8DoLckIe8nHtdkh4YXF2KoxY3y/C2Z/fdn+87/Zt9uyah1zb+9//ZDIgdu2AggUtJObWggq
BzLGQc8U905/Xz1323DkVqcvjDW3wCl16mTKpLSoIZc06BnKQQk4/Jud8kGaaTuWcVakIQgKEOs4
+s6p0ge+buZ6GqAkcdT5bZX2z2DcNr1dnpIQPTKoQ/daxsGDygdxqUhQyvpNEyCllijvlMtMBw0P
So5kf3u4HK2BihAXOEpM7l5AgjmS1Jhhs34qG1bNzqNAzKCQWcNXyUtLUoJ9QMh0WgmaIEpj0QiU
LiSl9FYcuQ47i8/FidOcwqyB1s8Ew0ndbhc1oitd6JHfWk7w8Uu1bbYAeaxzaGVSbpvQEif1S2xN
odOQxe2QpFhYLJKe3FCWKmElko+UGP5cIi3L2yeZRM57lKyQimAAKyanoZp4udssIoqVDOXKfpXB
S8gY8kNr71yEiGzmMPjZEQqyk/ZUzrqukpSeLkCkvjYvYe8LyOT6sWD66gmehTxCh69Cuz60VzmW
AjC03sYSC+6KRh6hYZpJOnLvKIdmpQaZ3bdMHshCCQPbl3JwW4stUs3xQe1ybeftjZDSx5QmBCQS
SXuNSJM1ZCBfJZpv8K8xROi+8nDgjkx9xAPiawuJfEm4eod+AvTGHAv40MSS0rFgV0ZNpi8ummRM
afaTSFCkW+3l86Bawg0qM+XUkmELVfHWP1OCTGRn4uEMb6NRRXPV8KjZ/OEZ0DrklfMNkMvsjgbk
Y+HXk0hrWxuYqV9CVvNL6/IwEwDJI0LpZxDkzhuEio5HGpiWZWu7p5vprnQEPNlEq7x9f5bDJA3G
TYsNW7PYDHfFLvmMHxzL3GWnaUbX0qbrUSpWgMYEileiKpU6lHvFTJrQsi1FX/M5GArOrbZ0IMJp
XMOCS1bINjrSHqY1FfRJ4ZTGnlITRDFXGgndhiKMfEv95ZNXx7K9g2aFPAsV41u6leqSuOsVlT3w
+QrvgdiW6LeLWarRz/sU7Z7v+uPh3BKcPjykFt+l93PcFJGIIvbQQ1O8hTdpVNv/J2I5pVO94cVX
/TWCojHf9dEo+jxTNp/W300weU8Cjlht2azt/vPCgH6qrNjpZsuzDOOEkxwyv8IF0MW2omdpx8bO
U9Y9uuJRZ7ONoSZv/AxsOOQqipiQ8qW76IZKfmTIrt6+6PwFeqIvIbnG9LfJA9aIuCSCV6y+/glE
9ipS8tGCv7uID3L3w4iBLdIMU8dsmXzL816ZUFa7LvBJhXvTYHDa9Cy82+EjWN373a+NnF8XTnsY
QL3rgr/EuL5odpI8gvhewtssDG0/X4jjcN96Mb/EzklyoqOCDt2ef5BQNzolQAJHAK3GsbohiLFX
YT9m0O7un21WbTGwWt/g7G+P1EN4WaQe43bwtMe9qKFXxGaYKulDWMfNwd/6U+leeK/zQAueyxTW
i1TRhDzholwVSY9pGnxOZ4voINO/Oz5fkOsWhLLUwzUQGnOLWRsf/acDxikmh5RMCBy1V/P2txdv
ffAlfVQc7zjQtoan/hdrxIiLOVEv+9EYcgCQ2ZQCUza25r9sX6wT476DZ18JSvWBXF9w5gkzmpEa
NFan0V5EsgjcicGbKS1QkEObDaXCHpb4wzqFZZjjckhO1mr57U832oGtb/FCaHg7jx5uuWFUDbGK
368J7BlfvaI/c2J0dDHYjnDJWToPdASX45qcc6ccONJot6xo57vSTkeySGINCww0mQC0/3nBnG9L
Patbi+FFrXp2uLqSDLyJjeZdmsrhFdsBeX0QPP+lz5Y9R/0+ffg7rDmRCeOAXtOjZtUpGk4L7Vuw
QOKHosBjUipE82odRWUuAo9yhvwO6e8FL91X9a14WPUuwsblWbFF6SW9UBRrANUsrzh8Yjdvn7e0
wZiNISi7k11fhwoHg2EBv/PTZa2q28XhQDTOBxEO4MhFqkXk7QDsG8QLOXf228QtzCcsMjKh4Wpm
MxrDt7tZTuelyo+lnjWeg9Ovrt18ldVNj+47J9rwOggZDFBsJ5OZ7SjogXs2oIOsgjj2CGoWIqPM
Onc3FiQZYyV/y1PQ2wPVroej92aX3PGGV5i+ozofdyWCNTWcqQBUQ3w0DTi3e1cCrGU/jXv5s8bA
m78BSZDfC/vMLxbIwx5GdAGNUriDuCN2Ob0aWamjDY5IYfMplvL2rBWZ73D7D34jczQahVGVtd64
y0Dl+fG2p55SHnpZzrvzidLxvzZ6KCUDUh8Ne2wIoVJJoDMmQL18Mk8u6jFFdGcTSQXiFQNyXbEm
vnLAJ5+y7nCcpXqtUbf26xVg5SsAerehuK86vwoCRu4fkTZAdQi+rAUwqTsn2afZ+NVBXQw5mJTN
L/pYBApMGYl6U5twAeSGfldJF8xyX56RgCwnrFOACeKphBBALWoe/ogFrl1ReYwex+sk2uCCo98Y
MaDnGGugFUo4+r6ZbMvYdxk0NzIXxlvLu/Rz71K6uD9ipgFn/PdTJwQLLQoeziyLKhAcOA5Ca013
CLI5VkmW7JH7Tp8iKNkOLTqPyq4v+5ASjJHZs3PpZhF++2pZN8VXEN5TsDR1uY44/UunBe/8NIAn
5fo6+odrrpegzsZEJ9Xi6h+/F0st78eXX/+PiYjLKqhxr2p0Eb3XXCHlpbDZWSd8vkIqanAAQsKd
F4wFP2zcM0rRGlu+bz89qKEy3c86OvWcz8hBZAMdr4AAixhEXgw5A3/iten329mzyAnUAMiqU0UG
eb1O70yTZs1EQMdo9oQRUleqh8cslw+do1zoPmImrxMnLPGGuUh7X+IyZk+DD3fNSN302sSI6n8H
2nQN33W2kh6mAV1d2pme7VQY3VfSRctnVLGEdS7unw1nFwMYUbiuyRmX+hJhO7vRIHqiM2u/Z0nk
KzQeEB+OLJT/H3ete3VmiWuBVsQo8P48VWnySH3hYtcuZaY39SIpnP2cHmViCy3ksIVu8CQZz1R4
FdtbAsG0y5zY99Sg4a4+tQlCUHAQMtGfkXckUUx9f25OGJsZIWtMRQk3NqQINxxlkPfhDvdYtUkV
ySBILCG2sE3FYK3IkHMYzcLybFq8oCeV/gAaEB+IYgIBtFmHcd19MKHlJ9Hk9kOVkmaZDKwD+Nl3
YLscQJ0JMyHsXnuwzSJVyoINu/xxrhdIqHaY11rCkyiT/SNBXXi6HW93Y2YLH81RFJXwUEmFH5ex
1OeQF8NXWYUxE1btS6J5Db8R+EHvyIqhw8EqvKi19V/SvCt3F3kSyc8kT+01Y7U0claP+tTadbT5
FnUTa+5biRBGUTbiwKScBMN3TDone1sGnvhwxfMsfDhqTGl4609Zdyio1UjIc/j6lNEMghKPja0I
R36I9LUoCndiGb8tLJMLOnW7pLX9PgWIWzNtLoJQUE86WmBynhfBX1zGSER4PpuGLT6s2rDDR3nL
qJ1qFCIW8sL6fnUTdNKq0oF5MgkraNu+3yK0hNmAWLAS5prjuzAUEshd/yV2azjbuuyAoZFJllc7
/Xc4FIkVoKZq+W73Yj0pYsCEMuP65pDhXjNBQEPR7aJEUC6btMNa+eh0+9og5+M2AaryLwRa0TgC
Z+NJoNt/+iMRcTy6ky7vR7wD/FBsql1+SIqCFLBdZjWJKVHhvleINmYZLUpTv4yh9rLNtkMDpGCx
uHglJiLqcH3asapAG2p6Zogt97wUv0MIBHb4Hv+FPU2QtJ1KzbUWqi55go/oRP5HT1gPAoKKfYe0
SaYFZYKFRgbEsIW+GBmTVUV4DnuzT8mtDVq+J4alwDIrB4DoPYGnUnk87vj52Amehy4YmLqNN73N
Zw9WMrsgX+vLcW1gKHh/0zBWjt5yHDzdjDpSu5Bk5vVf6Ws9QQ8H1YzT6kVlfObxh8T/IdlUtT3x
lqwlr5wB8jn17DMotyqIRFkbo2GkjRUW+8FDC9gxJ/WnxtER7cWIwPJL02HeQNsL9uS4MbynFDuM
AsvxLJp+0gIFI2PwoQ5GRisrE7rHf5v8Xh59quuCLQHMO/4g6kZZNOw23EQnCzrKfIphfOjklvQP
KLAj1aNMMKcMjmh/9OhSy5CcbT63UBQaF24Qav6nINKO9Y/zL5CsEvNQy4GWXkA/yzQu6CGb5Wol
ZAj+KQvletIwjnGH79DRk8z7N1RdXlNLZRGCwcE+upfrYTM74oNsDXd4wzrvDEkdXNFaSjX+FXWu
SwplmF3Apl7AOwH3v0MJuVXiQEjS+oltzHbxnEMPM0+FZjnjb0EgLfrHPaxQ+BiCSGI6Ouuv3jbp
KhiYuyhW75iARDAUAhxvC9pRYHl4dHB4YNariqBSO5fKkGZyk5MEhr8jmqdP1G8Gi+8TVMkHFg6o
7ooc02RHqGp3ykkshYDtSvq/JTEwUJgNV1fG2vKA1RjL2gkqA+ncQykv6WbTMJJlrvD4IsfJ2NxO
xvOT6scww+Q8Xqt/90cSNwghRi497X0ZkaTxwTHI27HTsDN/9yiZSJFNYEcQBB6n98svFg9v/PSz
9z5wcJzOqExGqjOxnBHW9+DvBXgyvAhaMfkY1DEONCh44ihOGYHWm0vs/ibDxHECUiQILyVEfwa+
0zETV79MHFjZyv40bLhwlINzH1aH7LiM+ykYZ7twiY7BkdaZL0mzO4ajDiSDIdASNSsnL/mTD+Wi
AwyzePly8JJX7jXqiuhXpokvCMGH0nIlgfIKbNnX6fSxERAEDkZZ5H3qalO+xX/NDkTxn6+cjvGa
bB4EE4504LUIcwdY+30FMo1jDDHin6hWHA1uSUN5wPjHVxhFgtp9UVRcMcN+GM2orN/r16vnOhWc
+SqMxKwABNi/qAFylyBWdzrS8/WocigB/aBR7nYXHEJVMuaGlQYD+j1knOyStlO3gVQSdl21R9CW
LyU+2d5sXuFJxuM3RB6OuRiGv2fql4sGkQp+dkhvMzWJ0PFa1JMNjE0bLiKwm4hMRC/2v/FUxib9
xsNX5c7yrwn+WVSvb9z47lSbyJ2EiXK/N+n2s/eSGq00rIKObm+1mNrnTaX/ypU9sdGzjq2lxxUJ
kl6CpB6ACPqc6ExC+YGgJuUlwcJC86WDRcvzY3/Qyi9lZ17XWoP7IhTPAbeIpj28AbvlAqcvKT9w
UessX/lO1xyBfo6KRgzWP/+JzupzybTKJj0REts6jBs9xaxTHUgO1MzApk4wgBii3a7/MVbhKMGc
x0UL+W8LssUjKYJymzgd58tO6IKBAW4w7k6nETdlfZuxDJSdEqruSvA2928QvCkaEMcxn0BgAlxI
bVG0vRa3cwheBv0T474h5BBbPCmZsYNPLBLvA+1iQr7fx+qpgm9Q0rGtVBIWFvzgyA1hqWQaViV8
DRloQi0/LynugYoKkiNdNFCMhuGKnlcGttEdHyfHMZEvFOdTUwF1BSz1fB1yrE/1gPOqpf+6OmBq
3oEVXV4dvOmiY8feW17XV/4fghN3Zp4ihAdkmI/GLOg24xjYDbDyiQKrj4CIV5kVcZxdqPln88O/
CZDI+fU/JaXOUuGVfyDjjDpAYdx3/qXXcppqLrjKHlj0lfTjt0VwW9LypLHGpLQfPF1fgeJ5HvBM
/7l6C2XKbtK+VE+IrZaCGrwux8OxSuK1CRfEkaSMQMHiCCDvgdU99isRIcbQhm+lICAI1Hbn3eyo
QCKv4tiV4ng97kZf/7z9+OCOcrTwUWnkcb/uhoSn4ccTHR3A634+gPgoKe3S3c4yZAGl0QqJ05Ph
iUPhblB9pH/4XsVkixF1fRj6GEv1pqIYDxk2pV24DF4FWhwXgL+MSEaW8hLnMjUwFTUIVBbwsc6i
Fmq04fupgsgSFQXmpqUTBMHh/Kx2XV+MqovULl7yJqVW+PBvr3eYoa1okwFY2a//ptswusAZgah9
nExnTuQ6U77e1K+TLofae+s+FZPTPygqTnwpF4iSfEAQJFVZ4PPwJf9/2mE58s5eEQ0ahR3Ov4CM
yWu57PG3WAztsKycBxhU8Tei6YVpQNpxhkemmnO16gDrLky0dkHDwm4k9qVK++krVKxw/9b5mtV3
8H1Fa5yNmTy8amMl2KmDtFbSnveiHkCyBbeYKLrkBS+r+5SjzpwoklRKkuB5So9MTu5J1FNsmAvi
UXtdx1xfQ+fzeN8kA6WLrsEcSBuhB0DbqsLTM0rDqIIOii4x+fgm4StxcreNTsXMwQlLEV2/bT6P
uRe9Hq0UeohLbSMPJ+cC+ciPnsqzgZa6nx52ipYP6bGTn2DhyVI8RdbVcfFtObrMDX+LMhO1IBq0
24qYjA+WyrVqfp6UNdoatwU/8FzvS5zBq5S8x6MTro10IDeP49c5uXRbdgCFvPUd7m96MQVx6jhn
w3oJBJsjR83fVoTlSSfJEjtRWWufaJQgXNsI1G38yqmTSJkNAVgfCaZj6rOUA6Zr7oeSqtrXyi2A
9BtLQOTYgpfooswiy3zCmK5eGi6/tXqg92LLLs8hB5R7svPGvz7qbG7s5d3wUxZH+F2y2cQ7dgT9
cmEEiyXqmBfPSxvoY/u6zSbRPiU10Tm0/K1cxRVpihwgyvVq4XYGspCZHqY8tGpuH7PLS5vKinPE
9fIU/5/TkXvyqzG5qyZdg5BVwKm2XZXySvz3Hu21iTcywMF2h4dtLnhVkNv0AMk6FOuAtI2v5BYX
e2csT9R77wd63nTeRorr3O0RnNPxKaQyYtfRW1RX0y9m5ei0gtZyo4BPCbioUPAlRfxc5Z1F3itW
IKEMCd0j/sAYYgEXvGuUHhezwtKy3aSEXpDGji7OvW4Su8OP43Uk2PW9BGuWIOTu7h16iJgs1bif
bJQascGiSZBUxCGI7aD34p2U9tExrSnb6aNTNyKA/evaIeVJX4EDf5oDqdZx+YkhgJmwBGbzickO
mIAztMEpvFmnFGt9AzIqBk0IhY5ZkJ9we2zuWj+EoWah+VrqbHmAbF/7YcEJJWakE359lgn/D2J3
xpfY+SgrMppvwpVpUIQrkeBSjYr2dKlq5h9SDSfzYmKwgKUH980M7flNHfx/otB//FDFqYfbg1+9
0R5QDkkGL30XOW/nxoOUil2x8pjZWlKFN6iYYy6ZpU4hIhBqisBHjohaA5iLWOqEFnzqUE2ZsFrY
DVTCtuKz+o5JbnQhpPDLa4pWAe2oPIjcURidhvIcRunlioWJEz7cS94SWrSDHwBPa3osP4y9CHr2
vsLxmYprS+V1WzYen7xRvFEU2cAEanQ49WEv6NRU9J2IM4M0wZW14Ao/dVyBpSBmRlOtFgnen9ns
UpwZpVFvHKQ6Y95YxYuziA/XmC5cJiTl3oBA78nlrstAOzj4o8EaDqGgEeFOddB2Hdrl0AFXCG/d
hp8wuqLE3ZuCWADmB/WhTkWmAvxEUMneOXDyEv7Fj4wxc1Q3JQVBweMQN4VlHpcI4s69TEBm66J+
WqWLiIc2fNv0GgdcGoIEtZwYih+OO8sRrCIklLM8RoN5ao+4oF10K6ry9+KNmtsQUHjp62Ssq886
pRT8c2zKaMZFc4JBZdt13Q5hNjiX1UXHE2TEQr2oqRKWyMOrYfJ7nFXTcAAhFdHQD2bJgnh4a6/F
gt/oz12iPNjPgNjBYiX6Kav3OCB0FLfCI+A6tgYu/YPrWaZbs9KejdYHB8vdXhZqr2oFrHeCl6Je
EiIv2Clmh41pvbITBOPtv5G05DG+K/eV9g5832Tni9p2j4dFOTgb7utdABSAfW43jLd8qqUBE76g
Uj54Bz4mHruxSZKrCJMO93+2QzFfXcKP3BBfRfpvtKUGGV++jE1ehBPwkP6/nEHAG9TfyPyOpJ4U
zOLLBRYsmwlH0ZLFJBFsLOwbqlrENCjCYmFKurZ6BZgXSyEmasp+4QcU3s73FMpJ2ZXlQbd1pXJu
ASO4Pve/pshxgEZH0hsnChhMJRzI5nWZ+X/RHi3rtSTIzp92kzLVI/3dWcr0iBYt4cCTg/tRsh54
PmqbB4kyhHIUGJvkwZ7lNSjqZknQC3z3X5a4ha+fRHeij7dFdXCKPWs5Q20fR5z6qFzNCMWfHLuU
2Ne1BrLCt2Efc44k87hOrwEmigeM0eLPc4EPvo1p+i3EslIqMDm4mVOzDAy10jwCJBfL9gKf9RCE
ST/wxNFqMhqk3bKsXfJk/MC7+9D+TNMCxFc+t/lZ7sSQ/EtIfhiHuJrahFBUM27D5qynYnf6owd/
nv5igDWPC4N+9pt6G99KAv/8gmDO4gq0IBZPrgiEtOvt+IoHhKyag2X112+1UMZiIqU6VMZgM9MR
tIf7xPaQhEF1xAUQiMDr0lrLs+sBGhGR/wlCiWz1EG9Abjni2G1ca5hCUHU9ajq/L88hjRZNVjd5
1/92bSQdV9A0O7n+k9ikJ6h/7DG4URIl7HHSc/OpkTGeGVy6KuBgoo0XwFKxfWSkIJi6AwxyuhV8
TSQb8EMIWaRUA+tuNZDoMIA1X9DZbIwhd+BGVGih4fRoYo1rI360cwG30AyvyzYJO8selTA/BjZE
ipe2FZF0AZeQNeA7oiodjjskUWhzDMlLkgPyOvn0slad5RFQZovsgKWrs5RgpKoLkIWRPGMuFP54
nF+6I5CdcHXcU4WjQTBTITsOcp2i7LSswzUA4vM9s1je29ExPNnYwuQdEtu5XsYC8FcL+nXyrJVS
QkE3wj3vAM293dE8O9BmVABH2GZduH2ML0y1hnqJkr1kwIiZbPB3Nlqv5DquHREmO/eMi02T+x7s
PoklNBykwnKgAwixDon7OgO6a/3i6TCh3OB0IIzynaC/ODSWIzz9lzLIpxf91oaFkyvzLa0OohQe
+aUQmDHWyAH0FubvoPiBDeZc+44C6b4q0t3qkSBFUGtJsWVne3felSpqzh1HkPkPHMWA5ZMsiZVC
G+pewFdNJXbrdOJtLZoTd48Qll6ydf/2zSceficGgA+ZlgoapqmZZGh7fLZz+zUpRpARufJmogat
vR8+QoMENewpoNYN+QNO9oljvPOM63NvOOYQdcJy+iVkePrtwMHpUZdpNv+oOK03h9ncevh54Efk
N9wF+Y66JGN1Eud/a7WP98B14LxalcVP1h1ZqYR4gwTqvWOwLLEX0NaDzTFTKl92qP1IwO4pdj6i
ZcdDEKGQFQ3YkmHYco4WJb4Ax4sSw+kHwSu2VuPFe99tvZTXWaSg9UeTGtmCWmsAIo4HtqThmr5C
WgTuRk+mDJcQNXB+eFKyIOiAyIyXNXmQqvsSOlkCjFShxieehELEUS/p8GhltMha5El9Onaa9Mrb
VThbzUjHu2zHmB/jUwTgpiIIp2ImvjojfhqvoApqZrsRBGg8RUwITdU0QoPcj7slQ/HSAkZunqze
Kw3H3TeBcRok9JaOsqi80Nx3+hJjxMhU6Q1D4N2mDg2Phcdv1wNZDhItaPeWTjN4ZFXmyjhwXdpM
H44Voz9CtVC7RA6AZqEgfEfokQSCP+MJEZMxTq420JVoXchRNfkJ/7jtVz8the16etIRtrR3Y0Ie
Ngne01CzdMG3PNZwg5rGX5KbpaKA64PoCc4ogmJDvUqhYUIkLAUYWVA/yhsu2YGEe0L5WTEdTvqO
lYTH6vpm3XNHVb9cR0872j9r2MgWPbobhnJYPdc+H/9XXtzCpwcQF9Np1hwOiHSh/1+f4He4aW/+
B4SQmO13iSWRdPRMEtj4Pdk15JI8M8EXYiSG8P0HSUMlbB6V8t4HtrsZtwyR8JdhnxQ9kKVQ7G5h
5+P4XzGtRXSVNLeIkWtIsq96Qp34XOwhRTCEhvJGVm4VajxWxNUmx0hYgLZFAlms8mMAYibc5o8D
0KBm/YisBCjwjvfj8s4QsbSFgA9KLyee98VEkiYEFdWpDr0hBj+8Mih1LtRVcIDRt8y8jz8iSGdf
tExtz1BTpYIoAoAzqLhFNB+MhoIrlfi9o6lpjvW48olv9ATYh52DXJwDnnupW2ZNG9QoYKRXDrns
P784J3qHHyZE3CWvA25z31Vb4HI74OJZBazUo633AYKzGXuIpf/txIxNqGO3xXeSbZoFN0FJbvlG
Hk8sk4YQA/ZGjF6LF7btCs+NK59eWi/N+CzX1o7bQTEB+d0xZVnGnfplyLNkKmh1y0Q4K2T+j/mB
6/s2eY3kkHnsREpE2IgToln4VxVzeUs2CN6GxNnww9Epa0Au4TG1YkomEP1ERLK2R3r8sh7scMs8
3izl+l93erfM9tDj0VfqdQecrL20KnD0IHDPYRj8317exMwIpFuhj0D9DaMAfagc/Fpn3WE9t0PY
i/EMhTZkDkUPlRB+TKqMsFXZ1IsRZ3DFnNwru2vaUMCxNmYoA0ZeTjjIWVDIl6rt8uv1UjF6nTGI
nusjgVLm0wMEsymRAAzcIRGgRAhiHcrbOMSwVIKoIbQm6d9ZVy8vExJfoUSnFuNVUVSHR6Xc0ZyA
XQEXAf9kNnTqfo8wI0TagVh/AnO7z/o9ftGIkfbph20zAuQ8yGlT9H+B+wcR3nkMFzJpmK5C4XH9
YnCtQPAeBuS15P339EJRyaHMD8X4zzNSSM0aCSnygvjSBQDc0hHbreQRZE9ub7GP2OXhLIbVKY/T
xXp/rOpCI6P5+NWHs7v/jo3p4dvFe5KOwxPO23Nkqvqnbc9LlBO0Zl3rORiVcZ6a3Ay6AgWJQCkG
DwENIYif4+ZJt9yxIX6vftFbC7+dcaVqGwkKiujCdC4SWZ8l4Mzai51oXlwKZVazi2iEJkKKQb7x
2bAIqrLoqtBivMyOQwS3R6p+uY7EuxSPNhR/mxi/nJzOaj1KWVb4EwgUTuB7raZ2mgkcxJwBur1M
ZrTgnFCFNeQdreZwSzZ1aXPzraSGYQbCvQ9enPoyh5JYIlPv0O9ohCy//nNvJ/K9VXXZiVQssdL8
QRzNWNyLMWN8USfvmis08VTjbODvaxu0lbkPdkdXsVUuDYfelFFRPzRDJad98AB5VwiR8zwVdA/y
8HSb7VIuSoTTDB7O7aJwHKl4n4wVvTZanL8i9qqfUW9f0+F1y6eexyU98TFI71W/C/Bv1xCejA1G
TqycnWIe9aiPqH/h+gzqfTqP5wenTNGna25CY77W25Pj4ozSrH4zUwjSvIhOqbqNQ6AFtkuonBjL
TAiMY3C2xDnpai8e1alf18dRf8+Z1/6gwHRzmw/cpFfr6Xp26KfHGwCC1Fnw7z1vbWAra0ubO4tk
+7O6cn+1g/tWUcMLjcwfvLEr5stcv6wKeLC4dfnrgiPxvILC1P3cr2cZ1ddall8i+tqve0Iesv4e
y0Iv0hgmhVON7r2CYPdhChjI8YrcpO4GKideUgs30MUzOJIr5vz7mMluL0QKcYoKRyQf5CeVMaid
GPhFjO2oUahOe81Iim6gL0F2ijy2KDhwBsggCV6FXgYmzKcKDNVIA+LtfSi/eS/YeR3no0IsizFy
Fdzh7pXC6UY92JnKdu3WKaRUhl2sKTCGWcLmEMMTiZI2d0Ioqt4Gw5fd/p5FnUleX+SSQ9MdMHE8
f/bRQOGTaYwknpQH5wXaO01c/InDnAIx3S9STrgra7kwojmZPgxrwYEnhoALijz25hVW5oRrAlXj
nYrVPgvIqr4e5Gj4R6zjDkU2QCetMddqG31XivI2a/rsPi5lAG7SY8Q8GiqhSNQhsU71CUSKOK+s
13vHofcEe2dbVH61DzaFNQVR6fcbJ+IpKIfXsAQcmIF0Bm79dkg3k3eVSLSKh1MB2inIXL/6sk2C
FnE592LPRQQxnKzCB3hqAt9XK5Z5szju4rSQlhyvgCbJ1cf+J9jspwm9vM7xtKYg5FtreGZtk0eO
QEUivUVC0hmCWPbvbYx719P1EFd6hsewkJxQhjVdrGDEYd8L7lgpvoSzygmgX5WiRJEiBokf6KYi
2b5Wij8RcgqhMFu2ugnyiAbHNt6pZrOvaRPeBbXLAQrwhKqKjLMktBdFIeBcCgo4iPNZf3RSF/q7
JdsD4ecwNaP1T1V2GdUv43t3X8mUNML26cShVHZaPZjXFeJ+5Zo0DhItCqeRKOJqgqBeHPRRNIqU
BQGoFfYMG53HoSL22Dyon8hvbXMckeKgXPcnfPyeHqa6IXU8lBsIrwUFXwdkbazefU6XtCcKTawl
972lJ1fLYqWfMnr0p0NdD3DjohZOU2lcH3hVBLi9kgM2GF0YcCIMYEgYx3EGUa9wJhJ92LYhykV0
jcbgDuvRhV35ymEq315IE0yszHZBoSQSiKPYTlKVH5+mjV3qrEL5oafnW/k3HcaeJHTzB4TPnoH8
UG9XMl119ED5fXKuWMZC5tfzleo4H66TB3UUEGvMXJwPMa5IMD+/JnLovK/kZI+Gpsz1ftI/kY0J
k4SDjYPhHJKnWruJ9Fbq7ZG7Jj9NyIVnXCZ1P3m0D8xkECmQWNFkzbNCHN1+gGDSYPFifUD1tZAF
XE6dL+k+VaHZO+JhWwFKB6p+az6tK3QeC/kNoPYlB8SLZprlZXfbg3gt3XvrjxmryYuwqHHy7GR6
NVbU98AXRflQH9Zc3zNEGDfFpXfUaF+5IK7Y867SMxmqVGGpBj18v/r0jmswh4lGXQEd+GE6wAld
W+qnsKif3AH2J1Vk8ZP6VvxXIxzose/i+NG67ZQOu66aZR6etncXjta8aEjxv6uGl3JQ8Wy83RMK
Q0qdqd3pKdzm9YGegMm3GrCnyF1+E61cT6/5+/oUnaqxnPvC/JcDxhrB/Rz6CLUa6HN85U6CAwcb
kH0wgnXSToJDT5tUW2Fb9ODQQ//EH4Q58+usc6Jjaw52bufs//cMZKJucCZNS0jTt6o7zjjMfSQM
GcV0pz8voXeSKnRvQbpW3Vf+X4c99BRlg8hzTwC9JJw/CAILeX0pqRwk3yskdIAExQ4hIUdK30OK
phh0HH/+21LJ6Y6EMLMY4xAFCtFGfK3AIVNV6Rcedpav7qgaH6UF3zuZMGke7Xn1CezOwqdYsFVp
AyYVxshlO9VcDIeezUhegG/COyg3A3k0ygfzyLkkrCAgpSA8AU6QDpXBwzhMlq9iy99uIlhygBXw
dxh7VyI7c2JUzgfmtPWG0U3krtBz+YNI8hIr/zNTZmYKCuH5hTos92Oc+WVgy/Zar9yS6duc1UHv
m3pOVB1oZkv+NgDyAAVu5kxDf2LN7ZVGjcUMuxpn6IOwWJqqwnjetB5lBGHJP57dyHXgE83k5EFQ
VEseGU6ai4euV/FiF+FGidS0x3ReeJfYFIStywfEscPCwjDlP30oRixcecEfuffC+KvXCz+MXySS
tx0A9nouMBiVYskMcugtYyvpxrHp4EYMlztiDx3rNh9NnnbKBXiBkfX+CDmRgZxkQcci9b0SK+eO
0X8Zo9H8mxSZZvo//Kzh8OdXOWT3Dz899mC8rFob+HtPZBphdWnPyCBeJ1PuGu7BFqGPNe+/F1HV
T7wUHrY0XU9b6XDBZ1Awrrd9IW+ouGD4J0X978VDgpSdXG9SlQJV2mTK+uQs1EU6qZMeQh8RXBMg
5+gRi0cBNmCiLcNOycAuwz9bzu5jOEvkvWd3HqEt3clmcHKLuLNynN8uc4lRCPc/pV+4kC/be36c
Q1X4r1we5CeFjLhNxN4bX/cfo8GSAt3qv93AgwXBT06jSf3miCQtgAxik5qJqKA81RKtXx5Xz4MF
M6fFOa8zIffMUF/xiriekGfDQVQ/gP19LrU1WAujjPz8FHwpmk/GiZklrTmkIX2deslYWxM7hLJL
jfMcq01FnqHlsZNdTn8I5JKybAraDSEHMFN95vUbS8gvQMmwcVVyKlWfMaJ9gZLl+BfhrYyu4xG+
08MqQSxeKeRTlH6EKxmaP8QgSPRAHWrLy1kS7W+hBOG31aKOPVXr730ew11CvlQhrkanXRfGE2qN
SsQOOg2f40jZwUXiXXFN0DlvINp7byexL+NIdpevsmIGgQdKrJ82W7lg+RH+Ckq8TypmLfTbZF5y
ZknoF6tKDa+VcRGjpJOo7wi9P3knFgd5PNTUO0rLom12ZM1+DTdEq4n44XCq03MSiDDf+ezVdiK0
ADp2lw+lSf5ROhDkDfClxAasqcrT3idO6/D3HpZ6zAHXPN1V0Ko8/x6760QKbw/aAihx9Qbke/Ib
7+whItprB87RvbMuUyQ4KZHTp/k7MeyEW9EdLPHm8pEVxfIEHtMYz/5OLI2UCIteluWj89bQiafv
HhaDzHC3fkFeuVsMcDQvhYu1T8BlyKDGu7HYIXk1qUdCM6t2pn/v65bLkViHWZjQ4fnqcRRB10/3
hjN9e4Slro3qV5GZp7bClMhNgTCChQinRUuF0/JR0ePY2Z6zFBtUlFG9WaPoyUV80zUuOGBidrgR
G7sWrgybSDZ6gwWgNfNmu0Jjeu3FKSC4QiZuOklTpegy5Dp6p1A0XISFWFm+kXiBguzE3zq2YQYu
R7cCYHMJFVcGsinLz0hN0p3RMwJdYvCKNDqIrziq60m+YhOxrSmLeDF+6T4y1IsTLuLOvpva5QuH
cSc0jAo1NuHzJnGlZLwp52LeU9HXzHHDtgYqj4+xKx90BvtmaAb7K08jCDnufb18OJnySItRkxyy
tOwvhd8KUWE2Bxj6F1WzbpDo6yMVu5yLqPssFNJZvNFVXyx7MRIWzG+DIexWxHw+iuYdGKXvjNqN
1yUGEhjrEfRdn5vKrTscMu5y1qndpOFdfTAqS/iLTgcQ9zveMmH6tqtdDZkqD9Yh/nuYtG5NbtFh
NZiZbR0WKheYgMrirvotunvtNEigZwV5TIcjDaLiS4NVIm60Q87HjdNlLbHnrbWb9P5WYHWRp+Ph
cKdYdDHiaju02NPZWZ4V04d7ZF8jXcb2OwyiNuoo/yT89cxwetMaUVSxnD1BdpGILgbJrRsEwUy1
SDz1tOBF/pW6Vk/I2dqnHuQXUBMsms92BU6NsT8AJGTJwemj6qWtWt8/fWI8va2+/gBKgbERPEmM
isMhs+PNTrpczm5jN19oWaJ/FX1UFvi6VhrRtoPL93eoNp3TkMo1vzREuFzYjw2l2DQP/wQhfiSq
NnG9MOZauCgFpb2PGnxkRyr1zORD191/XXyPcZAJ3icfZJNIVlWE2DcWFtCVkfEnETHGdBcqt5Vb
im8qaQjz6f9f6PgbA69tUVVS2NGlVF2oMPFvWaPdTiU0335vdc72IhG4eryGzCbBSW7QL+ASx/DU
kVUaLnu3rvy52xTSwy1saur0AXdmObx7A73YZLYK5JL8KWcUU8F6z1Ky1g+gPHYlAuwY3BDfGIl4
cxVwBnHPvtGgqXBEASpCHznrTeiBzDsnvIxyUENadIDj/bjyC3vo8oodYVHfoKkCMfpypyB1QD0H
N7Gi0FsmHbGWBrHUUauAYAA3dGg93JaN78cDipic0nOw/ID/A+WwYVBIntmVhQ3GqnlH6rPgeUs1
WPLMmTbGtVz53u2jWc5Lyrakt8+EkmunM0jQpZ/tVsiwuH+WZedPlKX1EGgNcCvIHhUtnTDY/GI+
0ED1WdfMEvz6UmT8EevU/O7J6AZUq8askSgCR+jzjZExrVGqB9AsWftAFJEl/8tjt8rH76TWkhcd
kzcyM3fq/LIWgi7RMlsq71GaNXyCTCIO2e1pBAVCWXgpwau78bWksVivVwyX3x5zVMUIspa8flu6
xOHx/bg3Zl8FKeGa3938kpc+xEWweCINM4B0taxjcdlFdy3nb67Eh4ioWhTAt0qK/Pdq4p8yaZ4J
JGEqBoQSXDwCd22L5u0LWZzJzmy3vjoBzubCe0uVeT1LJVY1j/qJAGZm8RI2aWyLEBIvuySsPnfT
3MVLSeOssnhE96/S3c5IlK8B87rJWiBz6dso65b+qE+4abq5Ue8vNcLItd7Z04wiIbdg1GwUXnLs
9pdELSUKWT7vZU68N1TqfYqpjD+UudCAixprBa52aXoQ9Zad5/GdqpZZflShRN4eJCo45Wc0+db0
F5rJAqYHB3Ze2XjoZCjgTLwFiow+NyD2A9NpgBuaBpvc1CvvDGF2vNJedvZKMqU7UX506hE/+PdO
7tZuoJRH+h2i2Q72f111sPrMaUs2hsff97ujP9t176NZCHxAtRd663IC2wmvt6u2UPojnUDdGgy8
fzgMyzC/zZHMSWevhQyUbA8o40IAhdIGGB18tmG3+euzs/JumdmaewZfpalm3GRK1+VUgpjF0H9x
UoXOdmsNq1H8ltzU5NIASrgz2GGcIv63GRbCLlE6NGl7v7vdvUAoL3zHOkJmMWhIJQpNydsfYElH
677YliEWxKH+7MF9OMCY6qlZjDtkZRg4V/lrsqfEx2mGQ+Tz/eNIzIJ8pEHOvbD8/d7Vsy67Ifz7
9QMqhK5ICLv3mwT402tDFBvyoPSyVpcNeQpve5IiR0VhV2JpSNuAPsXXFWJwGBJxrn8laJ5NjpRL
z+MuToCn3np/m3maZhR4h2rklFR7KH/v+VqvFX5l68Y+QKHVtY8SyJ0D5kf2EfwIH4Hfgp+W5f9L
qSjdfdFkV69//0B9hVgKG0UYnC29MZel0KsAihxBQ++6XTLvYdwoHVoEzyG6z5A14Wsy/e5gEJk8
PujARWiLHSjnljkBHJj4W6iu+jXvOfg8sAoRMv1bxSi1hHOdksR356h/6u/GUZo/0uZjsaI3URt9
npEKY5qp+y4VnW5fOCUC+N6n2xhAMFd4sSvq+K38seB2WN45VG9CUwDVWC2LSirMkrr3gz2EFj1y
uAMulcvESSvNlHkh0m/Fl+XlLEqKORLUsCxKra3LC+svrDZ1B12sM0rdAf9qCsUmCwpFEPseEAmW
mUf3pNZj4kPubztD/c+JLmoLjfpzx4Jy7ye1UFeacV+i3+7jfsIyfkrqujUBAUQcSKOwrcd171We
ZK3WqaMCEOkav9Itzsx5+XxYPGExCRLVpJ4mATmhuPuIOm6opu8zb+6RE6JorwzfcRdsa+DjJYRm
B6GU0dXZU4EuvVSqLfGdSONp/PRczzlzgbv6lpQiELFm40hhpvjTeEOgY34VhLAt5NCWlFAo4jcx
TxmVt5KrxrXbvjT5cafG5CWXfisGvDMJFMAHeFjOnh+InGJZjYNchh3LRz/0TeZ030Ga68tVG2S/
0WfDowf52JKePqlrIJvIKclZQsbRbrnFvkm9s/MA6ILQrnRJKA9vv5Nv+XxJWE1/7Ei0pJ7w/27I
zQdG1nY7c9rBNe8ongeaReLTnEmeX5t9WhnbUBl0g/7oAyGxUqDWTQcDBJkuZmkScm1jkhq1LR9m
itBblagyq/V+8rK4qf7zfKqj0xGa+G4jFNwnmH0zsI5zFt1296/zNrixeO5xOqwwT5thUtFteHGT
Vkx71zSFq1+EYqAJSWqqFoyAFrNauGUZSLlzWCi5fvtKFqLDxKI44gjZu32i3RDvh57f7bXDyiia
+6Q4mIW1Qf794DhG91oixe0AAUsPl8yImJpntCsB4AulIXlG4KVxAT+EDL2XSGIfxrorFcCoVvr9
QCbm5Ry47UZh9c0oly5pjRQFwTj9XbGGZk52bIiWok4M917LZChnMPM8vWLC3nyRC77/9LqDkyJR
fNlN9F0I9K4xhuISMEVShn/u/Sq/uVVEqrc7DvdX0OQ3WP7GkckbV95SMc1M/b69OKufdmgF9Opq
fQixTCI9jwJjj+iLBuijwyzYn1FDTGQBx5Xo+4ZUmZQv83Hsd7rXIcU1qVwCSwNXhjw/ClOkW8Cg
SvAkxOdPTJYuJysTiRiT10OcYAYXDRYSyEaJiW834RFjMzgNiaCSJ6FeoHR75gYP5FmJIjgbmTwD
XHzNhmTAgPvQ8+sCAoWQSMqvNhzak07oFG7zMnO8q0HFXjo2hKH/lBhdxVlhYaJgefnMdaYVCj7Q
9w9mZUalGbExxgw4KQB7bxi8+uQEmmv5wYngO0T1X7e/2tmvLLmsqAJBWwaJEQU/2Szk1pa6ya8H
JQb4lMbPbB7sD8NWATYnPYUaLHRk7qV0JU3QUhvN8NqDE8mPdlt5JC8tqGrUGJg39FzRPPPao/Dg
70Qd9+4Xvi5IYyaaK7u+5mta8ubgtXu6EoasCwLlL+LiYhU1qaWclTNqaNlqTrR3xgQXz4YDrzPs
aZg+vkY09JwiTqmDYyUA5363lDvnF7wzxtPRyuIgOtpBk4cGmetfoAdiyuujwOfXnWRTBCHa4A5V
tvqxO4VGTZ5HSNIVMXwb3EQiAARqAjOuE1Pcmphb6lzMo/+qxBkTDQhe9hblShQPyh43C5HSnWPP
GHPkDvxw7y2ov/0UQgBBG8Yms83RvVab+oZVzGNG3ZPP9dHDqV9xw+BkZR67EJHZWk0SzWWcOaZw
q0g5X1prsCw2fpFhxX4WofmwWd516wwztQ+WIkfGGZQKHQMohJIwavSAOyOXt0dk3X9MUmGpjK2l
/BsYhaEGPcztLgdwfN+NkLgToapdP0QLHsLscyQasy1xwA2vj35+mksiAdRXnWcZX9VMpuRvnHH9
FLsgv1cHBHBu6l1M3bSQAWCn+MDRid0Nv4g2QeH0WFXVAhnPeEKdINb1xRATa4n5rKsm1jZaGtUG
0xycPidoET1WVmBkjeTfuLGL8yWbr9v71z8GYm+hsQLf98RzKGuBc0R1q59G/khdYWkHNaGw1AB+
ArH+nOT89ygDSBt1Bl+gJWWyhVWIJ4hfx4VbPv9SW9pPAO5ON8b/2K5qpdgMtoOttBJ4cGLmqWar
YGWW8RfRsXPqiKsK+YtizQmyoYSyByz7AFyNpcxVwfcIGm+MLEzSBlSEPQmnF6OQ2QsZXp8+KmCw
diymtb67EpFA5DmIlVfh7w1UgNQ1LlN5UHmrQ+Op9ds+sZHfgeyeZTcM3Q/QKJWjtPl23bUTve4C
lyo4ZGA1PcvsJ39PAvcjNK8Kbl+EH9HC3SMiiTpCw2qz5Nqk9diM4qaR9LPJL63D92BSPHEugTzE
5El2psE9SRLq1hMCcstDe9KgPCXiD3VPEFcRXkKa98K/DfTt+UFsm0QK/fmzTd++AjESaG3bzjoA
yksf6P8KXTvF0V7hSnr2I0NOdyM45uwuZ/7tP4uafFbQP8KNPSreBnq3+uaeBDwwQ9En+zQAbOxM
AsmYqsiSJMoC88vm2bIRvXam7j2czNgRDnsFJCuzDeDe5rwAzVvRmXNfOh+xuKDYlfneTqubH3pS
zxyDyXWDM67+4HBh1E4oUCStEHFphGOcyF1lRYRK/HrdH9mD2TvMhMfXORAIms41sa+hPligsdU9
WGY1IVT+rTtfc0xQqcUpZdYe+OzjQJfNkeSGc9J9o8p3c0ekNWbkNhVZnW0mFGNndOk8RtebNzWX
VZS84fFttC6X5q9MIYOVAStPEJx7GN7mvgmw5Bsb77PbtiLke/HIl7rVo0RtNBIPajWHys3Y+kmC
ymFc6q0u7IFcd/GpJYAcyiKHVwAYgoPTue4v+vX9oNbV5CdSXmELT4+d2Dbnxp13lkH6hRgW6Haq
/3BkCgdpBOGpApMgVygYf5n9pV480vMWW/laR5jf4UTOa8NJzXXC5Iw/RHEYNseQgHXFv+nx7uEJ
tN4yuy2DvGrG2l4G23hL170jTGxlYKDzCVArZxIH/qBKDO9/ulY80n3Z+3ZVM+OSTQW4hI2ipzn/
TLCroLF63UDeZMKM6Igot5KqokW3ZTRxoSPl/4qozp1rs2ffT7jQAsMPlUaj3jw2mfGyPVb8M55/
/k64yYlhj3h9OYMqu2RpFtawCT8hvLkjKiFO4vP5XCEtzBYNgDMaxUM8HDay0epgjN7mY9SWsdFW
fwEbXZ3eBephugPR9CDcnAyBHKXNuiA/kN9kGa6izy/w/YfUsVMwoB+0oCKYYH5l7HrfRqruy0ZI
MKUKJcLpzQHIaOT/7HtjhCf4+cTtfWSYIEyOGuWRJV4N7PRoQpWkcVuGs+T6QCXLILaEFnaiG1SG
ZkKSDGD8hUujUZzGzqAosIGigqeKxc4G8/Ba4VAkgs+cP3+c3liGHqQQLF/brzOnnE41AY9ZuJr+
lP2KgkWRqGrSbMGkvR6CLofCdKUGcRUeSFyiqx2WbtbdI1/gXRehm0hr2m7Ef4INLGUXDU6l6GrV
cSWeiCfk2aAhjCsaeCWKX29saRCAKSSaP89mWfMkI2ETcXthhSp2DPUyAgm8u0IfGwTp78gQaTE9
/WDzGRSkNAkLM/JOA2ubvWqq97UCXr0z0HwIc4j+86eGk4a9721bswAng/0TzPXdjibuZXHvR9Ti
gPZJXssWFw1z8Md+kmxlqvQVdaE3Mh2Dj7ZMKF/GXyYCw/z2awoGar1AhlHD1Uc+TgtD14hBgOIB
vs0T+67Nm7FQjGQUbFt2/TkV6Vnr/FGcvd62+av8wJ85RViEMH6u8xZNp/SudHJxnUxMsHi8HoDu
80eBb5I+ONy0D1BkeIIwqLGOxlJBk0HRzGDL1EfyAGoJJ4Vs31VOkJGN2sur7gsC877qouehmP6J
5NvrEfcEaLQDq5BRsL8WC+JKtZDYY5Mgey8MIbjZr/+PtvQnd87Mx9Yv+CB4S0swcAgKMSn9ZCQT
NGLMwBG7Uk1M8dYQgOPfXRCX0KXOVl3gA0A2p1Q75yaKFBWyqUUER1kCvFEbmqVVkM/UTMytIn90
fqTubfp3yrarrpDUfUcOTXIYG3oDEzOjYjQT6kVpRv8QlXJQ17+xziXVcTaObP8Hv6L+7FGU7rhQ
XkQXW6u4GtoppwLPErqgDq1CSvUZ15eeYqDCP8x4Jod9R3Bvl6FjtUhC7uS//g6/ZOZaajPbvXeL
4CuYq7Lphztu1E6Oq7uHLBIFuHjjfyo+nfyD5F3BMX7SsdKwgttvVr6DrtvnZodJu3K+cUotcoJG
eOyFRCSUel16+Yjye94q4fVz7OnTyIms6IllGjgRTEcyeFcsG+bll2CXY26oSgQY8kUvibvp3shF
moSkrZK+OLMsL8ZvSRyeNwdZLaMcDj1AxQFy+f0qi2n06cfPE6pzS54b0qvcJVC3/ygg6ysGRBzn
vp2fKDP4UkjdDjIGtl57SS77g0GtK86RkbibOdkIZr7uiJGuIEzVf0IhCI84thMaL+AlBDRZXC4R
utiLGXL22zr6/UGxy2F7Vm1QxqZUWtpOH8huICabQoNEHMEZBfcbXfBUqoMeDwnGRZYipKznsoi3
e2FDsReF2iij6zcSBOA7uVDgjXdDn/CX1950iRNgR89QHdGJOZgvAO4JqqC+6t2cWWNUWycqpmJt
ECFzQDXmaqUppF7qiOidiFIs7kREQpu2f/Pp8LfKclooDSxQZ4BNYG6f9VELSL+aLKmvv/jRwuqt
0pNVmHUfXDvxgk9G022wM+BL8PeQ85txelrsmhqctdUqItCVs5mfCNhSMwDBbvgaYidUU5OUTBWR
qaYbK7GzgdLhXxkeanmUksoE8D7VDMd/huQTTOaj/kezIW/q2aBAhyTepS994+XBzroJrp9WP2F/
kwwwdCZ0JxHmzQ414IdmMwSr0A98PjRazXciaYUt6YGDdID8Tz2lGRG+VJBU7SMfceQwe08u2z2b
/PnztvBWu0+eFQdIU7Bz/dOj2nhx1C1ZtWB2E0rrhJSW7nHOYpqdNvbf0hZ2fbqx/Aa8Bm510jyz
SKCb8gIEqKDryQKyE6fFeyQ0fH3rBJ13DbeiaxcV6AEYfhHX8H18T5TI4YXgm1unu6I+1PA10Piv
cL8UrhonashwotaxBM6/aG9WdeQq9iCFhtQTiWTVZDJ6HyEQxKhwn5nFo8Oo9NKdm9fF/p8CRMxJ
qjgQbGzACAItGY5W/D4gD58c6rGCzeP87fmTrRGSuLLeF7CDpUOVt75f7ETTA4u/dKwcMKu5fJbY
Ez8g2rAF8wEyOSrwlijSMNWeDgPDxvICOU6mcx+kTHD/JTBdDNbzghIqAUmZWnJh3tMZMgZ2Tew3
Hgk+v/Z4g634Pp/vr3q6BEaeaJ8g4V3hd/xWvUJwvKqIbvY2CuH4kowSfh/OUQdvllFlbtKKGDmV
tPK/2PMkHGeDoOgj6XJYxBzNxAv+AD2r6/rFtZSgeAO+qQoiRQymLihIbgyIXKSj0ao87LmthKFv
UKJUVAKqESUBJBHqWZqkvPvEK/4ZlmjObQV7Bmh96FiJsCBdE/peA8i3DKvRzwrgSaL8lc0skiPD
nZY+A7X5jv22ftK7ANUC0r9GcaztxTEK5/DrMMg+95OOXMpLIgbbYOFY+aqM18uOsNSmkZIpKrX/
3x9mmT+CGsstYAfLjHztOQSlNOJIwc9405ucRbtKAkpG+FwpTFSbO0CclEvGhsJzjh7CjE8zaHxT
LtML5FvQO/b+8s3PNN9y2vmUcFF2pDYDTwJ7fbWKybVVuz4+gdsj4+6hRP6smCiOznOoaXZlV2Pt
ZdEwwvIyY1W3spXNO86KR04KCJqU/Rr2aEPe/CnUBn4T5avoYKGJup4vFk5i/h+l95Wr4cjbBBe8
bJJ97kDamh37AJcEhgnguv7XfJyDU5aM7c9uvNq1FkZHq5UhuWaDp/3LbPT1xWEk1j5BBoz4xldN
yzvotzDTwV/JtK5EnkFGolEY4Voyy6JRyhiDhS0TAR4czOWo1A2U6adkvoWVs4mWN5TjcJRI9NvG
PX5vk8sBz6Ip/pmawmJ1kwTIgrnkyAx56La1LeuCpIlSt6XRPzJW9ss6G9T2kezLd8iaMh4iye6G
ALHY+0DhtzVD/z+U083/kOmYZxMSLqw++WHZl6LJD02OyFUr8pQGtvm2K6RwctMBXd1724LhTmiS
8D6vqS2dGPUEpydcrrL+z0V+zSM90jJsNyahezwoSn05t+DkWnUMpxd1jxuh4QkLGGJgA+NwWp4g
etC/la7Vhx8g2MZ3Qwrs38taBwqFJLLl2zCERZilSV4z+p9fbcYjCSuObjNAJe5Gz9vVeROAGaYx
1fFhEcsFTUIwn8uffGK97Ynit1x80NTaPbppBEaHdpMB4pjSLao2bUBoByhMePwKUSAeQldyuHgk
lJnTk9I9/63w650S8m39tSBr4qo2QJAAWoj4BgbQIJsWpUFfx3GMSW0JLfjcj+ReioUpGerKesbi
m6dK6X2esAl/4UlKz+JoNWwMzcPuqneqPf/8/jksL3eiqmaJc00RES4JzY9HoyL+hH6xIWccIBWu
pyZzWcvMIArNB8QJ29bI9u4Qei0JJdxvgkV91ULh7HOgTbAO5VZc4y9zZtrWjDL5IB3zzR01ZxhD
UK/2LftdsscNcMlrkbkcLhV13YoPLL5ZCFk0S4MhPvRtb7llaGFeYVE7a5TKKrb7xxJzM82kzQrt
Nbknba7ojNaJYyeK+Jc1/h4A+y8nC9ycXQq3coazbwacgYnVHgo2g0lJx2PX8LowOM4JjzAZWZBp
hsugQrQpRavEy3eadxkrXLIKyidLTG/qUa+aA85fGptRlODKCE/yL03h1kiBajDG7EvzhK8d2+gW
EFcfn5P3EQ3EHL/0zEOIoMeAxc1eDV0ownfR97FSt4FJtjo3ngVyMquofMhY2tDF6Mi73rbzmfe2
5OwC5fDsj8i4Cgvoru3CjlXGFVc7MdX7CQWJpKTR4zi2z2WQaiblZ9L9OBxp+ffM0aDKcnwGoWZB
8pRsospBn9NJr2ABROxUCrhTC8DCejLHUs+nRlB8pjPkzh1AVLQf9cClgYR/VZCDHE7RqJKpyIlI
eVNEl/NJqp5euNVLhDAb77DiOZxvR1y1ngQKoka/pckUBYbqE8ecflB3WcuEUB5/MhEXjy1PAAr2
Y3CGZv6hPJMQbCwQaFySZ3iQBUqCp/tCHtXJ7H1OdH318hwdqTlxecurlIpSaDLxs+u1uwQqcVwf
kGP6SeUP37wfBrPcLmTQVEXr0cfn/3wPVG98RjdlLHEo+VyNFOM86B2WysdILBmpDlya3jSBCQIQ
xNkMqLEJUqA8c47NY5E88srlv7OQOmTIncNsBQdBezut+6S/pU1rwtsrT85MWSrltWRp63eZM9oN
I9LhGpHel1xco0VOmBzCaysDdtmyleOmkwt6wT8PhpaHgMrzlQnDm4V/4DAr4IuUW4z/eozYe4cN
2vsJK/HrVjo3m/CSOv9TCzgHqjrE35xBUhExEpTnL0gctd73Svn2Vf6iT6GpdpzgD19rQhuPt+Tx
TlcnZU+PnLEhuAqSJDkrM/vzeqwLxxU/dSf+1/D0m4WgpJVtVeSJGS0VaI7exfHN0slX9FMmoY6O
TEMZNyc22TBkG8p1FJ+sDKDJiWGiQbVMXM2x2bUcXBqQszUclMnceu1v+wB/cxISess2QW8/WpqB
f+mEeCPE46FgZcdtxZNt8f7LL9ldC7PTcwZTKU6Fk0KrJyjW56ffRRnVX6z8IeJ37fgc4sbVy9RF
9jU8Z2pQod4ROKzkgtHCkBDpsKFJ2SQYlhWzHe4YrTGNaCiRopUFppXLmmBUIXM/GxpPYllSryqU
7Ch/JSIf0GsUjLNwwqjXMNyUBm2NwYY5ZEKjcpwD8EEhd2IqOtqZQghA/yC9953Ej7eNcUf+Qqjf
1a/+05k+mzRgbGAMB0NhvlgXnn7p2cLaR+hQfyk5wEIlJLyBhufaOP0Rdo4lqG7MdWmyFg8Q8qxn
/OUgqyylZMioeP7eHMZQoUMDbs0w5ls0Sj6CzjmeTTk2gLKU+0xr3vwga5EXlcsuJFHGGGhWMviS
I3x2Vl/sxclpEBNZwheixwLFOWl6BJWwu2TY1jMdGxQiOPuluThYnTDi9ldmtuQgGfdrYhpBIKj3
xNbOqmgANoIL7sfbX1TLQWDUfT3lUALh0x9QwyIdCskODFioqIB0EF4vp1T6Ymhq/SYFXExHZU9X
wNlp9uN8blYFYeRnGFs0qBvQk+sOFDzJ3qspr6du04eXZPxDbiI9SvSuuUpiP4oT1P605zygIC/i
71Z6A1ctDOVJI69DYxtHHSZIhoBGgN8TuamFqmC93YWJXfYPk9gt2yqg9MopAwgs93+DpQcMMVix
XTSrWKrjeSEHjFHgZhX/Ox+h9GKY8DmponUf63pBpCPSHv7CV6i4juuSjqcwm1eQIrpYxRRaVMQQ
vv+3MNIFn+G8pGH+RNifJfymmJzxSxyaKDATMenSS7Z4ru9Fw4kVmbBlpQiz7BT2L5BUB7KNfZ6l
Ix406MKV68FlKvBb+qGDggAJUQgosNmkWY00btQGHI2W404Cng2WrdRpJpg9XqaBJyMShS+LErWE
w/Rif8FnO/ujIkcrg1bx1ajZco+VyN8+Ea82RbrlzyFdwb1T2W5DVBg234pbUb3ZdUlj139Ad1Ov
R7W55+ChaKghXjDUbgCpbRVjouTUAu+R1DlvZg00QmMy6b0ESS9KQpLgim0x6mdrdPbeBHD6EO4X
lYCKtxgCdEhVceqBF7ptZEHFLmdGqxqaM4P6Hdve3hHaKx6QPdY+nYkWikBy7ewwIXrsMJSbqBHA
pEuN2fM2xOn8JEmhNZBBd9TaoXfmCKDRCPZDO/0fb3/LB6hid6IjunWik3XhyWzLEcXeh5csbQ0r
iRCc7V1UMfwJ7idKBNsh2CwAMeLu5fRwXF0FLChR6vOYsqHitoFIbEoL5eelwWNdH2khqRA+Qb6K
SEhpW/y/uVXWeoHWQqE7194pAI50WLcwRH2MHpc4NISHi0hTpmpQZH+eyR6Umtenf5XianiUkP/7
AmUZ6FSPSr4pdnbqBgErubhdEGxdopYCDObPrqKUNpPaoXalAq83utgNNl3IgxNeTz+M9N+NtlRp
8b822iOmZhdsX11dwrELq4zBowuvuHEfYMGAtvr6TYoit13BH+pCCsJOlAqesdETeEQHTkuzoq5m
4b4v7fKjunevctb9LHDwSon5S9w5XY9gbqe17LW9b91fsOa/+i+XXGaSfyn2CJsn7HLL/vXes/8B
WjMqQh4TZiQMNCNRSGiqVVO6zMmdomSLj76iM5teipWQWOriU5N3G/4zXxXbaJ5Csb+wPS50SShV
FjW0wFFLF+/bvjrJ0MvtU1QGDIm7uSXu1SsJ8BLaU/VZyrnXEUufA3M+Q7fYieW1XEqiYtnDfb/q
7g/hfZ3C7pYEUr4AeR3I7P9fxn5bhbmTPPH7GYIS5Wa1hATPmC6ow5v6BDergLVtkmKQWla5G2+U
BGDtx76v2G1Q2ad9/macLidEjoAam+Nh/Hvy7ND6MO3t38o3E1YhnfhzjAyIyj45VaqGiwIJ1Mzd
DJOIgV8B8t+DiHZ9pKNm4X/kJH9mgP5ydWYKNglYbwyiIVvT8Mm49ja5+TcBW2EZ/Kpd3VxQs3ik
Qw6N28cGZ+lZ54tPp3QcfRdRYYbN1YNlgVJjSDcaEs4YJoEJsDn4pubxXzmD1diWI+nz6DlmTWH2
AEg9QttoARtgfzO3euKCiCQufFzL4lBuEWxTLW0rzJ/qgnv6ncc6mGkon/AmfetXjPYeAQKKoNEI
44zQp1KfbeU0zCmhSNOOTGOHJ+3kVKRaq85onuOYQ20ScUbHcufngGmSLavfvCkULOoYB93dKY+b
jMgp2KEWTBUXxyWlCp+0Itd3eMcNVW+G+6br0d58dlJj+hEfhyfNGI7wo/NM861CkqHmrekVI4B0
Fwz6iray1YoNV3YeSz5bnb2FqKFhw1Nwx7v0yUgVuj9p7kGXCpGBTz+uUwW7i16qW26eH6fvIg2G
7eemQMPWq295fgd2410BvcMSwhPAU9WI0Jy8keRgDESlbePat94KkGuibbGWh2AxzBDEGlHBHPU6
/f0kQI3XQ3zzN0RIyUsFCspA491PwKQDqmDHjEO+q4Ft5PlRB0dQ5UhboIf7DzTsqAQ0g9QwfAMU
4hPgQwV4OxecTN04/vw/ZkMCOvgsifA17NvYltUxiNKy4p9QQeIAatQeRgkRdjNFRPFXKPdTMLYc
R5huHZLlyJZYC2d4yFC/1DvdcxpXefDFk6iLOfchqJF+zrwBC/f5Ie1qo3JFOyjjnWqQkqrkI4BH
qAJfPDQjDKzXQdRkY2107WHbPMN/YQztLtIz+UB4VhvjeNM6sTAmdtw2OWRfLXxjTUzmz6/cSlxB
HEV4tC6yacUoBsVefMM8aAO1U8upbykCJBZjyzVIYz5VISPReTpSzXTqgr8+b1UWbAnsO9Wc1WOl
Tq1CsPKyQ671mlKGmhnzxO0lvra1a/0jtuWEicATfVhqAw2xfz2mC5LolarLDs8b0k7rstNemWfH
t7eJJvV/1Rbt7EHdFcqsNXHD1dNTt7TzdIK4AWvg4KGig/Yau1bZZSlPCF9lckkUKICfWCcN/C8y
mT0HFEjOOY+zUyY6Qwg4D0UqYEl2WBo2HVAc41Cxg0hBnkwwY0184RaqpOqlmnGEHwWsiUqSDB8j
8e9tq6tBAs3om6JC6LWeWUyXlgI2JuTcmoSdzXTGw0qk2KtWigu9RCQk4G9B5NqTZyJNzi8WKlwo
Jmcg3NI40p3Sbnfwddlrwseh2mJhG412LPprKqjUQKlGEOSxjZUMbLefnVmUk49CdzdEOlUC+xLv
N8V6IoGa7nChZ4Y3CefPE5TwTSf+qi6H/GPQSjSQ/D+Px0DKbofnMRtGuLld6IsTuP0eRfCv6Hop
OOUcrt6po8ZH3QTYyh2P7iJwT9Hrv9VRmeoGLYURAS843QMczONSjTgyE4z+Zfm9kdE7Zq4DLktB
ge57R+QrkzD4Hz0ApZ2BGp68FGqu10sToR4iqCefACIYLHE4LlEwZXC+4ZFq3ZxJPWRLFhaOQSjZ
CsRXeN5Bj+XrXz5kBaIRS5v64tdKeY1WiBVJBCCG9xDpSFw6qCui2S2q94VhIUX97k3/Nq1zCufm
2i7DnRpUp+UMiOrrp8YBsZnAKZDb/lpa2PAoaDhMKM6XBe4VcMf2P96xbUlzlVRaG4S/kyRSIWqJ
thqnlGWWZSxCR0eQT+rpRDGeZMM5gEj5rr+jirgUZpEnxZOdT8MtSITfXIkFtmBPP85AJDcw53Gf
+cjbBW7FwAQR1LsC1iUdRyZ+/Tsd0ks3GngCl+pGXnerBIpj6qHqvvcoZBmPRHLif9fjgGA9/276
cyTo56FiLdq9k6SmYQdQT8F2ySGak3qclaF1pwyoyROlQlxpsFaHUR+dE9wMRMFel76shm2laC4m
TGYnj8CL7XWGr8vB5GfcVKMHv48oegR0J3WtMykSsD6YVDDL8dqmYJatYMuQkRGtdaXzg2yt1YtN
BGzvHg701EIttfLcbi6hI4luzHFpeMosv6rINxqnVsS0Gs5uB9GDD+kvAsFS78esiyL+PxpHECM9
T+74Ca7jyKS0VZCTTRIEHpxrW13UAgNJKSxnnKnH3lvNnztcHBVLdcyXR+fcoPchTPYw9CaeOP5u
EKs+bgWwvz6uKo+wRc2Tl0qK2PpBPDZ27m97mfuN6VIx3W2/jCszAVaj4MRnDilTZwsOqq88syS2
FxadqsN7ftVLgBIRb4svk978cSvIRylLuYGZH6XvWXx+eQgHyMWbqukCs/cFM7lKoIw8oMeFa0S8
ZIuCXbExeRRfu5FnnIE5XbYTEIc++lTbjCxv8N9Z9UF7Wh74oA4Bmaa0MNkM3TbXJjb70B0orCKM
bZ78CTLtw6So8IDhCWdgP+ZJCWUqBeZHcoeiYqVUjFNfBZPcELnsnOcbp36zDmirXG+HF+v3VSCy
c4S/cSWDSIzCTVdalIxj4OL/tXinpf/k/azM2qgCU+PRzxBEmCs/FdndYJo5n4tC75miZ+j8Vwgu
YajozYaBTPUOii9w+Jo0TkcTXXAaU3UFI6cZMxigJHUclMoYmT5ImhsyhVAzDpjtkyqlPEcOFS+J
vA3WfriWZIk0o1xqpp7qm4ZyO3D5jQFdsvjyBHCugR86g6OrBt75X1wslo/jwYLhXm0yhUjp8YKi
+7LCjbDT+z8vJfXQ+WgziRWhQrdLo3PcLoHJOWXa/eewc5IxRBPzs36t3vRmvZ4JNPYerkJq6Hej
+d+tR/BGEpDLTC/1MDk9IYT2c0bu99c/ZEOEyYsFpHt5FfjbBoPqCH3eZZLsdjx2GFvTNdxTw330
FUFgGefDSx55f24oXJxhb9+zn75b18/krdOpEdjogYdM87N/j1iUqdq+mmOyganQnG4VhU3wQKqX
jCvNz4A3F5aLRodsFC7WKp8x4hFX1M1skTFiFi5xfTqMcttWDN6OMxlQ1UK6FXWCU5ddWqsAHpbD
i+blriRQOg+PeIOS9bDRUw0ZqZ/zARfI+AZXYqrrrqq+x9pzydIo6daoJZyHrJU68DAgK2T3ELuW
DeilOCGMMGkHiuWpaABDBp7Zth4gE8NbC/WTPvHDkXRzS0JBvmjvMcXR0Mi3v1ISa7RNZ+nzKrhJ
gJ1KOXl2imk9kscuZiUg3GilqNrcmgn7wQV23re9+woUYm9nRqyFXPoGoDFuO0WMk03zIC8syfxj
0Gt3Fl1o8piDP6VHYQgA9Cbr/+xsx6tku44qX1VJXTBAuarq/KrPjRffB8YNYWDOPOIiov5F+5lm
g5q4R81a52uq6ogm/r32wOWtmBh/fKehdV3vD9VvqTPqiUjceh7L2JVavoJUk47+XQyxI2mMLg54
4eKqGmKT2SxxMeafADOsCZ3Ss1GMq9Fw8XV8Pgcd+SLS7ujEXrZPj/phBvrIja+kOoLQJ6L3a/dZ
g69W282+a0uvMPo/NFGwoIJ+qlx9zIjf/nf4AuTe0Y9LZv6D3MQSbM1g1DoxQcwo+C2VT63onlWY
Swy5WFO+pL9vsULAPe1Hj9W9yx0xwu9O6tt8QXACEa1GJkXQ7ZQUHUoB25gPHuLq0jzmkeqFwfG7
GPCR6H9maXVNHmcQMHOYjQ8Kafd1RcWmP+/eq0rkUgSQr7ruAsIT/KreAUdIrnlccmC3tiGl7rXx
GpUioQ7y6FnvqQzPh4HDjglLgdTUGnVlsvsYW8gVc6aIkL+PX0aeOhlc/PlxRJlOH2ERUTOJJwRr
MRKryaOHo7lcp7n1V5Yy+lHc3ZmAek1rkxPfRszhndczahBw20YgfvyVrnb3gYcDUNP0TXAN7mlO
xl/HLQehz7ew11LmKP/5lZfZEmwVoomBLAYeuFtvz+QGtQF+qBY/VoKt2s08Um0PZI5hhVCjz7Rw
FuthoTg+w1ZUk8Aoe/p2ltYDjHF34NTbr0/I2Ck4tjR9leO+Diz7Gtqkdx1sIDZZIYuUQ1QuOhXA
yejzRfPQaliOeQZ5JzFZMvTqZ0IdcGekzQ2PWP45LKjJeHmRItDGMqr5QCqKtnXdH1rQtYBefp5E
0maKp5OehCHYTq5Ap1n95lfzisg/DsCIqHbfaeD31MbIqPYmZxqW1yV52rwU7NQE18PqgljKWbDH
o9v1ho3ZyWzT1Lw0iUT5kqAXM3p4B9Orxe29Sstfj0QHYp9//VrkbUn9EjYnssjaKzOm1uutrgE+
GpMMSYEO5EFmf1w2UG2jOcHsXEPzSzHlIp+95hwQ4YfaTTey660+RvyXTS0RKsDs/avyRvGSVZej
9YExn/Uuprwv8n2T2P+qm7sLe5msixbRDGGjy1eWKWPH+PMY3O2E09SMtF5kqETsUHIp82HaPM2L
7GdRjLmJCsjijYQntrfKJ5acBSrhuy+ELEQXhF4XdX/zXrfkfjesxiURgTIQl8+6ZvyxhSS/nPsN
kJqQ7OuWkm1V2iL55JaGjF5Vr6PMVXOnFUkHB/mQ/HQ8t0ZzeNgqmxMZp+jcDWZ8pZiVxknbYD6c
rypLmZmV83MCBbffnOHCYrb/9mC/GAkQk4Vx3xqFHkqLmaa++lxEFJUgmElb6CI/0EibEOyy7Cei
XuZJIO0ooug8vow7C5HVW/yJiYD3NaeOwHrtHxFlZU84YqbkYGZI3IBxdmRx1DIp/KJnBJ7FTo+d
Ue4XCLToI+ozdC4oHBfOxQbmt4MzkerltQ4PBg1AjUYOXEDR7EqSMWd+qzQZTL9X2x1/D810EvQJ
mSl0TVXDW1ld1wU30u0zhGXLnZSPtmINM9YWvphC0I0TJiLIKbpRizy3stqXbfyFfJE2LAwCX7rw
SK1p5kVZq5pmgHTouKp+MowfSspEkdfl8KY4HYuU2jxbwV6DFUd1H5cTpUegrhFPLgGRbmn4FyIa
VGwdrE6+7fcfX8X1QScnC+t6U6x5wepAlabDo8+xXO49u1TaPHNQp84Sd87m3bF6Nwwz70JtcSlr
uk0aSfJjz4LM3kvqnLlR/tq2LjYr4u7IMXfqK+38AKNyECc8P8tZ1RyNkKlshoPz0y/7iDdv7d6q
dWPlhMsSkJeRg5+X4TQS0uYxBRyvLCm79W0dmlhV6LoUZuxg3/WUShP6IGs6KNYrCLB1Mzcnmic6
eOiJKYEpcQCGLmPO9EFoBw8244AxJa2rDroUEyEyfYMGJa74zfN0Dcwz3wSCEQRMZUXZ4wrrYXRL
r9rawE5Oz4hqMqX3o5Ix/dSa+tSeA5lIhJgSHHFUnlDg80YzJEXWlDrn2xltP3G0mC4Z9ZRBOJ5r
bpzPP+tEPU0ZqW97rOGKfg3+k15+8lOKyGtoWg3q8tc8z7puHpdlBPjBke5TZBr9o784qBy/rExE
PtYpeLhLYRtZHfF8uNnGQJes3L5AjTDtTBF6DihjLrLtYXp3GnK85tUfo0lrOfCPO6LLE4SO9uBd
phNFU5XfFIB++0jp9ybFWkoIzU8YAWLdiIWXKZ73UqKNeHWA3YxgTiS9Lcdb6Y1riIntIK+EkQfE
DyGP9GqVQyzQZMm0x+S4yaS2+0nQRr7MSW1/AtwGSlZkk4MrWvR3Ca6srhfvnkiXNczoqqgexdyi
g50OOTVTHrEnmUOEKM2355PDygbFXHnUEtfo1u34Ndv3x6u4b9/hGCnhjc2vmq7w6vlZU8h2Fl3n
eWJgFU5u29yLa4a1pI00VjiuAliz7lGqu0XcwP+/qKozDsAT7dAACQnuO0Qa+saAalzMdfXbZHtA
l3UoU2EW/A8ZR1uQmiCXt7pb1Gx8WNl8FvhpuijODCF8fDmJLtkFWXkXlcr4h2Ve7Xu3GSVe4qE9
REvyY6TVZdbMZaZBXjlFSOlqRgQM+qp7pOQ0EOyLZZuEFUMNU3Xa9Sw75VQKre3iU252ngOz8qPC
o3x6IA56BIDSe5GTRq1x/3g0pZ/eQV/CeqANrW5CqNZuedodSi4YPmAvW27qy4knTv6oRttAbCN4
SEzY9FJe8igoIDcPlQjrz+XBBimpzYgE2p6YXQ4ekjbdoAP3RMhryKmldqkoBP7Sd0CrkgYZJPg5
PftZ9cBhfAIhHwpm4Mjf1pfr7kzf1iF8dUWb55KgjbL66OSLHIThAPxyGPp4Q5I7K9h1eQeshe20
9jgQko8gCGglzQq9C4xhFr9YTLpPYF+fMAp3EW5cdOu9TzWABRo/H9t0cfmGkwJsTdhTiiFx0BGo
8ao4wjFJNMzVjrimlqzd4NCxQM9RkK8p2lC+Lk6C+fZ719et+X05JCPRP0KoyQCPXpZiZam7VrtQ
q8ZcTeXGZ/m0LL0rA8SxEhZr249Js54R56S2Ui5drdGzY/SSdfEofom4FxJTNPtqs7hR2qwpgvdB
jAuR4wRPUwIj/b5WVVyWiMeXcbMIRWdfDsD9O4tJYfbah7yZG1UdVkf8jU17B7iAfB5T5KPN8BnW
bHF9xP8KHY5byYNnbCxol+FHYLsuG+7Q84LlCPSHAhEmIn2dYVAsTQ8aqo2se75iAWo4IvbauPE4
vdc2rTGUaaszMEgtVmyW/nbNc/1HcKGoXY+rgTDk82tNuPvhPSNgQFsv9bRhNRpZfWTpNM7asc26
fXENjx//UbsLgGPoxaoLLYUZkcluMuuFnJiL8XAp8CH78TxUCtJGgodq3sDyOrZsHpVyPvCM6RpZ
pTC2OK6GLcld/VllKpxB7SPT8eup2ylIiwfXGjzAqgsK2zbkXXGX9IaMVb68insl011+Hbsht8sX
w1QKbGYu8y6PSNZXkk/i95r8fJjccAgNkw3+pvfTxRtjcnCx6ngfVp+jQB7ujPOV3PzILf6coUeE
MxQi7irPbdPD5L1uMpWU1wnI4BnQ2s1aYvg3Qc40URJDnskGqjp6TF/06qgO0uDdne3sTJuEiMLU
hMdpfGC678klD81GTVED4fUB2HHQfy4al50wZv4dIN1UcXUYX9HLPCr2BUOVYmd5R5IhOqZFwnS2
CzklozMXUges7lE27SA6XDnbNC2BLQfR6x6SCfGXHk/njIgXMvgtoG9p7tNHICr3NwKi67zN+Zl/
8YHk1y6Ghqvkcv5Mw1Vq+UrlPl1UBpKBa51BjZnoQuzgRKbhL5CgesOr5SoI79iu2m8ngCByUBCk
Vf3ptDR/kzXBrsf48fS9V5OUvBBvMPCk3Dch7/5lwD9mXZrtrIXF/P0vvi5AGCCnB6T0ES75ni6C
HC99GOsZyr0Cf5trPtCFb2YiA+91uvr8Z3yEbtEZVQqhrageMSnmQetQ70muHsriuzb3BkXHqiW5
IT6XKeH/kExdzP/ERPsxm2cFV5SquCa2FOoZm2oeIJcW4EL7pwC1q9K5mQJ/CQ44+mYrDNCGfedV
2dItVJ2UjmKDppCFIZ8BKg02Ibgcch7MsMRRp/SjIgU5qmrFU5CnuCLzm1BQ0iLYBNr2+bsflpNi
ks0Tsxa7Ue0hYRX03kQIw3NIFqObfKJgjLb5O7493tZzeO0T9bV7vb4HQLktDlx2pck/KYPdcdU+
ijE+WePm44rIsToEsbIOexYGL4rDCSoCbHpdVwJC904P6HPpw6fw22IkwK2jT0xf6fYGwq2VwKzh
fJoJy9FKIUPmM4TtuPNJ0P+PgGa84v0jzIrVw9qmIwl6xgQUtTu6sZn/4KK0A4uWiH/1Z9X6TflD
n+Q0FhrCRg8lW7XtpYr3/nQOnDE2KrNSV4Q4eaybfl6Juf9jvQ0+tuSeQLLKA2TbDMDFk9fyhcQ4
VzNjzEm3Sh/S+EN94cG9A07XtAhit5uh97v2hFySbxRVhCxNkPCrYceEwEOvQuA2T+/d/rs8fZEI
mW2CruuJOwUiOPi+W3n8gf7PQLdbRy3JCL/Rh0Setj2/ZHGt6TMJzQxZsEOy6rBll+DzsO7nOe5a
XQiAyKjkEl5spO0Gt7qcAmMZI7Ogw9n7q4MhA8I28GWmZeK+7+uEcjLYdwiiHnnxsRAI3QPFlKVf
9M18GbybzgQwiHF7vGIIPszMODyIfzkOYQbIno0eyEZXB9VeKIGxC+ljEhJ56qeghUAmYXJvmjVr
bTJjgb8QDYnTOVf3ldX5dA4ayRyNUepHofpxCTJDGn+y+Ad+TnvjbXLiFd5ChhYH90t4xLkNTvCt
szN0p16hiKfhUOR+K2uwZQJtU0himHXxC/vYkBedm3VYTou2DpCZrh0dCiZtOYkfd5xwPiBAGh4v
nT2TkH0r/CJnFfd2in3pEKU4bDMG56wq6YaTduV8brvfKQoUDVLf1PIMhZ7u0XMHg0fa9U0qxhiP
02xhNN9nF8j8z5ZA+ePcsbo5xPO3eeR3QEIXolQbGKk/RsYQTzAEDC3ODkXcgGquXZ+16Vh4i4QO
QurvP2RQOYNHEgNagBmYih757bHY2cUmF5CYPI9KwxpjAvS02T77OtxP7XPTqBsTzrIO7v9FRJqh
loNPHxP8XzAa1AWcxhaKbbrg3h7UEY3s1zy0qtodfJUrvVRR4V/O9AuVIpZioXRC51vkUQ5+/gj0
jdb5wLC1XWvhFP2uxE64q1X36Ar+/+2+9URxuCMpC0jv47QIEof5JsBfjq/6XzlbUPeOiSR812ll
xdNa6Si62v7NHRgXa6BT7VyACSqrU8tHIX3c0Ee1DkOFoY7w1mDxm6c7Hf+AztUQRGi1mD+jv022
vWJR7/nNiq4I27trMOy/ILYn/7QU59JUnIb0vWS3/4bmdjmtwY4A+Rw9KkVZjClRM7FFUrFfhtDr
iwRDrDXzgO29XOGo5BGXp/5KOWZH7eA+ey3Z70O0SToAZya63GGwbOuVOzsc49GOH7N3XMYti4XZ
O25WlixdKz7hfHWwkUfX8vnuUhA4Fse/DtWcuAS8NLNNwMjguPk7FY7HXBVqGRGNP+OWHTx+Ee2h
wQBtEVzSvorStY6qIY031PEk1k/B1doBKDNZ58nav25F3KB3ZYe9YStrthE2itbEBGjs8es6e0Zo
1zLBDhj+NJIl7U8NmXmxRmxosVPdwI/aBRvLR+CFNU/FIb+ZwpiSkcohsqyu1HpRx2uY7dyZmcov
UusgvBfg5huvfa5Kp0XUWs7wl2sM+7moJVqxqOBMvvtWfVzFZeWYzTuf+dIsjRzB0OHZ1OoDHcoY
P9wlRdMbFYKwlSzIcEMUu4bb9SqaiRxwtNnyFGrvFa03+h5LcYlXmqf2ob5hfp9yKdW8Xys5Y3n9
bx7MUEqO1Rblr4e/CR3Wljg2/n4dhKrijE2sKCvTjr5AFBPbpnZykHd6T5uyWeunUMN1bNy8nGYc
pC80klkKkxAVNFVukXiR/ILHIHkhIpE2GMdySbudvElVXpP79JthyzB5aKw57i7pIhXvLdBV0M1b
Kb0zNCcZ8K+lH5ERig1JFXrXo9lMIuwDpoP1dBfgm63qmu14PbSRzPKZT719JxcnY2+U5beXIdYF
k+UC3wkxsRvFcQYAs8EaYL74rOjJ9p/7USecFNmonAEY2jaXUyFo73rof/hyuTHcvKTsf5+RgXX2
b+WechgGInJHq0iq4WdDVhI3Iyjj/FmcNrY05hDoJ48fpkSphi3SL0llzw9+b4ALBNnqiRUzEsbV
ymk9LXq+/jFlOjdlAMzTITjruMNyVCfUUj4LXNXFGT4UdPm4WMdKk6pO1qR8wxWT39aOSi6kvVio
vdNLxymAxZZzCDg1ppHCxOz6hoJr7bNqUAJvFCIr4/UmWVm/rYc+nrHxrvGBsazTRnAiJehtnx55
y95LO9QrH4uefFrCEJov6q7p2KeFVZntqgSIRld7g8Jqu5ZXN0hr6abd8jblqefKXUbRLFPeiZ3O
zJfUY6IReGpm1yJGfG0L4R/lgOTl8f7d1njTYG0dD37454F06thQb7z3ENM5olvu0ClUHzYw77Ih
l800d9oH2Q/4uFpbdnYJy7mcSUnwkO1asWiiPPXvXtkqc5QumzNsGWl6gU83N8DKu0kM+ToZPiDw
OyV85oDS+eMq7L7WZawqEQ44BxUlehNh2zuJjcmZPCH4qQeum+1tF3vJeOvU4bCnFAOyzVzXkxpN
GeaX5CcOsMQ0SQoZwUL1l+MhZvidi7ab44IMRZfAna0NK5uGpE2IuOBamE3e4XSVBxz0LkC3znZ2
F2oFM3td4mLmbslzYnwxB2WflwMCNbEXc9h5EDq3HNzHHKoQ5sBO7Yyq9JoCk25k8sEvLBkgkHyk
nY0LtcXTfSnbOZBv99jGk+4y37f/8ouagYLqzrrWUO8HsHdGvGyzO3OaWPBXchgLHpkkshcBfjfQ
jG0rg9XB/rugiPlA6Pza3pkYwFKUDhaobral0J85H9+B5ouf0Ws9SGkCNqn2FKlr9FpBzRe5Fydo
7LlUqRC1I9hEu/rCDNY0q2IKEKzMR7ycRoA4XOwp5mWPlWRMTv37lKCQmODWbOv2HMr5IvohuA+4
F/5a2+UfhVeHsseroPOCUez5wOHvNoEp2qJ+Ctq1guROkiEeTrEx4IuMerVIpiGLBjGchwhuO0FH
oDrNYvxVk/xDdgCKxHhfcB11Zs1tHzEJu4/nzNdBXr+094B/woDP1SPEo1fPabxMJ9XT5h4YmD5R
c0qZQlKgqOUD7tZ5gR9SbK5scnC4V8lq34ouYuRyxYzPxGeF5JGLZLv3uWIe5bToEFogFPjl27z3
+mN4y3t37fjz5LTZVH8RuGYs/bwuB05cetLHFG2WaiZxP3LcZe7VZIyoXCaFCFINDWGV37/rm4vu
NOrrGtd4sX6Ug6JOODOyj3gwaGMJWf8gNApZqvk984aObDzKqP/R2ucEqS9jUw0NCjPtg+PYyf0k
XRJ6jGJhLEnglt66CR3ne3p0jYa/a/lv4stSH2V1yv43Vw7Vsmo2TrZLnQdO45guCfD/6tzfM1fW
TF3cn9v7SR53lU4rFljd3qeh7TWyhR4yAU0rx85NbsfuMN8C5EfNCYyJATvUFQlHRgihxgZUPdnH
m1cFetUxRlZk4SjQaZL2OvdK3d2s1pbv8tSavIaRb00OgmbhiEmo6EShuc4oEccG/dpfzRz2h/nL
/k5LIw1S4mN51YSpk7zLt+THy1qQ4NW1OJpWOTr3DsADKqvBNn9SsD50pEJCbypCpQSTq2b/TGiM
FfTAbno7KFBz5grRdK4y6dYIjXRHmLk71P4+JVVr/JloScenG0Qp5Da8baAZ1+quBQVYG7P1rUVc
6Bh2JNXgPVHyi6CRjW5aSEPbhfzEYciAsXstoNM0BwgzOIyjwlEQV8hzKriN2z/91VV2HoipnUqZ
/DDp7WquEg6+EOWUvl8zKwiwsfugpUyTixJ6GYl7TMEgKCwcZhZOltMDTrqJ8/qWJ+uBMihv6wVz
2GQippxTBD6jEEcJt99sk/q4y+kjfOD+0pEZUI2rsu3kQ5l1/3wBNm5FT+1/yK/MhqE9sjCt67KQ
kAzm0F6uC6cPt7sO1/RkjGgfMHgnrM2Pkq4UJFrbM25YUPaHMJMd93LpDLtzT2zL8pRim19OOenX
RBj6nZItdPG7JxDbC1zglRwMbSYnZ2V7krlmfoSiTavxGLBDT4MVhCup/AVF8wssFrYkTj0AwGGn
N+4JwOszClckcspOsifGX6o0xPEUNfff1MWgjmoXKnxkjRRcR8Uf9osBDy5AeIwf7b8zte9iGb/a
pq/06xb1lI8pauW3vdi8SYTgm/dHfok/83OATQs7rQsY11OProAxBwph4nOK1nPSeo8AcLosLHA0
GjEHq9zGXAiWgAMnq9IqW+S72vcDYHtBgw4KNyBBb+gpBmBTysynnHTsccqfN9hPLlShuVazF+Vl
roDMAki/QnjibXysHduA8EEmxQsB3NXu1GV98+C9tswgUtlBZ8T4k2s69R2y+hyabQ/qjnkNFXPi
EL/rF8JpSc+r8t93eAnxRehsUvyZokc3LXlLkD0AwKufbBDxnnGM39ssH+lD2lQYiwax3PyvVJFk
cyeWORV8ueegES4FG55322WTKSVlkFe5u5vf1Zy+SKFR4StaWIKB9apP0nnJDFeGFDuESbQnw2br
CSghFdJE3EXGYFrv36/ojsEovo0PEcnd8i3HQnNBNN8x5OkdEGC2Ve0eHdr3gutnoJw+Kd7LBCLG
tkJUSD2Oi6rzIBDYFikzgIR4EqNAtIXzhs/XDC2jdp6nPW3Z730T4B20diIBHrZ6Kvw2jjcdxcJ4
I1sg75P6bsj8x6yJx0jvGKm3atASYk211oB3OIjPb4GFO5oHsaOpd+0f4dtAqjsHYStgd8mRiglQ
T5dI+H+WYMyxElMPzSBbhU+0XYrqAsYlBGOA/poP6vHuAKW6aM8pNSGNKLrJk1RzJDuDS73UL0oh
VYrUWvv4XThKIWpaCh8UNRsQJQ3vD1o36o8oo0hIO/SRhHTlFC6x69RDTS0z3TnhemC0kaOJLq8d
e7gkPOoiL/KJdIF3i5oXcW8YXoPSi34gMCfgWf4GbLqgHoZLq5mbFHV1R9rSLM1MZ8Xr58aFv01f
BUn0UuO9kkVCyOY04Nh+/nTioC2IppLMTRLnBB+NPKal9Bm8+uvopK8i8TqPR6chSdsj6lm4Il65
rROUS02q+/cW6KKzdQsKWk3RqXfpKrClOICH/NvbyK3S/53okvprU14oEpMmL1OnO5RpGXvtrHbi
Z3eouHiPj8eQZn9glFA10RTp3dT6L6TH/37TTLMj2pmX0ib7oppsJMJbF9TwHJVsknTP8vC8tCqO
RPYLmbPEyBiKzKZ4IVlNQ4hxZzatzXwYbhlGUOkiXZBCVODCRm0sSFSsEto0RwPWNwYdIAF0hHY4
RWlg+RfYrBYVM81f2AxHpuV9XTylAFwuEa4FHnWNlshMqqZ6vU/SNojXIrfMzKfeMeeHmJdhfZhZ
JdlVj+cRSXEMlBWaH7nFWJN+/vewT7GNvBBLbXQ3AYqz/iqUaofkKH/XMODAqLEYKAl2+GdNHuTS
fGUlroD6lOR8PdGLBdQ+NolsR8CLLzKBJkLTigPaNL/eNR+zORAUKo8rzGptcIJXKHUbqy0rgpE9
e1z4lRCj0orC9q/T/xfeYavaaW++xgFg83ZIVyYVxzvpym4xutvMjiZZTP7LDB1zpbwpTLlzeT6N
VvEyAzrsriwzr7VxKHmZjHNUezYfeGYz6fQRKUbdjKAjs6ldkM2BwyOEV4WNFw5/SmTGDgM+oW2U
79sDSKbY2MF4HHxuZ8WhpW2Bbsfd3K1pbbjHnVNgivX+HRhIsJBdJdNk8Ino2LhcKKWfhzwYrpgb
L9zjHXQuWcQJccNDnldHtqNB3pcU6OogKF4Bg8SJZCwsCXWk4wfwRs8LA+fpB2gVEx7sa6D6RcME
NyHGE+oJz4wleT3mOIx5VNOsRb6gFEhmyE05+7Bsdeb5oQ5GfGvUoKI1at9D4nnml7/WqBKdtK87
0PzhZjsDWNjM46dCxsDqzHl3FMUo1U9J2dNT1zVOP/ximKIg+8MUL3bmknUqq1hNCDO4jtQ1Vv1E
qrBJKQT3lNl0D+2nuTGBAeAVZ7TQNSgeMf4OdH2/tj46QxrqUI716/ZAQYvyDnDOR4ginFREM3DG
4dsapcjzhZLKrDhTDA8B4CreKlgg1yP44+lOKYG/YeTwnCO2ghnDr1+QAapY6SSCuai3PSlSPOJs
NpOO8pwpClFaZ+anClTzbfvUzONaCxhcky6SZffNc0E3NVY0L1HZ30jb0F/90sgfZ5PwBnnmYQaA
Qvu1pcHHG0HSNLeL+4YujplkeaRmW17AHdrY3JvUhduCwumqcexT3/wdxFwhQUE8W46qWCzsAvCF
mttXe9+rrCluQ6JaDWeS7udG+K9uP6PdVpApge3PDxxNCEXAlM5k55dHiuIlc/y9nzpPeB3ms2pN
F1MIjzBZvzMgyBflU5N1F9mAtky1mbXIQEL5a443tiMg2U1Spaw6+2KIm0GA+ciFe8nW4fQWaP7D
HUASs0VOMKkSJLvmENMCiO7PFEj5MRsKQ5kB6hXy+tS/Ciid0eCi5Qj1HoiEw+tYE3QTfPRUPDAh
8SsaC5qXe89QClqO/7orWaPNvs6bLqZyaa7X5WjpyYH2un6lHjEgU0vjq5/JEwMbB21djkqzuBwG
OI8CdAP4bUW41ueTYNA3d3Z5H3Hh96sU1Q1UJGAaj+/VARl/IQ+UE/eP21XIufNqhUA7fDxHwDWA
gmQ3hvD5XZkY+4SDQdGZkynwNmKdyp6gKcwwBTsiCxmVcgxFodgQEXZdreQ+YVbsNEGeboSF3jem
l3T9JyGDVtEETP/TLKHy/YWvxwSOoK4g+jTNFzK95MexGyoxdDZ1XA5M0zT/Ou9PvPEuo4ytc3hH
lNnkVPmJNb7kWaJDYVBeOsUWL2cimKXbaFbhqyb2vh6mBGURbp2XSOuyNevMq+qDb2/fJvGDQevs
hfudbTR3Ue5gnSw+y8TLGJ+36aLqgqc5mrpHtYRUuhfxBn+5atZ6uXFkn/WYEKU/f57pwUfA0Y89
FyFidQFPrOjbRSgCn0l1Inwm3hpCJzn7zCz+Z5oi0vIrRklkuQ1KOSsSxFXX6CUR8qmeJkMc+Su0
69F2ZkZzStpaFtz9xr4/uhDZyWIa8qCPjPp/RRDCST/F4462ZcwejMPiT/YZ+dudUTnZqknZnlST
j2vy0sjG+S2MloHCXCC6Q4LVSMQ5dz/BEhMRgb5WusMA/v++LWmJFoXL+9RfKD3pMYVPyl6kI/4m
bqrUx/MjWRUVIHwOAbIWaIL0uhw1bbcd7aons/HtWfZYfSbtt/qMgKwzM+THQuO9Q056lpkQlSOV
yLl8Z121gACSqeWndJo/SnuURcHJrSCbnKyeOwbDloERguXjk5YXq4NAmToNzZp1Kcb5tF9pgWwa
oBbXbHkZd0DsBBhlbYTxBB0NVz7Y9loCUUTjBVYLE41gbIXqTFr4iHjgnb1FM9+q2JBWZmV2HLLq
oJs0U2mUSmTIXr9ByWgv1S1gdMtPDck6V6sGzQjiaO5TIMSqnuRk+bCHFRjy9z7k27UboSABJBUR
lmBj/4Ib3NkdKXfbkBvxwiomgiiPQ1z6rK1mDZCypBhtHbAsaeue7FLuWHjRpuiJSob3sHLNhzce
d2Q1P+VVb97gOkbqc8g0xFH2DIK2Rd7dmGHH+2qQiq7dQyPJtBb1WpvChSKUH9p0RISVKMj4tOMB
A6HehwyK7Hjbiq6SAdrTE2I+zsUbPuv1S6Mz8wZ/YnzdVVRuI6Jpa4UYWJAZfwwZ5SG+h28nrysC
ng5hdtCKK8XfiMiF/EEU1jrhGpaexhFf/g5/kMSCV/AJLeUkEFiO3Mw3/0R0Q+2+dStwyrvoNRNW
F7lfCx7z2XG0LIL1BWqvIPl0n+cc0hOu1ARluthAQ+VWMVRORKmzGm06xC6I8K8W0DeSNG+1KH9A
KmYHBg3x72cYPDAZ+X/YYh4twX+0BNQwpBS+mVl2LFUAh1Eky6sTjEdCrYbQ857YkeohyNGZZCAz
vktHuGefkn7DQ1i/HLX1xRWeStmh6Dw8rKmkpsrxL2FAboAWdoxaJYEiqVbAhuZoulAaEFbjq2Lq
Yx789SXqKja/m5MYEAVE2mUDd0tzC7eIxY2+Ey571iW0Jztw1DrshbqYQvEFcljMgEt72W0joKBw
1ip85o2Ip18PJOUsHFaLX0pM0pCCAecSuYoQrMTr6l5XXUT4bvzcefifC396oYLcUNR6Jk+/JF7O
9txGePlRSikJOoxkrXjfzNQvf6hSFK5otLBO2CVcs67M5DQJy6Eqm1bDVWNtADc31D7cqY5FNG8b
zN+oGc98SGrlSyRGkc3ObTjccMGnzpgEk2CDsYzqiuz56QmA3+3RhBq6OkYIxZg55ugJAUYi7EGo
0JxZIBsPc8/IgM3Pv1t26R2I+nIS9hqf06L6Y8YJdc2mvOZbeAfcAOWPhD3rWUuukg6Gs1qijZ7a
++1hUHdiLm6SP5LfaQ3lNZU0SZeKeUfPBqNUDJuP4nPw8eliVrhYPitGWHKX9dTE9fbYrxf9+0zQ
bcACKVV8ipFIEHUqC+uVh9UJfqYBtv8URl7D72IopFCY6AFwuOunqsUDpbMz/sNZz3HH+6n4s5Nu
K+h6fIVH6jhtaeAsi1CejcNjXfmibNkte9LpmPlQRtnX0jQDi5T29TlIBXwhLYd4GxBb+Fx4i+IH
uLom3nMEnwehY/6OPCwhtnvwChI+09xep4UsJKeFhcd5Vehfewn1bvNUycMVBu1Ss42M5W9aeI6q
QvOwGnPqS/FKS6vyGjSgs9XSnSxD/TWpI1CHJau8FCS0v6m9vI3ScIDL+Vi5MdcskrzQjZfOjR64
a7571n3BFqvYwzvoYwlPW9KKYwlu6P//upYgaqhL5cuaCCslMFkcnZoK+HI+RQbSlg46ExDznz2A
LQG13rORJioWJJdes/gktfQuWQe3ed/ieBjWfKgplTf3jPcVfQPpYStdhldIE3BoXF1v9mucqj/c
DxR0NC8C2ILneMPYsB1frdH/HtatiPdW172yNLr/MVngsOmI7uUCUQumhBbI1ssGajtm/RrS3fyA
wtLGWiNaZKtoV2cclsgVDmu5PChCmIHOMpXsu+DPY6xbR5MUNGQ+NUBX2DkdPyDBomm6+n0mtRmM
Hz9flKSwz+BltVnGiSY6fOcopTAfVjTkhUbZFzmag5R8ijROk39v4H3KkRe1evw1WtG6e6c5UMTr
B091Md3p0io3cZ/ZfHhla5zDkRQEJ3gs0fBL05HhjOvbyXmJEYKwqLFRdpTy9E7djdfAiyDEelWP
NqGL+9RdG9qmu11uA5Jceofemvr9+EYyZFDWFyNlG46tDAQQJxKLHtwcI4khNlwFNigxFOjEwwza
66kRIJR4QA2LWlkupDzgch0Kr9IMZ03vYRwC5WKNkLUbJtp6eZz6YOfrVV84KkI8seZ6f2j/7Rfg
2c0Bhoqe42l1MQaa2YKvQZUj+r0nwLogTmt7p0B+7mEy2c6eT5/P6lAZWulvm555FrRhyWic4pQO
HDwjdKRHnm6jMJLJCVO05Vdz0/ljCvH5ytpLphXaqEHoRXtPDa0FqV1rde/vXi8XD2fCn5J5rsDM
UglpfV95vbDj6U2oYZfJZ2nBUc0Bch30C5B06435v8jUzIAmuegCcpS1mJOe6Px/zaGxKkHKy/a5
CbNKoRXWITGSfxvyGbcfHdN7HcWkWHpgMMUD49f7QiBYn11RHKrLdq3V0AM45YPwThdjKRKDx6xR
MAkkt79kwjkef8PFhO1K7bbIt++CSlVo2Pg4RmYW4k2+Ra76/lx6CXF/k+ve2yR4F2wLKCKWvniA
B95Lgxg2gQEg40xOrRANZZFxCvGazPS3zp7p5jiOQ/otCkoBLgRlrwgkYDz0KrnvmrClNluOFdNM
7eN8ykBMN/EMiryqvIPk+ZdDlrcUqFv9iMJddBI7Ghgye1vV9kavKwb4vwRJPYgvvaqJpsCTvMfG
0akEaSltZfqreEicUMgcdwA65SXk4PZ8xOsoyFJzKnzFklBTxB40B4XfgQ1VuK6dRRK77/C6QDhr
71C4SrASPPoJA1ub1oFAPSw2hbU0OeZXUkqGByGfPk7FdPB6hPT8y1pJ2VQzVw63lO85XijeUv21
UPt0DhleCGR4nQuNDt7faxx9Ta19qhYMkl3m5KjlcIuG3s9nLE2NMl2+zAAZ2VmbcuIjIp0huiQh
GyBx7atXq0Nc18EnlRT7+TBe8iUkn7tN5WFw7mSwsHW9w3LCg52eQHmPBmc5nexM2JE1olIZdIcQ
GYSdLk4+TdMx0O6KlWxQqQlfu4v49qf+Zvb7PK5tqobMM+85jQ7/z8uD36AMyJX5T1oq+gCuSnkM
hp3C+ydSF8cvYV6KZCapt58b+P9qVpg59Vh41/cFTzkJllpD/kp8ABp4M+NYrnWNMnQfSOhj1gaD
chSouLBR/7K6Bx0IeSKLaCUpIWySExI+i2JIT3jN4IGWhcMyrNGg97odBIO+NO7H7OOPW9880YQ8
8r1Lh/2sI3+Rzz0WgbI2XBhiAFGsyZe9RU7CDaPDcRQjAjsqrSLDD7kiNHiTOP+wTlPIz8TP/GD1
s5DVHAHId8J3Xngh6wT3vi1xM4mYI3QYfwpkLVGrAKeDJQqnN4LxCgS1H7N1XMP31PBB6bgbKHdD
0yZeq+qcKkWlq/nQUdA5A+n3kOszrBNfc341v3wvy/2ruvZ1T4A6x9zeXmcFd6wg9oz6splN1pXI
HoOaail97c3Y6/FNmV5L973w4lAQ8lUfJ7oODwODOEFitBkuvZS+Zl1b2rVQ7JqlwYL2uhXZg7mf
9cAzqcwqnFSIC5X56S3+ObQf0hemptH+ylcqfk0T70MIkxX/ye+meWQy8/Bkz7I98hYxxTqOZ2me
zF83CvhZVnBrrpc4QCP3/jXFynATqr8vepsUS8lUuGpKTUhbcIXYxwgPj8K2ywZ1hhBcoOrp33Ov
+i/pZ8BuzJsJRy9zYgfSFsTiHNGf9v7/2CpNX+2rCyjNbx4i0ulgQVbtm7e21/jQZp8FXRwrp8HE
M11HjqNRsAoKlGf/zU4HSZsV9NspJGJESr0t10RBNIWSaR2gDolcieeSUgDrQvWGPaLU4dJz+/qd
HzAjqnUBCP1ydQuYfIrb8msSgLWM8VaMZ10+aNzocSnfIEKgjYVCgH3F3i32O859AmU0JGxlWy+/
oU5XdxKa79SwVvNt+Tup524G6k/Y+IKL+ViVuiQg5MNM6FQ+Vl2AA8nu7x9bk5+RDqLT4aUj45XJ
ijQD8Dxnxh//zJ7MBC2HXfHpV1vQSTGZtfpiYpsdJUPjtmTQZjxExCzeUGhFc+H3C2XQRQ7XC/yn
/oSODAG/9YN1vCPPLWCkn23hjfcu7dPfhnQe4HaPx9RLtxzkGlJzM0M8XQpa4r4xVPpQaoQMj0zd
Vrg1qsNp2j/qXM1V3Pz4hMruL5o9SLrl4Yt6W6Jh2RfGdnVPb5uLKJ+QHA2GvAVOn15rvr1GN3YO
eX2U+Pi/lMytxkuwhTALAzVsA1FsQjD7B8QEcOFCQDHJ8zwIL5DjWAenhZh6YSNdTd9qOQ2JSngi
zCNyOzVpM2m1v9lIfq0BpfTKeMHQE2H6rSYGU020EXq4Om8I0t1eAHK/GsCPGJpQ2KtJEZMvHvxv
uD3XMXwlZ5QVED5BhRbO7CUUqS4Vl2MdAi6jBQwsp3WiIoqg6VCXB6tSSh22Vbh5IM5IyJRtfvgW
m/KlQWlYEISiI75+LVXxXj102oaGDG4rMrVqCMNpza853pkWvz4avnLOSfcvYgdJhhfegvnWOW9u
dA0m/zSbNOpV7oepAa7FEfFXCYb3QL97S0HxtEUoAPb+8KGN0c1a1BZ8WsI6dYzgTOVyZ9HXVClZ
0SNGtIR3y1VSBTQ8dsmd/oFkXNjkcLKHYlFFTQkAgAtJGFiYPiG41UXGqpkYCEgTPSy8wnHeaBxY
VQt/SyuSMiXoStiRBCUj+Jhq/3zfiJwCS8j9Rn/etVML1kJR7XtBQYZQ+tRcFnm1ndhrxeD2bA9T
aIkwUU+/HlLQkYwBwxkYHmwMNFOSk0abuSW+3MneS8uvfM+YwB4hXh29j/tCd5E9zcCFZTd9I//c
ZQ5+epx34YJGD+VQ51Frl27YGFxxtacDqMRoH1Oil0wtYGXl7Ij+zXuUgGiSO5iqy1qcNcz9OpTh
ZxRChAHfK3osERi7Am4fGYSg8C2R32dFjGQ39vgJiNLE/d8iLG8ucA2jseLBVA4UzfBNLS6wLUlp
WVX8qHLIkzhGrjVo1SfZWq7f/tTQ01+gFyyHsfCAf4HuWNKAmq1uT/76ozN8/f5e5boFzZeUn4DH
22vpuhA1EDqLrtlkYwegVeL/FAcbzb3VceRk4/YIwlCmKNfS5cQvVhw5z2igVo7kAyvmvB2QHDcX
yN2PJzdM7wo1jA/2AzyB259vl76NOteCyblBRy92yeIITg4HS5DZylHnbcBM6VqYzBmHK98EkQwe
M7w7g97ZSSbe5TIni/uOZ7cQ39yclbXi4HCJEVeaTnbg1OEMr4xd03aEW8IX8ztFTyWIJyHkpEmS
S+3gv8Ad10yl9/ORH43m6bxFRWlwVyUAPnyxWuEc42iXAayaoME1BUkLAsaactjZty6XXFBGTtpb
nDnX3gjg3EGuqP/DX3UPZmbuSH2P5sEFJMHI7m0Nzh7qx+qTpKYz4pqS49CLI46TvXgmPqNIocBv
9T8ohXSuuDifBtAPiOCQA7tcCO6iRQxEpDfb9bNI9/DARN12Qe21FBsUZ7YQwlU8uHEKkysZg/Hg
GSNsCC4IrRssseZEhQFjQlqxZwKtR6SWCFhYPsIIajUxTLjFWAXjONTILG6nuxlyResI4Af84qra
ay1Yfe7Rgc6MIXMIxFz79pj6OS2ZnNT2iCAJvQgoA9+w9tQ4sOGubFujKbq01o6Zq5PwpFOoSLib
SbFkI5rEB2cVCUFv3u8+JyXmKe/NM9QHDVYWp4GUUM8pzDW8kTU8slivKeB81ISal3/w2PZYFqjn
fUUQ1rn1wy992I4crp7F7myVmNehKs3OSkk/M7uNrc0hcsiSD/flGXoFdu4wTNzQHdbYOLSt7GBc
o8Cchqv7RRuHE6JL8rBtEzZ63ZvAxYjFk+HWQvei+wGPW0bS6FFNmI3/PEIi0QYGxXUdKNmD6j6U
zwrvtnlTschHADE3PLCiL1QRDN4A8JjJ2hXa4qwJ31tFRs4tSSiOUVxWUn79XzANDR5OI/nblhpp
3V0+x+4IoDcQj6DmdKFy+kwaaOjbVxf9gn+7wXtW478u56ltigDzkGCkkKEqCo7Z1xFrQM8y84M8
AVFmep46z4LpkkaAgDv67U1VkkW4IZ4OrLyeglVHYGs5uv1WD85kXdsDeD4nJehv0mK+L4NDUYA5
sG4Iswtpa2yj7iusSYVolzcQ6EhrPNCZi59mmNBkeQSMJfyNmK21ynzuKI1jnMiJFxq3OTZ732+y
1N8It/k9FgZX10Tbtak2xdFENLa3ZPxBtmDmB8R3KKZAfMA6KR40FAxyEKSanyXLzld4gTbc9cEZ
8wEE5zyBEVNsq+MPw8oLR3i9oDBNMlto5dB4bR+MP0ulMEy2XpfPTkifuqxUjhzQN5iZEh1fGooo
4QsFkjEGAQnxeC4hAfHmXweeif624QSplRuLZoPVihkeieXV5PfoWRXnb/2EcHhI52tb8ENTPwv5
EWLxHk+vYFXekSVVGbW53/VOSLsBTSkUR9U3+MmTYRQRu8iuveKeP07zoi+ei9HiueJuq+AEOWE9
1gQa8EhRJQRxGU3/h+Yj8V+EHpkcKBS9LOLFSWLs5ORw6tpN6oH3r+Cdu70WiGt7AEZfw7OT74Aq
l2uvOHHsAVv6qo7RGdBg5K25i6JewjvAdq6yckVN4f+GBBkKBGcxLZIRj89z1Wy4HA53+nYWGqwj
lzCrulS8RG26TP0unvSNGPkBMKJ0g1MP2UABa4y/bRg100LCpY8W+S6vBrt6/0bg2T2kcPN4gNuP
30+F2cOlCSCgZp8KhXYzTof3w61+Hl8JOqErCXQE79i1tAzk7eG8WFS/bmtgfmYSE6xNy/AQ4Xfd
6JMamQR0rm3ezUhMJO4E+1IEFae6rlbp/UPFuebo2q2BGUo4plwMyB9i1zZ7X/2YUwLGeN0/W28x
dZN//MVs987pME0BUsWLxFCDLZWV/N9GktMD+5nCTtR5mRiiCuT3LmThyBpebK27B+Zg0l8xMExP
51HvpyGHBlR2Z7xzQbc/5p0ul+HbEV6guh9YHZk9MMVRu4MiLe9vMCzTL3ir4idIFywihE+5nWZP
NKkYxr7JRSREBaUCWwFwjpczsGcF6fr/Ne7cOn0KeB1fk/tD6fGItW3g8q8aD/ZEuuOp/TSE0Mt6
Gf32FZLBESq8WBUi7ye1GpFrFLZaxb531wNlUnXYmjjxPOCSVDDDiP7FHlGkobPZQdlWRbTnZ38R
AJcdzwet0L9RwVQteXfmj1OLI7z8GVMe3EYDzqawi3GGUF1fX3Z3tBjEB8VHEFUVi5Qlafnn6Gms
F80waXGUJKUsau4RQt0kX2p4i0nUd/9zMaLzAFZKQJPtQ06pKzb1fWFWLjKs4/SXljoinrdkufQR
kbtxYDanfV95rj0fuMsUbzVeW258e8b27QZRKxJCysVy4av+gdetef03PJCDjffyxP37lnaxQo22
4lD6NnehmaNgF4LK/0eou89jOAW8vmEsyTwT/8apfqductOrSB8Fw/T4C9fP73ZDcNWldODUm2ZY
dhHWAXDELEZpGzsQnRC/tXbU8vjuC2IyLRLMUHfQ2pK92QoOxZxcXh5uPHugeCGn36xsSZAjOVTS
WcEUpB07ti0Hea9Nek3fG/reqw5Wx9xVdhWcoAU2UklMOlFVwXTNbyOpGb62FTN61/AnvIto+gpR
KCalzbdPuVHQ1Sfi2+mofe0+9YiBj4QlZNpgPhJLJgWlEJLSo09kz/VNw+fQ61lxwQeEegYYewj+
TZvzDWEGjgnSD/DC1bOVldwFNUDuVj7zED2tqzTdlYQeko7JsufWlyJ2GTrERBM3RLH5+LEFp5ZM
5Iyc2GrWQtASazUo5lNbhn6FqRahK63ocZjn7ORQKUr+IfceDbSoDapDGW7LR3m3slDF9lFQUTfP
bIXCAU9TbQ8kZ4aHIwuDhKkU+KxH7lXtLQep+vaW/X9AInLrXk2cfKAD5JFEHCH7hJGgN08QxG4e
2Qfsq+Fb/Dd86GQTDJNRVWY3aZdrDHe8e5LsmjC3VtQmK3HA2VLLBRXPghKwE0eKdWSi++3yA9xs
1uTCiw4te1CndvCQd6Yl4pEnVFZURTxz8axqRIVt99GenDi5PfJEHL4J/DTozIYS0IPWsgU5Vj1x
aMlTiQglp8rKw645OWZatINgrHFWjmYJMKcDEk6z97k6VurFqFoaUHs1C/yiEy6ZAHassgp6HyR4
3gMv48pLhr8BYS1Rr+LPT/2f4modQaNSwUrzTYdcySrF2A4JKaHxeoxZOD1aCaiERQzHgNQX1iUl
iv4hGS4axynWNRftgh7DBCd9ZmUrglnbO66/kMWAEKhXObJC1Mduq0seG1inV/WNtV6laUNENGiQ
QGTc91n1pkTkNcrpHc088azV03VhtTU1VoPvkI6A/6OcNI/wb/gkjndVG0gWoKz1iK9lm6ftsUgN
x206RR4rMOMCbhfZiuJbl3jeay3bo4Wtczn7rsWgEa4UjJHBfW/fjtj7mVcxtJPBxJ8QKIKssYIL
NY7GU72mholk+JgBB6UdygRehCaRVO445IbGipP11OWkZKGOtep0qIpQfd0OOWkPc7EhTZ6zIP9s
xsZrf1tVxDe5Azh7hvtVYrPtmSixEYe9gkjEIqnueiOG+vd8r8N5DjrxXvwJpksrRF3UuZr2ox5K
ajLx+cdvPbsSUc+9U0yABIjFfkB9JJVvlm/9T0WZQf5F1U+1PMGzqJZbyziX+CJXJzpz3PXZZI9u
5H6qz5D0Jfh4+gSINxYdxr3gXmatv/gPaCbHhfaMolk/0opXUmj87Pro2z227F1+nS9Gds34PC9u
9N7GaFXDwjnAyN+eIohh97MqB7ph1PnfBqpvFUuS/kvfqJ07KCix/Au5BSyfXOTnnZNVWgMGGuWh
B3CAEeN8VI83jL0uVV4INlyZL2KOqYgNYQqjlacnM/3kRolvaaVtWJBtrvcSsuSaTQ6imXox6BAD
lEmTzNvRH+HGKjayc/ihrxHKM/tiia5BEvCKQigiLd8lfC9r494GebZOyNVs7Q7LbqPsC9cA++fP
j1faZJBXEdeneDAgOXPBwcHslyIeQa2JVKR/mBIdl3Qc21XqGuw2NnBU9XDHTIaARWNs2TVIpPUr
f1lwqlU+nNbl65CZGLcfZEq/0zA8FOU4PioI2UA9MfuOF0CisyZq05RmOhb4c0Y1KepudbAWofbF
6aserbEqjeJLzzkH/5275Q8UkH0b92/fV9uDGVskFkNKF4T6kkzHe7H8xxsd+bRFdok2qka03HY5
4L5t76bU2+Dm4FEIW45KP6/v5K/Upc/96N94md2tgdycw8+TziWhaFLBha+IJqI5JL5naWEbiiq/
ZmcXaOCJ8WfgX5VSnWTIKZ0AzJfSiBL4/IWVKq/5e9AvvQF5P+eVSVvp8iUX2AbTeNMGDb1N+y8P
yb71jFsKSCYBi+CKD6Rhmp7soYy/H5vKPFk2KghO7J/vz786C2ZLQFLmer6/RQpM0rJ3n1De6tQf
tBgCoeHrcmQ+ZBi2LBhZjCjdf+8NxvzXEWuC13tDT3soB1dL0BgIyO/038vQW/5fJSLEwzmSraN/
lg8oyWERUTt/4K6Jaqk7E2zM2Uq7EQ1jUdB1pdfWcQq3+qTttv8p/kF7O0eeeFbV2K7DrMnZyGrg
W+8wj6oTdzf8kUFeA2pVihv0gw47b35I1msHMio1LywLiSTLE6oTAxzzW1MK05SMs6iaYSQb5lkJ
N536N8L6AQU8TMgEzuOa4wvc87brPkpskP7jw9XfhryU8Y9BbNyXWwCikF8NEabSUmzfTCnzU/ta
pHzFB5vVxv5YERdlMNIZuicXV9/pVLrwn+exf/3PTOGW+BpMJoGJ6Lh7jNJiM1do6sCG81ACs1qE
PpPMpPbZgXP1eaItbxmyMkKIT+g+IUymKBKTsoyghy9THjkQqHBubacNcGhotpCH0azyLddgJuXP
ec6hJ90XhMQBtp81SF51fwyAQYvoNF1k2duCOJzio58ne/COew8NV2uNVTT/YvW9bmIGlTZZ6zjS
+uqetusY/5OhorNhpPGtNBRkmQRfA3vy62/WOo3CBtPPZVjPxiwK6cQXxMNx9kDBFxg8ojEqt0sc
MRlzrjlLrFd9pcZbGhiiDbKpGBG/56PN1o3WkYuqGnN0kJAJmQanv2yWF4fb1rPrlaUu6VEUwXd/
3lPfxJD5JE6YGuFjJ9FbXuyw5HyZtRf/7ghbW+Dwawr4ywDmHBL6Nyc/eDWvU5A89elPbZwXAoXX
ahlHfYYnsIl2EQRgZI6oluOXomZauawv3kisFjXWrO6s05xLrf6MHP9OI8hQu+1RIFe3zV1kE4Gq
3jpfpBw+L+634/VXlXrvpnA/1ryw9/ckhPOtO60MM1dk+e8bKxLeY2pWwZnZmHR+jkkpV/dtO74P
rCdPjEUt/iRJaf9seEC8OrEfk/3kKOH0D9Hoy48hPGrHiIOXBAH+pqmbIHiBCa4xF3qAfSWLNIQI
58eHGFf2SahZTXtUE4DsmWRawyMw/sGj9qqz1Pjbn01oIcl+FoDbLv9iZfD/mIpGw5v8WIFrdSOS
ElHMRC+MaIgjQ+Kmp70geJrSIfq2yiR1OZ8yTSzRHNnjmDauwsI0NuH5rUe1U32K2qM1MRTGEF4j
Os+f+d7Oqe7eOzDMfiNwLJ3HBaz9UTEDz3iX1bQpAbcpF3OMEQnzJfutJuuDLJVkN4868vd4V7rV
8qzXpsFyotYY1Q2ytSnSMDi10dvgt+P0JX2bQsWPAYQs7BkZwtG3n5ikC4iUF2lawfqGv7zY0VK9
iz3U8GBpsdx9heqU0PmdvcZZSYZtSC0W+FdF4Gf+ipVzaAztsJxwuN7qxoqkD+HUVojMOZodLK2D
3zO8TiDM3FVhs3Gjy2+a7V10DpDPnNhuTbZhPbVItInnWqQrfkzGM4pRni6ANcVSF/v7uep2eviX
T5cf70yuqMds0VEco1cJ154QtopGxrQ8wwUBN+V1/C6lmpFX4VEQP4n54GXI+FAJ/eiQOB5l4zgX
EfPM8ALhB3K8RhQ5Uc3TwGBdD7uVdSVEALsW7jJzyzGQe0hymFGBxapne4yMUI6sasAFRnRe1vES
p0r2g8WjLZVvFVpRdbdVNI5gZGYLW51tPaWMACNkv4MS6cP3ybRw+E5oGG7qNt2e08xxRIv9P4E3
oplmwdopWzdOa29M96nS5QROlxK8KxUFhOKhIOO5BpGtnc899K31xe/73qRlbtNvtohBV1612+5v
YRuMTYso2NRQJf9d6XiDggZbR5jLRlpnoafS7G9xQ7u933lazknozyV7fOloleEgY6XOzzkvXi6A
q5BddZNAOi5cOGVdz3oqn4EO+UJknrET28QDHOcjGcMXKI3YaaNUay2FNHmrXn8PG3XXk7oehl4Y
v5hqWL+rj00J5hb/3nHVkI7nc7qbc9PTdep4PDDGP01w1J8EvIxxPWHeOfDbEBQ3YxZ46yYzcKEU
9fS1YVszikUEJmXjjwad7lDUgfcxMgh1K8BKdDF48iPpYLqsAQ2djLYsU2c1NJ+bd9u8gbqzxB1K
xqn54XhOTN9w+Qs/IAQlA/v3plQ1tkIvYz+l0+zUj/NlX0GY/0wQNEWhfZHqWWqsi1XDVEfiXEkh
P9lx/5NLp4jTZZUd5a1fNexraK8Fbz8m/JC8qd3vixKhSysoBZbzTGDJBzPbjA0Vkod4WTh8SkWv
16ebLHB2BDZDnFyvvYhfeo185F5o8Hh+Z4bWGvTjR9lbmPUa3VvbUztHYgIXAPReLrGDVnJ6HcRm
K/Zgc9i/JDNMkT31z2aoiUoPFiMeNVOWLQbrRIleq+aOSYO2BYyoVqOGUk5dNMarCjcsbn451HuA
DDEWVu+SY4mbVJ7heMtpuSE7HQKV5XQPK8IE3mYU/pBf2r+yL2MnnFZiUrmcIwqm+p8DRV1/Wl6+
N4LYD5bcSXMABSSysR1oPPIGtFJmwXZj2fwtAeJ5HX34JYTq1pWYiQCb0WGuSOPXFJb/dxwVjHAm
1pLOjAYWG9lrfQ/j6ua8yIw2uTo5FQDNkzdiX56hk6OAEdGkomyxd8ChL3rwf7U+RY0k85cwvaLi
/iilbITpBpaldCY0c0HloO/L2/ZT5sUlM2apPOH5Pf0B4st20K+NC8RPVskcTUvW4TFuEXW6yig1
x1If2azkq4InTM1/VzatyJIHPBuGp1v+t1jMOWUbwmCNHecoeGoZ7UNlbcd8yLfBbxoBc9VHsoFg
3FlvwDZh6PNoLhreGhyUir65ATq4FJIgVYflfGaonCPLJBC2e+xDXDGg1InD11CSAdI1mji10E6K
GoGQ3Ae7vhsPccI/OIc2VvviE/106ym/k81scMRJUUUJafkSQgflcUA94ZDQ+z7HS60oe5tDerk6
hZ3msOGhiFd/tHLXAvzAiBDeEzYJ85dZnRDCJtB8OKETnYMFcDkgFI+7FscMJ8KtA9Ozg9iQKJsV
X93IzmhZeLrUU/flFhUnboYOb99afz4AjSGVKdmx/q7FOGoItVbacjowVJeokg45dpiNolki2gjV
9xGMu5dI4SmSvdp/8Kz42c1OTEiCUmJELxz6RbmpfLS91xmU1YprkRfVkAkoy/v7/mZPA+8QZUUP
nvmkpAKXp867TL6bqMi2mqlFAvy3DZU8VMNG6D1x5ZO0iJHHRK5mA7DcHqGh+rdn7BmlimL5Eano
UOn0aXiaU+OK6SSbqbaFfYsd+Wkw+2kKr0Rdrth+Ydz1mxQRwdX3UC8ZG7WYZwsAGKMsiO98BETC
XpqA3NgbSu1ONrXulPr4BmgBBK2N0ofVWU0vXI5gXsATAIxt7XLoU27d4zk9YYKdk/rh6qVqN7CO
y5LMyHEsmiyb+NbxTQdNHc3ym5dT7MuDzukonmpakGtsDyZHE4c23ZSdYCcBsu/MoVq/ziJ0vsbL
NZnEMzbJOu+mVvhmzNcBSaHh13YEeH2Yy6ae0dTEZ1Ky6qtGzhAIoUJcuyHaJcHasn9fu6Az3tIl
wAsQHXugBDKVCp7WJrbnCbpsMmRcqImGJudwA2Mj1urtcHN2mSJ8kcihz0io9uglKBR1DGdtvqh4
8eIwXPXWta+1FWXa/qhXRpLiUU1sTRFJuofhpkYp02DjKnUIKbXloi/6wU7N7pFic0M7r54PbMVB
oU19kHqb9PG7SwSzl4/DMzwsrFz+mXlqrbyVQmfCUglLAwcgX1hSZzWhNZOqkhWLC4zp6i2D4YVt
SC8e7TAH+l0WJGdT3xqz8i2rUZPpWw8jR0IBOfCVAoIRSMfJ5rqWYXH12wS+SrOGOxXAj2+X9KPG
iS1Y41r5NPMHJ/LKVhUvvGb5ekLrhZV72Q0V6ffK7O06TQwNh7sRUy2IBnVKbwoMrwsSVrItfFr1
tdjoCkxzbIJHehWKe4V0w/pV/a63noN7uhzRJm3yIUrsWe3xaXVIxzTlmO+tGxu6F+StnuhN15IW
BJ5h+ejVvgbmxKVrqaNLLAwq4gd+DcdGFXdqWCVukgM5XPl0YoHXPnZvBPPfaZn3Jk/6zp3bBNkA
iB86aDobNw+L6dKNbV3aPjdW8no8V3G6HDEXlOAgpJYIJhMo14Mg2yKu76Ff+4ORBXe4KQ0FAO0Z
7ZZGIO+zh9ZpTh4fB5BgQ29ajDmiU2gxwi2KnvCy2C4WmK4Uq+xAbdwKNuF7kSuiDo20JE2BielI
DCj91zrXiajPymSH2MfR0JU6hjTzUxILdbzDaDCik6G4OQDm8dTT9+x3AvaoZ8apgYnrTDjTA3Km
1/b39nml+ZlOJrvO/376907s2r6d/uG0TBpDV8aZo3hGasm3u0X/ZUbv+xkp6Ph1IZU4A6f7RhhF
9Xe0O5Gvp42M7ceq5siuESSVgK5UIPi0Kfft4AwvBY2m6Fi8+iUh/YpCxV3ebl/XIy1DogBIIAO+
CRoxelQhDJH0EcxeZSwGaYba5KGFGfUlu90yXcgBhf4frMYylUPzLbftbrbrrAY8A+Ez6uw1qy6Y
DPsrdtpsl/3SHR59wXML8YuX0VKU+UHUFF3FI/7ZsK1cpVzyKB0isdWwLRSM9Epo3zIKuMhuLksC
AFdDc9bf03AGwO+KyI7+2ioUHOcHb+e4Yda3x1rE9jUJVjaCjKSFZD12xmT+5T3a6Zitt41KIdH7
+Ntlf813QNgl9X8AP7QJvyJUgZiFx/2jr5sCSQcO8d3dKv8S3rAgGiXkGDluEzl0YD3xzOt6DTqe
8xvtYROPMBpBa2c7awYYnwZiy+MpH+kCW31sh2CbLzyGcsBBa3WXoL6Hcq7fSxa8s8++qH7SNEe7
Z1B7PaVDKqo479daJM+Iq86eZTY7ILS/c+40rGubw5LKnvKRtzKHfcYpTglbCDMorx3D33lJmUpZ
oCWYQ0UdZyo5e3xck6baY8HlE+h6o3wwgn0AluWWIvVnq6iI46dLSWaaN1KruQQHUNwtevlLjAnA
oLldPLsrTmnWSYJmNOJJrc/E2x4K5DUlECM+48gFEComsPqByJdGtUEnn3hKy2Z/6QzSc+qCP+eV
gMBuo3gGf7jovFnvlXNVjaCA8fLkSAFH1j2IBixcV+3czqtnNcdD2QNBzQ6tn8bPithAwrbEtoCJ
3pjQvcJxJ3BjexevbcIUGf6Jlsn5pWokkZ9YmAqig45c1qyewZ5WbIyJOFdmVIx1BGctKY3AiSyc
H6LOmP+mVj8n12uHlO7hyb0wYKdIdz1kHc8mPjeP3Rll/p2QyjAc5lvsQgKv1U6dN5TjIZGUOrGQ
KXzTDCVku0qab3XkBv/MEEOrTgUYBQwLQFGsLEmZf5p3SWk2Pwm0PS8OeyZjjaF+CeANQpYoEtPm
2WFFjapNaQYNcvVYcMuYLVi6d6LxRoISzN4JQOZou6M0kKBYE9dn3X+Vhy0543/qsmg/odjs7TvD
UC7EV0SS3+JoUxhBi6cFIZ8qhxrScokRqJm4sKltTN910tsrBjmwvZ9s5ggS0q7L+6iu4IOgCc3V
RSzj3wPRbearNh4s+vFbvMM0t7aeuuPq/1ck/nNmmJrXh+TuAJuSFbbOIC+KmagJKJxS7x+p7BOX
sZSMQq8JwHUzXw27dsYJG+uSHIEIU+VkxVJNKzGUzEYlXT1Y3J+6fMuxhcN9IkInV3PcHi0SGxaC
FxqWO4mBvIm86Qf2mgEqdY3SxeIjBxtqBTGaFr5xs/CkFqR2X21cBPGBl+yB9ZZZZVMsXxtSaZlg
1BVrEPX0dv5x41OwVuVqtkpLhT/XpugDlEN4yrSalHYwHLrVRIuakIffzfKAx1/bGLkymm6TbP72
8QaRLJaWb63zMlHQtnSBa/SAXavjwei4VoXx6eaxkfTdZMT9ZamWL97+xE0ALJijW0sgB/jdMseC
B6Tz9OkHPZYeZWo8X+rVoF1pXmR7i3k4yw0zDcUwU+KakypJNbPoQ/P07alVjlUwpwj6AQBKwIvA
wcwQqSLn8lyQhV+N6bD3/jgaFUEfw5TDUu5w42dLBGqh7pdwbPEA9rgahXlOfJD6uskC/vbcQxzt
kzO8SvBxxE3zNLZkIw/U5/aArb43sO1DA932L7yPEeDp+2nZ6ooCZVW0vou3d0angzlnLQ68579f
eMhUsCWnuVHJOsUiiCCQxyMd0uhfU4C7hwkjAvCa+Ga/PAOXoXoWUDxC07W9RgWXvLhXnBfNen85
HAGqvqd84v5DfD6bCQclDArWW0urg+rtBr48Cx5RG7hzAaYzzc72SHfsIGdsNurmd9cCYOMwjBLC
TkGqe9NYXl1gGgHJoKH/jNdGSInNquPExROShQjLIsnaaz7vOFTkjdQ69im86oXMY2iJkL1jeCJg
0TnjT8oTe/V2zxwWtBiLqAE6cHB1D/Qto/21mgpk6cuzs9rVpXRYxX2jKzszNZz4d0P5uXlC5tIE
CjKNp3eaQjFNnKkS9CNSzJTGJCbWqUgQEehvYxjewFrfzk6AL8GEZ5I8BWme+l4Y2p+hVMddJoEN
XOOW0nI/yWdjI/FBNGLyrQrzAOZe1Ay3PmB1vdPGjWN3vVDpc1F6V7uQYtw6WFqqkJkrId0tqi49
71R347IYkl7OuG2tTHu9VitF7EutTNl2jFF+KA+Arb/joMWIhZVayEWAXx7fKS7AAvYTBoLxsRst
/cLeT+voFGPX8/QIWSurAQ/yMD3yXFyZgoQ6ujLEFdM5hA1qiKBvaaN7RBiSBY534QCQ34veCJQm
Ie+OtP9mZtRvrmEnuWM217pXeDp4N260zMnpsjcEyHYtR/WB37bpAEKLgsWx3LAg3SZiKkXjuCKI
ez5kJ+ZbIwW68LpACbrhD3cSIz/l+lDewegAYuRoM5T01M+2ln6XuFxE4DdC16A9GA7qMAtk7rjT
GyDecxpIQN0Mg72tV+Eekmj1K5zjAAb+k28LEnEB/h6gj/lViJgtclRfSrHDDtypCLt/0pGKPYMH
RfhYf9M/exMPrVoiOFfkNsa4gf50wBtVGfiC0I3LEubPA0QybTSyVnRzdOlRVHnch4WWfQKZ3k9y
e5oUYrvjSRRqfcXe0taHDmNecpiulfFjNJC/W49YxK4DL8dRxGQdTKdt5mmFrRL6jvm6uXSawc9u
jMaSdZEEJSGcxcvRqpZfT3+hYGhFvzaFn7K5/I6wJe0Qg7PokFtkzqOkOxg0n8g+XCpmSgiTOL34
+5JiH+0Hkzf/JTmAtnz/1jsnc1LWEH3dP1X1D827luY+C0SWhcgsdpnCmcFzQybe+sstXTxwo72v
QtXgVJfjNOY0ExIXB8GoV6KLPse3YPep4H93J+TAthhXWpce6y9YX0yuloXZ7FE+PoseoGg+h+PD
YlgYC6Wp50s39/P2jUVsZI8JM+xkeCfLI67EathpGvTBR2buqK7+mtJouey5WYk2zS9eIBvOCb3I
yrpJONrT4WoUoJGwjsHpX9fEKnMX4qeZxOGdqQT6dy9A7G6xQHP5WAJ4IQq9gOnL1mXuHeksWRJT
hKHok6idHPdzAfYJ7G1BX2lT69xooiFhpUSirPFVyly+/zO8knkzfHUUm+kClOF9shF1HFDiQ2X6
X6TtM+qqBsjsdXxjvtqLsHmUCYOaX6vsAfJAyeYkz6Ov7k6nSDDNvedq2QmzrmI+wRrMiMvEYHYm
Q7MigCixfgpZaD/Y5TgTseWZRWkDtOroMPHd+w06H83oy54MpOGBsQE/k4/YSsXx/dOJSD/k/KVM
ytQa7/x4I2FZXiURHyb3cHmJSuhOiNLaWrPd6sktZ2cIfLJNa8TtMo1TBugk9tT15bo8mltUzygJ
2UJw2fjmcPmN0p19weqBKFcRG9I2Q3dAyF/NcpsUUMhxBcwRQj7Sphfi2QJeVHEuGkUHG4BYMRr6
JNioWfkWdnqPJKs18uMNrdB4cs0Lo41qMTcgevqTsCxXljViOsxEl/ZGmFbX3gmzLXKkJ7VlGcpI
E0w4+XfkCYx4672d0Xf//9p9q2nL71QKoKKYXz4cc3y9QQ3At6AnIQdc6HWLjtUHac73iGf8uej8
CFKGgsaIXSHgeeY3BS+LhBqpHhDNGrnZTSV7dL0TT8d5cgMxJlmPz9gWaMHAMMssv6M8ch4Elfpv
6zDyHyjc/Q05KNn4+JNy/NFJ9HkmgKgUqnFT+9GRMsCYzBAkQ4qaJw6qvEcMgMkVTyuBIlp8dkKI
XKRCx6MukDhqEGc658lTOfTwhnhrk684RlydTyXJutj7H4vF2o+O0ZHd27r4G6FKAWkflMwAD1dm
c9IAYizW8IyAqwbfnJnYBdaBeA13A4YUIdVXLORcmanBeXop9bUxaq0vJSxKsNxYecZeVcqmbEj4
fReiB4CIxfUU6dI4CgkcFUtzoGXeztcxR9hK9HRi1nIRficeI+Hu+I2+oU6I3ofSJwwGulBkO14r
sSO3k5+idFup3zUP755EXz8IVnSk+tKGXxVyJkdkJ/W3icZ6mzXnUEwVooZeqcotoJJdUHeeGpid
g7lbYHkVDliItuyy0V0glyso0XcUDTJFj5KXw+D4aiUZiQYWETAV44UE94nXwSWqIvPTw3I43bb7
oSIEnhbNmDOdAmQFWF5f+XjuLWuabkEaFBMfrRMKEB0X8BItK3d67/MpElGvtw8coaHhm/cXo6kF
+XL+KoQ2SHPUPTCApqIpZg2aFTaXJyDSR1ezn0qy0yCmHa99qgJoHyofj2Xd5EObWfSJ8LNZea76
Q1M6YTr9bK4YCW8052sGYU7HsuNk5UpTeekjCE908DTf1e4Mg8cCFy062ImHxDzF2/eiHug6HeT5
+fcLBA0UfppigEs4xxjq8/pNL1Olp3QpGfLUcCIsymyoa+7yh9J0eVf7cv14lU+uoQhfE2JDDp7b
pkmrM3Uob8fzc4YokiNSH1oFzSypKBt1XSZoRj62i6cwhp6PDhPrAAoiAVrQkoS1hq9rowYnUeG0
vYMukyTjbc7ANFz4cZ0Egf5XGIz+MysZ3j+2ET8B+kh94iPyNICPUB4StZpH2PSN4Z+9u0YV9HRX
ykt3E7gP1xSOs6NRTUc5VeFaCRQk/sKPbCeuidMlfQC2NsMJJNGRIQTHO851qZv5SILvjxmse4qQ
uRRydm9NSlfumY4CmihKzObiaSgOHZhXPb07x+MScu7iv9DrveYZhx772m4dJBau8LUmK2oAwBb0
dTusFxKYSh5ZNQrPBJ89yqEugU6B89XDyrCk23pgZ/zy+UEo/wikFSMOc2qyBNvMQEPBpJM/kuwE
9mW+LTE/scz7mW/U8nwCeCnBVUyW9/sDBOU3a3yogHyMZSN6HCW2nUrIBcaUttyu80cAMfSpLn7u
AofcRVBivftJOeqlGQb7cdTSnkg5NpwjkFNBZsaNKYiaLOr9Ts0k+UP8xCaVO6kXIYEubRX5ZogL
KBqC3lo+bAsna6iZb/eIyeCAK358pU/vv0vNwdLG5dlUJjjMexeif6TjH7SDxH/J1MpIyygCkOeG
viPtfuGH2/mqhmx98oAwKzWjiqN+l0cSv5kQklFCbWGcw1DNYnDHJS/6Hrmq+Yfv+FXglY3R8stF
/g7FR14yfM+i8CwJXb3ci3fILp5IMjSl2G7SG5zo0pf8b8HmZE4l463DWfco+CuW3YClbziTSa/w
pCOmOPQvkGpo52dA9z1iEf/bzwghf3LldjPwxDM6K14y2f5nnoSmjU58cxa9ARhdRbvfG9DV/MVP
cYqwO+iaBGzSfbNld2SDa7zUD1bIN4gBMUFiQFUcKHCOuI5wDtcrSJyU04P3kCZLtl4yF4e5Ia35
N4idg5lAwGhnJz1FfRzCDV1qETOLmoFiLGdXH2LykAc6mieKp1SZ51/fDr/DLpWDBvGbyVL2xFyS
uZBn4g+DfOhlm80jRm0d3HVwaTTHnkkl98h4hEkBCirSasVgSPSSgnLwDFDcsqSEeoNybgjcaMG5
QZ/CRklTCjf6qplrdBhl2P6GtXZt7glmaRkCjYfQuCb+3HNOf7uUUL3T379JoYb6dL+N8eG8aoMh
dyvQLBgFl0sP5wD4Ay1aPOtcofHXkQXVeeXEyPjv1jO13u31ngKJbP1UTkoGHIH+/QOqy+kc5Dqz
lQ+Grdq5wATIwD//T7I8cFZmLVUjlILmrAbm4MiJbSyEVdlm4/24Sx2FPEPpg4129MM1BN0JV/E4
NbNAe1bGGQk1EV45Y4WRqUqyWzHCvRcSq6hDwrvp2K4wdSRQTxdcF/CongF0FBp9y+PMrs9xygtv
sFuQBdWXSqxsw99+pTCc6Vk6n/h4q2dZjolv8bSl5fO2luhNW9KPNfPz4PIMkPhnD/UwcAkErSsx
B/ppq5R1Av3mGfvdJstw11elEyFTQM9wUrvlfYMHvdVCYmMpN3e81F7E7lbAxE22kqceeGIryU+d
6B5R52SgQXdbf3+0PLL0dOtXm3EqnAfbd6FnItg+bWuGnFCI1QPOoHa8SCrjBefCwFUdijfBx9l1
RdH8dhLQKWxGdoxtCJVXP444D5t97XxzOgL+fZ7CrPu7pnYwZ2pNJcDFdq435I/OKb2ejHavURBg
iNgXtjLpFAW4nePlP79eqPaGhSIJkftKzM8QvIJnZU46g5v276luR6RqGqUn+EljyrUdZ5wi+Gkp
7TVwFs6UEONBD9mxWJUR+xm1bbAHzsZZ/1AERq6dXLOJbvzyZpfVdb0pK7mYd9sjSiccOItSj+iJ
z6jX6yhVvf1IETwZeuTD24uXPxP01JrWHwUI67Bgbf8kxBaEJYGMYreDU+GwQou6e3wHFTyHWMjW
j5rHPlawgVsV7A1ZQpIVg8+wcdMKRSthMutzFGhxu0zsxIUYIi5+rxeoyfR+ouljyyBnsYjiDTJe
zX/jBN1zZJsJTQFIyKi0mBvTwSaENqtopCWlQEgOknXMfNyG9Z77sCkO7OSifckiScOS3x51zHcK
t8UcFlXKq5s0AbKi0jda8tEYOORaUyYQSnI8amzsu21pLdmnvz2WKVlcVuYqVIiFEWrUizah//cZ
MThrjDvvI2EPD8rw5WfcRRVD183AFG5sUE5a+jro7mXXu6fyrXuR9FltECHhUUS402nttuRo0879
gP/hQUDAGrfFHZDl3IF44DP3Btn8321zCdL0exG+Lm54yn/1zUPZ/S2ZX3bfmMirkGl0iRLHCQuH
o0k6WBatFeIaaqsBU5xvkU6OcURKje0PlFC21InItYyOWCBq0yNB7UEOPpMumwcafhdKAyZJ9oQP
r2RX2/WFHdSexzNdSd2h58boz6+uYZxRll5oJICDx+6njbwS7+ghxZkr9BhUGYLOQ7XweZ0C91gg
e2x3yPDixDXxCLuX7BFJZw9TyGjcAlQ4dp+C1H+T+4OucCLIfzITjI47wSXyEnNbXvI49VKLaSME
BxIT5OFUEFq55+UYcFGjxfbQ7Gu3Di5zDVa25NyCsKJfyfSG6DkGfDxfcbFl3mZrvJIubhdEQzsr
9eglpPm0+F8ln0hRPTIHfwrlWPpCwUeGGsf7drNmAaNTOD5kWZqU+bsHTlEtyC8yeHeeY2COBGsL
TapHYMc6o14/aoDwfLL4V8iWadr1Nzrploygn7LztrTWniVnuOZ2VvYcL+QyfyclW/w0EswJqywS
2KxnlOZCOlTnLjFIq44GvnGGE8aP9jsltMikxH1ZG3YzipjuaDiYJimwFv4MOurTqUckxKp4b/r+
l4ra9dGiNFM3ia6wMJyS8DJPCaiD3kEnBlix/RyV/b9NJaepkaMyH0oarfGiR6Gskp4hkIPvaGek
pts6XY7A0ugm78Obl0653OyLMsO3SbRDc4eIBzRI4bD7a9r4j/1LZIE1haBxAtrmgyUdYd82WLO2
aFlrXaIlyrR23N/xZyPO4ol3jwl1OfH01YDJ2oQhLko/5o1c9qe9T/oNFkdf89N/U4vYyTWOmto0
urKyHKEeFPOEAWDKOznzgJseusMnmnT3VU58eh1XVG9P2vW1OvpQm5JtHquwJdtDPLbJ6UCOwGN0
vxD05dQGPsfwH+3tovcXqDkC4grYwS0Uq1VMEnADujpTrFyIN8vmlLlk7iG+UU7q5pmggzmuQDSX
rIu9nkYmgoxXIiY4cZWLWmWdNNH1jxrb3BOPwbuld8+Xi6kbl3AfAcrrGnyxXYavi8gfl+5A1YqN
W7YCqKuZZmGSNE0qJmVANDZgBaeOhY31Dcu9ycBW7onkV/OWu8iSzJQquCh/xO5w0pD7CElX2T1i
L5NZ7lnWL1DhjPnldwPx4qviksVIkCLkDazpge1dsJbW7hvaFExIc3yW68Uuaa6euVRpLOIPcmK1
Rk7dT+aRPj0WRftLFSbX57AHIBEL0M0rZU51wvrlv2zFo/grO90zjDxj19eE/XDkYXqlIykvvvKJ
czLsOZs/+g2hSAXyefNOH1WLoPaVccO0UaPksS5Y4OcEB+q5a8mEFVZB8oqr+/NHXOHQtFpbWwlv
QA6DEp3jLT0Ik9idT0MsbMeunK+xxEaEed/bM6275HFevr0MZvLHxL1KrW4EMQCprzPuKPNDR/Ow
RLJZAB1FPbDPZmmViK+Eri1JarlPLdz8dbOjDT+QYFf1PQVzz30exdyXfKrUUL93w+ygO0hAMzjX
pK00NZ04tVTnCB2KPjG2JS2iYPFVBhNR8yloTPjGjCn6s/xVySQm12ZxTzquILZUyrUd+e5hWLEC
YmFTQ7Vl91sdnxO15377/OaC1CJXr1ej3tLlNGHA9Pl1xxtP6v7rCZWoCHN2YtnV1xvIHIAA5ZUz
4ZTaLyS7rMAQo6Ecczd/VGkG08BScDGGhEh5O+BRDiYHNqM5RUFC2blMXBOptXXEnceM8ObtUmzz
M8h1GXNlUeFcsOZZUtpCOYgVQNUKfiZCJ6ohwIqD0dDvZvJtobGlNLFYXl3qeACxhIuwZfjUMF6p
n0nPeGwjzHydL8LNYl1YBLeGriIlgr/xLahYqr2FGw3NK1YlvU7Cc9auo/O1GI74jwA9UOwimSR2
O1olVKf2vRjOMuwMzywrz0aN+yLr58WWyYL7Oya5DQ3EdwlGv7GH0Sa+HRk2cVaRW9AzEKfZxPt6
Qqzznf6ReILMMlQDJAMMPJtalhU3aiLtSe0RrROUJdWck6EHsct4I+KtC5g0CiqBuYJ3zvRQLG8+
0CN6fk7ZS8qBsc1D8krpZ9vz4OXqX01ptgVkGvGUI4p51n2QDQZJnAyjSbkcfbVjRqpIsIuv/lKV
HXhBgWwjn4TBFovWrhMIhSQ7Hn/OgmpV34R9Z82xRjgddpwlE8GK/4Q6A4ZZDDAhtj1ce8mbBy8k
6DtEiOriHxbBz27nyLi/jo9G6x3D6YikRCH5H/OeKhkHRc7RMlla+2uR3o7Zd/TyM2Rnr12eao2D
B8YaIXXDoyF/GPLcpxM+XL1NZWOi3Fs8fQoXIiXYCP5tiLwlioFRZfYaVsRQjeZX1LKlgTBmtzHm
BLzUEFovTQqOqz+G4pj8SKiVrL+HlGu8naId4jX0f5mwxJFpu+miyPrYMk3Pvi/X11gCLbK3+v/i
4QwlSlHB8ootK1DtwelaJMeVVkmqj3JlEjgCb3mATg5k0OFtwa6zOUa43/HNDZpyL07T3pbGSRjC
IJrJMexvLoMjjL8iuj5JIYdBZcBJpJIbT7h1pVrgitfpxgpzDzuJqYtOrEnWdRgoPIBubzLiKrGu
ehPsVx+8CvL6xMOAu4pgOLwfITEnKiHVtCv6inqD744bpjQZYLPq1AObmpsoUQvOeK0v9OinYLEZ
RGAWMw1VO9Ul67IFHbRIQ1VV6ChhiP1HdpymGVamHWpQvD+hyJVEbn/kYPQOa7BrC1xKOyddWB54
fGhsBwvR8BVD7q/yTy/d5PJaCy5JqfxhzuNTgjLqBJknuLyJY1n9cjOe2JAvGTnrwKYlFvHwNxJ/
nsAl0Z2QpA6FXKPskqVFBbEnB3hAHd8BsN9e1DrWu4cM1pnXhIV+17McpSXYmrbHw+VOEO433FD4
yv12nd0c9ho84+5T4//ypQ9VGy1AvvNmXVkrTWL7x3aa7kL/rscJtkRKQzPhhoIhttfN5yr8v2Z9
l6cNs/k6e68QI2TLQYGci87RD2/12f+Eq5wGL3oUZeYObzcFHdU13/7wG8aqOJBn2/UD8hHjNVlP
3VHIAvfIZxUfFSKrJEqXBOrbUSISyWrXOOSU1VFOLizVAMFqZzp8I7DRyI4cD5DFqRc68tG7m0XJ
1tWNo4FB6Ap9mOPVGkW8/XnbjAkqPVCulz2cddcFVBHCnEHy3blndyMMdLJoy2Aycl9YwAFxReUE
g/mCMKEVmcemGXM2/HNOZle79CTcpBDw3T9rEfB5p/B7y2V4Y+tsmMmlJ3E6mlx4zJMKgcSAwO71
sPhv/cuePjomiIjCqPiVXM8BIC7164FymW8d+wcGO8RNTOaakhhZ2QxGQLDGrNpL4mPeifNcCzrA
cUlNDaf3FVyLVypzfk8XYJeGrhqIu22merLn8Qa8b2v/Jv4Nmjo/XaLZYMmXheLsdSdyUV1xa+kt
nhugtX/OC+ZY15Zxp8mgUCNW0nyjpMJZMlnYbRpQOdwRLlwSlYMjfbq/S93oEc/J8fPs0Ix1Ouv2
UhyCcu/apgWGv9Zam1Z/FtF4Wws491KKdb7SHvGZIFDu6bigBpi9ggZRGhRtSfPv0JabclPQbd2v
pzRgicH4td4n+g90adSOz0I7gIHVnsy8MIM6bGDr8O1YLjJFEZBv65xdQquusR4sR9/NfYYQZZYK
TM7mv9jxD0jIFxtQpEab0RYUsb8Ps5zOTLzm0LPPPkl2Gbrnk7EFs1V0gx8y3A5Umf8vniyFe5Ty
2/AFqrOFaELzNG64W7ULfSBw6VSs79pGKA0ZhQtCLtRygzzK+wKfZ4mrXFs0ndjr8TAWf7mp8xN8
bNs1hdsqT8NdkzGjoW3PZi4GPSVpWPB6POgdBGjDN8UIG7SqrETBgL9apgyvbEGv0HXuaQLeGnqk
S9jFSxu6KrOE2E4yiNhSEE6F4q137UhP5oBlxCPpzu1GmlCXn7id/fKKYS5TAdvCt8jmuBDxcwmN
25PZBdhV44fi75Mz2ee19sia7dajrWHfoODQ9stadxCgQ4HIR4dsEz8K5NGOtqpJ+sE89wOClgkn
x8Wyfq0R8+yjA+/Un9BKXhGRx9hL69fUKKw+ONr3QXN3uT5Ze5yxbMueZv1F0eNrUnhMZArfziEX
P5L2wW7kDu02r3fVGzETMBsAvmtIVlf9ap1JCtXtfRsYJDoEO5rVX2MtCq8ZJX/A2JbXH6Hi4ii4
e+ImapdFLNiI4lesI/c/pawWUGUhvXypCWc4fSVz73Vx3cWYidqT8ROiuAItOL9cmNa3SC98q5FR
OkdGaKH5eVxSa8Rrra35C+a/za4y0uDv1/s3//Mh+0i5sXN7j2JYV+fQ7poMyWZ6pTyXY/vRI6jS
8VZnlG6M5FL8oO5DhsRhzj2hz6WO9VW1t1Fw95G4pZtolM52TYStaC7TNAwbwTNEPRImxY7rB+bE
ZzUE43H9PO3D0ULsSsoyvflwUrFL17PhOlRujnoc8R0iSW+JrLiZpDWZ6BbsPGmOwLwoYEZHiNM/
mY9oihxFlO4oR/drPCpXVKGKweUL7HUtZMY3zaH88ZRG5LMkaCKRN5LzdWaqpKUoIpcnOTJXunUj
eDtcCiAcgICn3fslHMszlIFkd4015/y28LM9SLyOQca/9AgCOLvOB3c2kGe5F0KR8sZCT0VaOEAF
/sfmsszDyBi3K6B4OwYj77nE0r4EcVtLnETuS/kuRNzVQF3Mm+GbOPJpWDz46zVd76sOxLGDW/Di
vpXoDWLWdOUaCFsbIyKwD6LTHZXIZbKNXPDBjgJZjwhbO5RTnPqch/T841eYXOeLDa9mLFS0l3EA
2B97xKtA6v3a0xQkAriyw/51XpE4A/XN9I0NvY/kOCWK78je3AHoWWr2hwTlT2E/2tO20LzUd2YL
iHiuQrAJq0MVLkiDbidgk+Yc9QAQRaEp0UMtzY8dG72btFU3C1JJMaM5cyq6nLkAH5DfxwDF4Hqf
lYr4zrbBNa2Q1EHm6jEm5pZGRi/idQbdeZvIInQXGmhU2gHELnVWcYryzgCNpzC2h4k4eRNZ9Sft
ylix/CNNA4UecPfohimKMz2L0JfgcaSLgWmqEjBszxB2yShLyX4gbZJIWenup7cgTlIcxyoU8lNm
/0tJ1hcUed2IkHXyfBvAvnQmuc24X8PcZdHEwj7x0c303CmXnEOcFvxZZZAwXtPfy+dDOerlMIYS
GYXK4N3eJqBopJ0PakWhhPY5qpmggImqXOHBn1nV8SACygj4MYZz6sqRqLyQ3C2n/5JvS2jVw0dp
wiUgoAeQboXbObQnbExRq1HCXpq+HcqLyq1JaK8EcvOBRqvvuJ8uJtRBsrmD5MvwfHj+5qoRmSWx
tr4fRg3RTTgf0WQ5nHAqpXK5RZyD/+x05t3vzVoKellXXGhDqZJ0y02zsx8YxfddeOgRalNwkW+4
G2f1717BYos2nzvK+Y2uZKv7eZYjb+DY6qTJyR47wxbp3Fzd4t04Lr4Mq9zDOn6//T7kCfMz18WE
DkrJBQ+7vu6qz9l4DO3ElI6pQH60GdX6Lu4h/a7aAV5Qxepljw2GwpSv0PI7sRxldLD8JV8IhEmV
acikt0UFkOcwNHpDyHGB3a2d7trBldCtY2f5Y/Z9gAO+g7keqfZ+Zq9ZIGG9m6l+/SuRsxuF8MAS
lreH+yCSJD6GCJlGDgVXwI5rqw1OXHxKiikvrD/YQaHLuA6TRbeV4v3FEZr+jzrrVBREXjnVfOWm
jHB+5Qgf+espKLseLbrqcPDnvQGn6x+WrjI4DUNd/zmO8PXHa8Z22n4gYG/zrKg1d94GCAWzOkxz
PDZUP9aPBHkq722K6jCON2cVhD4kzBtw3+vTLMlr5agE9DZvavZUFLnSto962kZ6Bq82xxor5xpd
a9z3f0xGnzCCG/ghTj2RHvwreuNkAAzWv21ewLtsXFgjEO3dUVZToNoACvF4XlQzpUyyk0hzo3cG
5kzPipr/YPnhwhGuF8SrV5QU3mx395E5MR/tgrj+gnh57h65st0ZMii5SEJQTY8ctFzdwbrCoK7I
lkhfCxyPNmuEoVDABdz5NQutxNLcHahhzcGcgtKl7xQy9cQ/jhBoUm7OOjLnh4F39La15VeNjjP1
crc85X93mEzCEbPoBTg1VGGE+FCTGwSaDEF808PMqcyWGKUo00BbrO8R08oFTMCH/ZtEEdd7EDOA
sLWXBbZZ36H7kCdIzKRMLHc0uRAEPYmC/zAWOYAJsfkYaKqsLq/rPsyo2zEEfBHbA/gRX4x1j1r4
3qmu55dgEzsVe13dq8c4Dz4zkSvEIqcHCewfftY9HI0GelwHafQETC8LWX0bjhxi1nZQHW2pyB33
BFKSXcQjpRL8G5cx/UvnY7wky8ZGwoyyF2pYXoAMJc6cHyBxkWa4WZjMzXgI/hj47BO+DtUxeY3z
l1pFcLZe4sbOT7LlKH2mw/tvckHNvhXN3gefJRQKWNQ4pUq/FTpTtiR7BTsjZhIAHnJ9Fh5OO+UF
THJgEY7IuJVP2Pg0vm+nM28bzoNgqXuyG8MDcTpLi3/aP6U/s0zhmbD157CamcmfAwmY6o0QvvNh
MOpqySvPCm1prJmu14OUCXHaknZSnCVW3+xsBc8u/DCEFBcwSQQJc4oaOFN5YOErPWdVkcLQczzS
2iwdpOEopLDrBw19EKtG3FtZ9i7jrisTQd3AThPM6OHjIGtFKnLkpgSTfoGDGQB/By42wv5wyAzq
QlrO6z5XRcdY0SFy/Y8SmHcufgcD6dtcmHNJkpiS9aB4UWYLj4tbnEvYmWUvFPDBtIBMCFvbp7jz
dZr0WxFI6k10YrvZ29UczoL6hmFknl4+jI+fSmoC+zYo0ivMJYX23yuia0Ug8mcLpx4nO/dWKmrg
0BtyuRO2Bm16fymmuBatA7AldGwzwBU+Y1JYJlQ1L4P8Owa0sx3W0J9bU27zVMrKTLwNRjWy8Qez
KwHJaX2DBpHpkSgpyQ/Pg3u0pb8LyKKTicl22mBmLk8f4dKtaVpmEaX8ZEh0/+NK4+RveQQkdX44
ksdSvzmOlIDQe4J0uTBaK29vVpQTcdET5pOXOLCav1UbYHkzT/+gQz8G9O1L1m9GFIckZIdDjN2n
MSRePBBLCPDgpUODYHewajxTTfZwqDtVWGl2kAW0vIiyyvm6ogzNClgYzNIjOYqBMgG3JxyqnSkw
RGeMyhlMgaskYyO+SpkWMgy/CKHsXyTmQ7d4gpMFvLnyRtx0/lsjhNlnIYXuyYtJhQMYsyZI5ZBS
lHm7KFtB1yBTgLhT+3MBaP3eDhKgU+QknNxBDxRU/wukDbSETwAlCgKHP9CZoKpJ6S8Y+w5huAr1
Nzi6gablA4j9sWUaE5Z3bSNfbSNFBnKt0yMsF35n5SkoKLhpkeGGse0XpVUFbmd2xUL8/3J62v2I
l2EEZp7qzohfbqs6T1JJplabQ1RMLo9uHfcoYDk5uY58E2Ulj7LcefSXMmZWrqXFLs+bUCske8Nz
g4Na3l8Wrss2XOr/v4mQse3X2w0aL1mg2cOY5rqsRwro4ob4w4XK38Czbqc++JRsJpWQjZpVnDnk
/s4DkOzDtbnTG2nrfmChGHYL6gaSRNHyGrY9d9A9Oz7I8cVXtm7I8eNPfJ7lc5sKmfToV1KQ7g+5
yydi7g3y24MJJLpB6wOCzY+evTp6C+c1EGkdpTIXuoJTBWc5FWRHyH8XO0asyOGS1f3yUaW4ZLkl
zPBmn/jANtl08gZEbx70rzr/Y3Ijcu0sefG6k4w5T0AZKPqGd+K5T0X1JGvU91Ss1MdCIuuOkRu9
iVsngd8W1QvdCyk943FNnb1xl1eMy+R/tSFzPbnX7x5w5Z72E/aLIbavqSWszGfQAkBXWDrHH9l/
VJ6FG4cGMJ6EnP8Ntd1mdQt719ZdYJQBRss4gxrBKWvQ2va9GaC1aG/jMTp729uBrcXmRfnPl+sV
tcdjHcaDUa55iG+wsL0K3PcHCUJVseXptoTDkU/eIYI8c+XIiNE43JU9lQwIFkJ7WQCH+p/ihjF4
oyfa8qN4yEn4YSwDz4E0EdLJvt5aVZrnTqobibt+xniMBx07Nc+i7LL69xOV+H2Q0epGDDY9Vy7b
O8xApztI23+WBanyLCDzfxYLUakKqf/mjZXwmvqxLClrVN7Uu+7chP3iVHee1AY5Uj4oiCtchIFP
c8jxO4OugJyoHACGYEVxRGV96qoV+h+ZgcA0+M3u8rMBJVJJByUSzO6XcZp3Vi1vekJfnmq9RytN
ABt00Ld9zrieROF/lMAnXfpnp8/f8KwSGqPlaPRuapbmeyEFj38SPqhI2Vq0w0JB840YTp0AdWxu
gWx/PWscQ81OAFPyevhqYGYoRI/a5pLnMwv57sRKDUZVKTHwyyYXDLhOivYAjAZqEvnT/aSHTSJ0
AFHA21KJXLIdg+v5MFTkbTFXWh3Q6oQfoJrae6aw0IvOXEHNFZq8YeZgTd28WZr/p57ohOMk9Wxz
QWxudEJlK/r7CKApyI0jsTkr+xHAIJ4ZWbir1KGxbGrL3mh2AQzuUS+LTqAi0iVv4dYldLi7ANSn
rfk/RqLFbA7S88C7LtlnsXDOZ+UJK70c8OJfMyW/ErqXwUGO9rd1LH9H1Ao9p3j29ZpGUoqMf/Xh
lO74Vs7kA0bZpvMZDBtWEQAsb9Zt09A+lVz6KWrQdtU+fbFic/0GqIoVrkBurTa2+lH8lRW1cJfU
jODKHZvsa/aSjtBEZfIeTDdh66SpqTeraruShCJjrluHULpWIZDRhvYMQtIuWbNrMePVmzRRL/ZP
wiNxPj5S8RkAiVdzrHLI02oHtD1ykHa60GRE99lxnhgfkvc5eymV4vb8RgJZpQh2cdG+QQUA3ku0
g2zQgA1p9XS9RyDrRaqrnMnlfqOttQkpc2qnJQrv7zO4ieGw88Z8VkDzHP+SUKjPvHU1PJhN3bD8
zRvJPS3nbisK8yPF55jZKh9tOwSo9vuO7JllFfEs1aZaeG1tBCZC3tJXyTTw8mnt6/iWmyQHq2MF
ovNbJkMySMxDZzH0EBJaqEGETMoR8GYx+1PflBRDFrSUsQ8EDFnkPI3jNba5DvVTRxTDd7ZgB/qd
DVZAI7A8hSVH3RH3hwTpO1Ey/BQVCzkMGlBa5FFQWqMKfn0kjiHXDmho6IXJMHp7gDIV+00qnocY
S6MdG6Ti7vNZuL/6L2ZYE3UiPSxza5Lp23TQqY2SQsci+oQ4Tk8OERo63pMO//0PBmGt4Ew8lKqN
v4emp3cxijXZFGid4t+Q+zd6KwM9aTd/cTdyKOl2j0U5BIweBEyNNC5f14UsjphOLmtFPJfoaZGT
P/Iv23w4CdC3FwvtDs5HJQJrIFAkgoQRWnwI4PwUwHAjVPJcoMxCDwYpjPU2LOo3wXK5XmxMTYrC
pMbJrQXDanY1yzqAHuSPbtQw1ns/nfG6Pn6weQ8ABtEoP63ndhmexSB+YF+vdRol0nPzc/jkQzr5
3o4bB3ob+eaXB1exdRCjRvNloeSrY+f834afqMXUVWX+G3gIu5AivEk8Bem6TBCziiuoKAzpvRel
uy258RMsaJBQPrZ60fWfwjaEmoMW6BKEbnkE5d7VtYUgoF/CrmLHI75qe+Qtq9M2gUCDuSpgtD1d
Vr7QXx+3ww1e9LOzxm9+pX7vl4tmdaSofrQeeSrxmKoG1af4FgfL0CzFWQkZxShKvfxdoFtzIGjZ
4tQkiWC0oNsnlzIxttD8NMLX/ijKUeT+AGuuclQ5Lq0TO53i0c7/jF03Qrqk9WpQ1OROdCPsm+Ap
cLtTsDFvWh4z515j2kQbM+rRkmS9OeT928OSW0e+NGJAS2NtC4xXg7Dc/Xp4d33TXCAANtijcSeP
TnbMZGz9JBZAnyVsv1dnXY0R6J8JMfX3gjumZul1sWfVsTrxnsw7RlswY8mHReF9OcaI15DxLEoo
J1Mn+GROM9SG2VolVrAY4N9toDpuKaF3/zVMFofnSqglorfCISFOhQGKgLElxOVvVt2L7sy4KV3F
B5fCzym38yC9JOls2cQo/U8Aa78yoRf//IV1O0dSZqzsrP7r071OYm+KNvxNlQ7cx5bJY0DsDLOf
8r4t0KsOmW7JO+ZN1WvFdxnEJ1kQ/Ty8YYzGsakZtvnuxaJFY/JsfCM2Flb7DIl7XW4eIQ+uGVvs
6FMAtctr17LKsj3TUdEgtRUn48HxHrSD30Rl0FvTM36Xga1yZOwkTM6bvywTI1loG5nOzl9INQ2w
u2rsloHMSFv+W9gSiz4cPBTMUyn0ZynR+r63AQFQpQR7ClhrwWRf24YXkEdORNLocpITbAZKullT
+Ew90JyIAxIueJ1VjqrmHi/lwXeod2em3Eidjfxp+ue1DsHcx9lISel4WefgaNa/zbf7/V84kl6o
kbYrZGXrELIZiOS4UabLmPDnuLO8cMcfYq3sjdstfyumFsqTCg64kuiRzHoCt3PpRz1SRi+Cww+I
q+FWNFfT3yfXhPKZ/J8rzLb/iJhfcVsJWIXLHt7/Ov+M4owVOMiH0ppDdmWCXB7PIJ2RatEppKpS
IMnFkh3ELWidYGb3uhGZM6qt5DbYx5ZMl9yNLZ7vYdXL8GnyEwS6cFmL8E5n5u+6cHzo2X1AUW1r
WeDmqTFaFVUoz0kgljedwBTzvC4sjXiKyvtQIStid/bTueipmIXq5vLoVzW3WzWx32JOXWx1gVFR
dn/B8cVz4S8Ci4xDbvuYlvCSZ5AlSvdakCZuJXMsWB0MyDhamQKi8TRj8jVHTjJLGk0yJ/Bnj71g
C0rMWTtkQPq4eXc81za+tV2efjixCeOQ3KOhhota0d0GshSzzsGX2MT925XJeN33fHx7J/0GY6y0
ci9GrDWxEhOgBN0ElXeqZuSDDa0xSYfkPJIBnW2d+g7RS2ocNATN5rGOalQF9dWdcZrbFZRGFiRk
wc7nIWA0VF+2YEtWRL8v6i418DqNKw8wNx41oynqeotkyMU1h8MlDpV/Cil3rryy6c0SiQZy/w4J
GHgvMq0ALnmKAvpuPQPkg/pbvTL6fHzsaMl0fifvU417O7icfsszldkHpVaXIYVpfW10gnJs4op0
wiRBu2PpY2D69vKKZuXja21W93SgACvG94W0153MpjD4GaP/2IwVXW6+XMjaOO8XbbJfsSs5w3Oz
9sM+CHle/y8/SBgBWgz336+FeED9wlxltGjZU+jMENMwA/SI4KTeXxMxy9JItHNX9Hdh28H66bkB
tWAWGL4akTJL3OuZo+wlhxfmjQHqDW1GwbIHuE441GP642B6sJTZmSTws5Jqb+RjHwOdStO6fEK6
twLdebmjVNRHHnbi1cV9fRGEshuitMm94AXA7VKj3iOeO7PZQRQu2qIw2hbjc0Hj3oDpHe+AlLpl
V4DBPLokjMclRSqx7dWYMmRXJ3Sz3Tb+fFrB3Lx9DvI1H10C8Eu/kl4u/kSNDmAZgcj7lpTBEQbA
0k59rwg3M6yr3NtAjIvLCz/KRdla0FkilXb9p3v0vgDB60QPQ/X4kMbnm8J70+7R6CBq33imj60n
0f8iyasCmQhfcrxED7jupv+w058Iy7fMuEhZDK9L8HolPMCIlfBkp4mYL4WpQcoK/jnAxGxy2LrJ
ihJ86++nwIoGFN2c+H2slwljbJzTJaYlxh7VMdf1sQtMHaOV0lph6yo49B94RkbKN+vZLgir5z7L
vx8NAx5SUts2oiK2FKmQnrtzXuyGhtfXdycBdp3WUEAQIo7fDM+ew2F6sUbmN25sU1EA9FynqwAh
y2z3vUlzn2R4QkLWJBdvlln6B7nWzQuxk0QLYateQHnOhHBrxJfAvUrsmONQUUuV9RgXaqgLM4Iq
iDfiCG0qyF5FoWNDCySH6Mz9Uz0knJDyJKCQ1Tqy+moJWhjj/c5heackf1KyVDuWtcN5baWvhMpq
HBiWYKmc48ap8dfGt/gBXnLDHgVXFC6hBFiJeGEnRegWNbGl13YEJFg2CPLczxT6045TZ/7Y66Bc
9FW43Nm5h3bokMwgpDwMfLE6AumV3aV0WsOb3FwUO/cZmc8BEl+tfVy1hTSOyfbsJ19o7xVnGmef
gfKsSUJPepa5wpSIRnYTTFO4Vrz0G5C6RTBnqFIU+OCqHULX3ShoFxjGlIn14wG27IXxPFmSaW3x
il2kyGzOHw7M+nKPBQDe0ptjGaLF96/jRJXda/T9DOz8M2xdzo/ctc5h3DVtdprdzzLSW3tMkTzr
n8s9HxtWl7QXV47DbPr5WzR5beQ+di/kzPpwxcu+DWcZHxt5us2tXRVRo08IA+QUylqXylywOwPQ
U86NAIiey+wPS9nWEiSa3UqPi1bJUOpE0OTk0HTO+r8CCSJjvArMLujykgaVd3IVpGiTSsWMHeWK
a4AgRzUV5pmEI2zrQ9xXhnTUpKbya6yPZJsTj5dUC5ta0+R4lBVsyuxzJQtxCTLOdfKWqxzwnZNa
H4uzbgoKVXLKAwwkQxpc4kjJVQUh7PvCu0aF6BqnanMMl37aBdMQimbxKfmNMHHAY5KfMJ7j+5u5
s+dGMPCJjBkFa0M6LqmlbOuQiRj7c4bkB623+ZMITa57NS6AQsP1bLDHJeKdtPwKu2is0xghwCx/
PgIqaLIzkkk1r90ROIa7RKcNeJmK0D+0v4cyM83Iwb1OfXJTL9p57K6FAT0qsaXjB105n0MtCkdg
GD9mmT5aYGFUeOWHG9j0f0BXgBjP65khDTNTWa9V4GJfDlixtaShC8plccla5rsklcp1xjgDwjDe
zTss5eEx+cjQOgn1IKANw5JMJNbMeUZLw8vfMiBj6p0HQo1MP94qJN3fXmarlWIhUk+Eu4jBfyaO
3cANj5Q4vyv5YwYyTOXTjqwOokuxLNJahsOzJ2+CA0FZOqW27JnOjKDuusOZZ1UptkZqe6aJe4gS
G1YNqWRXNJUfKhmAo/2UlZovwybEoGYtf0+TUdQUaNqoUqPhVZC4rUcCVOnKplDHCseQ8XTcHi//
wDkXyXaq2AtM7udB9dSlEFtnS7VyeU9Gnkap+KO34MRkl9aODGnGNdY6AqBgF9JL34X19zm7jh28
rfNMe4ij9RzDB6+rogXxUXq5eQmvdGdpLTAjm6jaOu1vYLaPFamZcnwtNxkxt52EVD3qoFJeCwiD
PTnPFVt3QUdzPhgycguJcOTCvMSph/dDISeXkZof0SkCsJUuVUrfABRDAz0BTt9l3Thyytqb6C/8
pvNqSdmq3+8dVBnOHKLN0ByADjKjYmXdCmtx749+DYSWZZgUQMCjlZ9sjhWto/UeEJs9jWJjdpB0
6XDFeuPtqPmh8DA7zvWgyqUzzblTXoNr75XrLD905tV6iywzhdEHyMEB0cXwB7KKeKaa+Z/JRxYC
/b/KzYUcP3jTDlKQ4WH87WINp4chTedsyTLlLiws+u7mQ+drWPLXXZ3NU7gLsBuIdmm7GOeS3EIa
/OPPVrB1lX7e8tFp0Sd920SI7vzlO7UjgrLvSQBchboXztcGAjG+ngLw8cOnvB+TP4kXT7ucxhq1
0bW0FqNhG3aOcAuH/peNQ/yNajDl28pvblsu0HRReOZNJT7UFDZFO6xxsgqZkfU7zT3k0TZgKzZj
cMzkYc22o6oD+KkuySLH0yykTOR8XzgT1byr4a5Oxuynqffo2KZ23d1GCWFMFQIUtwPDaPiwUklh
bbVSJpnlx4bK8ePq/3n/fPYUMtoWi893WuGwfbb7JdEy0Kw70Q3lnSntYZUiTd95uH6IxQrFLwvi
Jz3isTqM5uOiOZ4lo2sKgAYQj39Ej9r3dAlnikYd56IKoP8mxp4p09RnGNO6hV6SN5tyiP6a5We9
aX/svthzuHNyVqlyR9yMCHqk19gM+c+EjSob92UowJdai0A9ntkHiAlnDei1dT2CVn2vQ/1vfYMM
9kyWZLqjV/BTijILaleIxxU7exsluISqSvbozTYhFBGunWLGqdqlE/KdB3fWOrg7i5Vy3x/Xkri6
hCLC+wjezdHOdK/2UrDGr1JpNWhmS7W3UIWET2W62W2Gk9qzWPMfgFhw6Cu+WnIqOlXkJ27nUcIl
8imHsgycbDjK2pQ2Z3Zfj2beOykrsKtzihawd2fkmS5RrkMSNkrYfIalykCcOJDGSMGXYh6g/D1J
1oKM0HOJfd3mAweoqjeWHdTuKJHEscZh6COcgDvnW64w1T0GMwibJ9bURd50fkj5SkND5GlrsjkI
rWaIt4kq3C4rdI6eDDFt20GUP9kP79KsSb9vlTcDXnKZ6vPSSEfDUZ+lza+72R3AstaVql5XKQXA
lo+XDyL+j5d9VNsMq6q/OYROfNWu7cjfl+gcmkCctRabIHXY9ymy3IOtNfoHpR16BsgiNYIJCCRV
v0YHNWahSJ2YWqkAMRzo4XIX+ZJnIxTRf5IV1aClYmFKVm/OUAu+5jNXDFXnry1VUxEKSdrCDnJe
Kw+GnCiHDtBTv0SZ+lAjPllQWik/UmLN4gT+d/1fpvh6fu/MpbaoD4SpUMQ9cJdpamJjJS7iCVfo
7OaDF8bhnf7jMxIavFq43Mk3aXxZjN+8O1+fCntF+vdSwZW6T3fceHaJhXbhL5xgmljo5rlDrA9/
2qpimzdS4U/EgAeoa7UkPA+zhnF4jzYcvD80j9ulU+/Ch4MZZBNygeQ/VydI6/iX3vxdBD5yzC8J
Ga6/Vt0rbE0s5Q4s0Hjrqe7TvvH1hcQP4VwNI2KEJaxy5p5i9W9faAF6N+KOEnZNcsnyn1DoKW7z
JAfuTACzXV6WStk023Tu2zI63M2ZS6YrVH/CbUcOFV6skiNX7Gjt4NqFVQ2WZ3dzjHuTfdhHAlSM
jPR5w4wKoe9m1HBXKQG2phuo1e3cLFwGYSdhLtVggPr8SfvRLAMFqHqODdAOOMpFbaXaN/eK6I3a
i+HHnt61UbY5MQWC6GWUCPeuYk0gMqgcweB22cFRZD8/pQs/h877/mvjv1IoY1HpbU58t58gwoyO
LQcSN01frnoCyfyIKLVf5rEIajLua1C2EcmdRvxUh+SipXY1oHnM+rNUL0B1UkFmSYQZOL7BxZon
rhFYvyNInjsmyrFoPNTdLC2qYoUmp8RG4WBFjJML6/FTNwkqlZfnxgmBvBoUrk1+Dic/+INORcUH
GlfgnfiA3JWgA7v66JteDU3QuzwnEwLp/4HYx9M2LAnBNmTzB5obv9lnHwojVcy/a78WpWmzfBUc
LZmdKwl8Ni+Jw4CWmWB9b/m6j/FhBHuPbjwIdfJjs6gdMz+w9tX9avBgQFq/WAb13PCAyFursmXm
EpTY7E9UJBaDwx2rkAulMC5D5NZmPNIveRQU5SFCT20tZOHhU37cxN2xIjneJKiJTf5AHdZzRUol
TTH5HHO8bH/OHLgLYa2fLztMydcl9Ra0xgA05SSyZBKlbHWLQh7rr3sVU6u4P44LtVK3r6Kjp0HS
0ExUWCYT8+AwpElbgNl7lOu/Bp2PQTO3pV+OagmlPza9/RdgxWC6xfnUPx96p6sndwF7zWnei7vp
fCK/erhf6d0KnnWZ1VAYCgQ2Hh+58srQqJQwDdrpocSu5AXXiaWYRmWBuzx9RYfVnv+k5r3nCgC6
MGu/mApkzanXxKsDYDPoLcjyRFRxl24fwAE9N6VlLqwZk6yFqXuSdzNrziJt62d7vu08fapLi4a+
iaSvW9nlrYAjQkbkYUKTVzV9zL/HpU+8qH98YRsFp1jOryPI7JduGZq0Ha2gg0hJSdIJRYYWYvlF
jdFNYyZ2ZzwjK8WnEggqAuZD6bPqUy0VHhI+5IFgTac2RLTGin0UGNIW7q5gJf0qGG5riu2pJ7oq
Mma2WIxxilM745xrt7FHJoAIs6iNuWZjqhx3efnO6KT93OEsJsRNhDGyMTTiOKfMMJNupthMJlHb
NtKFhSyy3YKdUF4Q77/jw5+TdppIOw0LKwKLe/CtAyMcsXK1TUCX+I370nwhZSx6UPiGNdBgweeI
3X/Tt0kdxCHarSGbnJBc78EBCjnzrP1vC/+VRIaO2yzQBVj2cdkOZ45absFaw0EsfDMwl0NDSNDT
pPNFnRWrWUIxTBpNt9bPjv62rpT24zhkeGiNx2Eo+5HR/CsACXwN/b4qaHbj9C1Tind11hzc9fKW
X69OXFmpipRvnRzQm37zEYopZ6Px32OQGO/XSSNl8kPk9bct4vuaQQ+AXNLLZX2LPMQ6FeiZa7g3
8nkB6TNgz2+ht/aN/WQUezBD35v9zqPc+Omv2L/xDPePEw6K3eyvamE5MDORtuWiVsn6NdmjR851
02IYysI+GXB8jHr9xw0bz4LvsaSXeOszzkmr3VixhvmkK5ny7DDmBnv4J5sA7VRfDkcYOh72cpjB
IROWQ03fzWhP/iPcrAoXlnKppGB+8cRYjaZNj3I41l/jSMtpnfvLevGixe0JNip8RnEdsgA1fxvW
MtPecFoNH9BiE7rhjF+1/wEIdP9uDDJT6LaOJKVr6hKQb3HpttnVAvNRmUbW04VpzL0drXm7YcIS
mA4laGcmet2pyp7jOQ5Q2pLL26BIaelKtohMcxPetIE6HOfH8A0ECl68ZqOBHoZtUYAf8/VmWlnz
bKZdFdMO2MI3e5POIMCUtqhsaEKji3piDnwumYAALupO4faoKp7j3uJ8MsIJ68hmfDeO3FyLJgcj
q/xFjMQ/gimgR0O196H+OO2XCXBck+dfRxB4bBKr+teN1IRL1IPtG8dp/Hpp36WkonFVx5t3l0nV
3IwdS/hQuJ3Yk5MRtvL9V6kZYA/wP8Z57LQmfE5JDuQw0MdA4vPglITrIN8ctLVcSEkaEAq/MjUQ
Lcj2/qhWBjGDQThde9hqVRrmNWvQygAfrT98VVo0dOCaqzmgMSsgxsQcUExKL2oifilBRFbWyuQ7
DYumZKkSLfAJScQoM8vcBbd19AqHU+/5Xwh+rSNd6XKe5jcay+RyH+1f9JLGQp/iJB3mTjNZ43hW
om16J9gIBbVJUz3vpd8LPVbYvDXz0vCsoLx6mKvjpamwDbWETbaQyQc+PMGr6sgz+HJmEsYF+Uo7
ApBE5MiQrD6q7r/P8Er7cL2iSXB9/u/XXz5osFemW9+jBThuIhukzuUp049rbq0MTPyRDelWvo7T
H1IutuoyJUTqjF7kZScK7udZpjm0CLXG03GPYUKGKAn1ZFks5O/EQPOsQdBCHnJOCimsqcRc6Rpx
qqodFPc/Mo7gtZDgF59Bt7hM1H2Ie1Mgow1QZm1f3PMn1Y72CuHP336tLa/qM6poWrH0Qk2wv2Bu
RcnaSaQftIN/ApoLWWcPZkUx6CeJjJdDwpdbHsRkGBPDIe8DWRpDhaKqQ/q1Kd2xsX4V+gh26UUF
SJKkdWmJqS2e1W0B3oi6ZgNudlPS3Jh718xH+jqz0fC9uppiROvI8pLkwwFsMyRwmSHIXv3tqcJc
aewDqlB2toOCtazxr8xmXwktJ9z77bnvRgfml6Q2SrgCElS16SfIA9EegarCZBptkqwowHT84Zok
FqnUstMyr6UQppXS5EZL4H+hLeL5e/JC35YggKjfZlQzll0IIwb9JhpF9BVDM2PW17Gf4PyRUqS5
oZJZUctNxZaLZrYoUB/9y8yNtVtRXFUSv3DiDDmv55CYGQ7/0EePV6/LeLBKTPW8dD9loYpjGBJj
SCGQhMcphjWcWzJHxzD4kcHinh5Y8CBlJJBDPsuuimqM/S75kXObhvr+7tCY3D9QdkLLxnO1XoKr
6MbFfXJzPkvZtuvwUOFrOsD/DwxR8zO42U1I+tphsc8a/PjcQ+BkYgopDh0AqhIAvGO/SVjFvIF5
d2LKdhO2l7TuQ1FrIEv80qeb5HRvYxTIWmuScpsVEnEgd2QOE79DWfWO+L9pb1Inbkq/kSsjoLlL
36h0SuXvdfoaEPicCBhyZfjUfqBb/70vEcKlhABOMi0K0NiqMshHjgB9gamCkrqptrrrK+4Ydaf2
NOBYMMXTkhf0iAj7LLlhCfABrQVKpo1tpsXF2Eu0V+TsTG3zLEziIADVLwvlpYgtwFIsxiOqf9K1
EWgMmDmbwIJAJHhsvuR2Oc+Ru5zjQRA7uPwDZg3qGUrl8JlufgXyIzj3dodQFDVZgAB0YfVkBmqR
kZDojqAWxnML7CrwceNIQDvaVycpVVidKKJuym7ejksokRaqm/1uKa4KaKiUbsP2qVMOaTF9hQfD
4s00akZlFFmpWQmRuht9n7oEr+ElxMVdBNDT7X8K3T87o0VkibdtpHEpPTzWKz2zmQnnHnb7wPtb
Ohdys8gjdlrcx+vDyR+fhC8ZCv1b7fYiTEdee5VtNZeyzqCeJXwRZQ9xqdgGTStuZFzMu74ruwqW
QJh8Yd9419PmzZz2DDIPZkU6efqOmezFH1qH98Ogy5Vh1JGzcU8MAqC4IaNCkaMXo9/g0Ge8GGPG
UheePS68M+a4wtZvQI++uivtgXA2lP8nAy55kWdRhaLOzbyRvo+5wFwCSi+A+9STBD2MJ89KAxUL
UTElQj/AUIhOLVbqrHAQ9fgtdvLJx5Thp2JsY0cfNw3b+K/swWKlQw9MSnVMaHipf/2M3dCgJj51
y1pZErzIO5kNgreH8Mm7GUtkurUs4OllILc0YV8xw6urV7+BwhosAxuDe/YpeWyi/EjPIki0PwUc
iRkMO8XOW+zRimhXiLDoq9XMeL0aRs35qyasIWPW4MnubTBxyfLm6gONXoiemqrnz+kwRC/+gIKK
2LwS6O+WiTGQGWBs+Wbon0fax/O7xIIT0De02ZecohInrXR7GTS0YYl4X1p5XIsgCfqeYPnG9BdC
y6T0ZNTotBhOI1UHC6eyIlXnQ12M90sGV2C4iwF5lDlnp9ybTGJK0IT+7F43hVO8L7/H+ZANmr2T
2RRbCNh3hQg/o8LHYVdYZZL4kmJLsaKyNO9bFzPUcRy1+Loc45O/aEdC+Ca3YZ4xfuTRy2hi40Zw
QykQaYnGssBZio/93qGHyRuuEW0rhnVslg9XJyGCR6GWFyKUPuaUVGcwd/i6f3UfoK0MTszEB+OK
F/4Q73Cbtc8j4c3JZeX7nUiCuNdYw5C3jEQFdFVdW9QgV8xtSI+BFBV/4LfPJC/bWr4Ti9EMfyPn
m1xmKC5Z/xmEBfd0/6Anbi4DZ8H4jivQOg2ebNXyXCUWwv0/C7CUACheJam7ne+u4ApsagjnpuJA
6MnbcAjZFGw2ldDodh7pOxfxTYDvwo9Sjdd2D+dGaWQWbBQeehsxk80k/JH97bE4qklEonRiNP2E
yy2XDn0rOZt+g8PyywxgZ4dVlRFbO8eIUloW5fQpVXrFzKB4i96jL0M7WEZo07UUGNBCPfwgmIZZ
SD+Okmb6WPTkHsGjP/ASBY+cBLY92pHt80Y+XlvhcyEFbUKw3KpJQE0e/nnzgsfYX//WW/uDfcNe
AGXvsP8b5AY/F8l53WFNBUu37kpsuTnRmYPoWVIh0gptWV8LP3i96BPodbQuFBETByMZabOX7DF3
djdWrthaQYZeqduus8eSe5QCmfuNWsfgehprdCRKXRMO27f8qeqHc/O1Jecq1VoLKNb1JHxBkqWE
uchGti/wAmEvl16utt0+0FNBZ2jwnkT8V0ZMeZ5dS5WdevYTfiVTvag8mJllvTTdJrjWaIkTtC5V
S2H32ozu0VlEUYbt2wZRMcsCpayGbSpPDj8LJCUMHHqj28wNLmdAEiybIVcSJOvQiDlNREtY3V3o
CVHZgdIE3xpOs41lR9M05T7iP/5uQou2SoPaSRj9zmRkrK3QbIGPYhNNI4Y2ZRWNfHWN3es9QFdE
ByGMrlptOCBndlWCz7BM5k4TOREZOHQxVzaFiNdp4WnAybJMxLcGftM9AD4y6ZN1zltl+Occkpv6
zORfqnFONKtp+Se16L92jnZSQjj+LpPV6LC1ft0E3Kdz7pKK3BmHxZ87s9phgmrbbUVbLUqOs2gU
iZs9YXIok4YTn2MhewBRH1Q0mCktnPNhPEpphU/Y+XCf4nezJqOMmn5au2jbC/eRobeqJEcy6xWQ
qF4a6aLpWtHbz5BmGp4LmgNuPRpOJT3PpAqVQcPy31ynSKO/Ry0Bn5ydddQT7u1yjpLalsSmH7yF
PPvEKo1U8seXipKq24wauDdFoftanvC7mBvb9qxdSr6rBaj9yaGjLk0NDpfHK9M5A2pck3GNjE2v
X3tmhr/Y8rSIU8+2JLMdx2MLWQX+WBoxm7WWb74s9qlvMokg8q0FolAWSqJJzYXDLIRD3sm856N8
M0heAAcBe3k2LCTnjDXwUUaLrgeio12lE+YNtPZoCBWywPBlt1kwwBVqsNGS5BfPqI5wJ7nMuhAR
fq//GaWd0Eoq3c6rkjZdFS+fRBTk9QIDXvveB54RdONVdUlLRLgOT9rdbQ9l08gDcgxiTfDE1Ncj
7dZ1bYhj/cioLUkFhMzEB+apCr/FqjZ18/DflFQeBZFEfUhXI/rIK7VBR54M4FvT2u+uR//BmIN5
yRcf6yPNsouFeSEKnEo4q5CvesdN0EzT4kmkGHKisIaDhcOFSJOuSv2SsSGtJbqbePn8fEy/FAo0
pG3Ewp66Ze/RhK2VfDy1ZqeO5rjGR5PNYCtvCr1MYxp02ZtiiTsngDrZpmwrt8xCQ/kuSjABwi6Y
qx9GcpHyPHgqdBA+RvSoH+nX3w9s+TA0Y2tuTTynW+RbJp1DdEV2F74y1NSewj9jW3RCMjM9CdlN
SkZABXI70sFqePigrPqBjkl5i83QiEC6/VWbBONLfY38oKbrHyJj0MpEi01QtG9/uLOxgUp/fqwI
9v1rfeQ7qvCsyoCRBE75Zcju501s5taxAnpoOfgu8sNfEqI28c8LMQPeB2xMPDl5PepGH7oSVXeR
NIUi5MNjQ9eUvWUrev85jlPwW1MPsZfr+hDO0oKkUR7qseNHqLR5M+EzeUXgS8+mAQ54vmwlVpLC
lknueX696NCKs6jqmvraJN0l5tutaiBW6q3R23YRlF3vloTiJTOfXD4LtMRoxNnCoznAKWj6Id2/
s/4uKJi+jDAhBYbnqaPZR94FI5AM/R+X3jLCd5h+n+4e2HyztM3wXysmVN4TOxSIoSHhDKhD3Jet
kIA2EBj/681Khq0dCGFmBWCy4tBlJ0TLBaYxRuh+YAtwLf/8EGuPv5TYwbFYFnlcznvl0sL7SaQx
iT1Yf9m/VbBH9fDd7oAoo80n4AJ7TOqb6oXDJzJDSuUxqyqu3Grl1+lR8fv2IvOeP9AzaTxPqqU6
aE898FvOJCWwvQCsdZdc1RiHaqDzeIsPR22+kEsp64YVdpUj2DlYLD7nkJasPAoNIOyUaZtkSNRu
lM51KCjwy3R06WhJfNmXlx/C3Qap9ZWv2r2aXpXV3yS8NrbsjMP/e1NRDaw3WhfDS9uV3HXOaK2Q
sW8E/duePvBIo967EEuv9Qe6bN+D5ranOwgx1uTqfrdaCH/2dExfi+QlWqbLJmXMSWTyzy+exm3x
gGuERsJihp4oGjrbt8cJ0JlfvAdE5BcAORiPd1K5iuFGNrUdPg3ThUuMcaSzNsgmnAcitKtnTNrU
nhwGj2fBxI+U1M32w3lIaZQsXoqGiL4sdc5TEeEAAlRNfbpV5R/DdRlsexsT4YNV5nUA/DG/o3ga
kZccnM9x4H3HOUbk4cqWni7R+il6bhQF19ttyOlbJjZQL73/ecwo3e4K1zIAu6TPqpzhUSwLQN6M
s4Mh7DQbGpEsrZ7egxBZ0YM68M9mpEwdQb4Uxe/dKw5mas7UpQayXczsXFOf41uGvIq01Nm7BGPB
YpWEykG5ZigR56McDeP8U6kb3qoS4O5ZPOi7kNUQ0dM3C9mVNgHbrsqzLZs7EIhHMF/jxHp0DREY
GyHZgcLx79PvVClVDVlwXdLEMRODpY8Xtg30QcltmAWPDbQ3j+NJgza3TNN8f+WpVz3MMVYwpJis
XnPm0aHJk48QbtXZYzzfcj0rt+g6cu2IYAULvj77QvNwOqL5JXDSXCF7pZBsWZvBkhb+vHn7Xu48
v4amWvQu/Vbh6QajoSXwL9CsYisuS2Os1Q+OX9zd7Umf5E5IgLhm+S5KIps+hc6msVCUVx1mImve
PhLm88W2ys/jQZp6HmiiQCO98xYSJm4sM0xE4e3t9t91Ty/+DJgaPj1BbXj6eYi5YUYi6XObtVkw
Lg0ES5aHRWjW4qkXH5FtHl2hL8er26U6di3M4yQZomug8Mrc+TaghzmGW+PR/crjge5josFjIiR5
UHaG7uDSZeFhp1pXBqsvUQhMbqMF8vutKQPEfQNQB6FNwLFWx6KJAghP1eorFxD6HT94qRqtPyTt
OgWbb4GZoXBwa45Uao9q6bShTiQU8CVeUds3ROV2zbPEHaDWANTHBJPaSqfW+U1YwAmhKV56nF3N
scJpptqO/fvuHfS53v8EVohu7//8tK3Y4UFMnoy8niHfgd0PUPdhg2sWXJWbKDmec77mmzfTNr8s
/gyadJtkP9H+ZUWbs5eVdO+kjymGO3LBmxxDElOV1mpgd3179rHGhVjBbUS79i0l0ZWxQkLlA8lH
XzHBSIm9I8BoU3X1tiys06EITgGDTPf6iZL8m8F59BjlNUR8hV2sJykLsvlosstdbsUNb4C4wnV5
CufGN9qirLkd8KbUTCSj2R1qprQFaRX/7ZF1ID3AqhD4PRUqW4Jpx5/LaRb3Ap8F+qKfZG0QHyTH
I9M2UaYj3GweUwgiismHaT1bTcNFhoP+YvZZQDrCXt2G63uAIGYetx+VOEqczRhfeD+G8vW71DL3
mDOWioXl/HSyQ/BqkcnbiXRyotJZg85tWDDRSbfP7kOxK2nva0n2BC1TbA58VSajR+o5wI1aNHDm
M3ZW7KqYdsP2pX7PG+dE9bph/IySkscm3REK8xdBOQVhAfWOiDRa1XPaYAALv/yh7YmCSX7xQOOq
BL2Wyyx3hES6d6Z1EN7vlPTrMcrTad47y2oc1BBKZxMcUFjHwubVnJ5oYWOXxxE1yRD3rNihgF8Y
AKV8G0v3jdts9rTCdLbfPdVsFSLnUrXp/ynO3ouemwYYAfpcj64egDqO9YJuRqUmmQvOpnAVgZ4V
ZwsU8kzL/dxJec/syif+wfj4iDMTLm7kTCthMJ/MMHlf6c2SZ+jYrJ2xJ1TFWgbOHqmSsE6YLxW2
gh5vd4kuZ4cbLKH6goEW4Ed6RrPFWYQRvqVH3ddOLuDHjZMKoYNpc/CbGpdMftJ7k8HYgacw6e7N
RSjUTrtD7zfwMfqykh+IkxYkeeR3p48H33WQNWQz/uue3GLb5j/rqJS2fHzO0fEaqvS8KxbLmqOY
3XswcHqBugX/zK1XXaOOS5qsUkvIkOdOu7kSqimmzpFErKeI/7f99IoEGyMWq/+UwJTLE1z7P77X
Q488RR8c5WE4E56Qh9CbhftxwdVbRJksTXDqXc1IoA45gGN4RaRZ+CPDUp7kZnCCUFBR2VUzwfSx
RdJwbWRsi5I8qiiibX6eTohctRVBLjFwhIrz9g1VUzMe9xLJ5Jv6s8hdXgDEj+ATxgUI2GPjj7rc
29111S3Rw4PjYVQ5s2rxBWXkq+FiNK3aHLpXWnujit4pTipXGC5myKjiEBM9KK7jTNBQN4Pfzkic
dWwJFyUdEBXfeqAMnmWgnV7hRnC0sRhHgRcrNqFIKFapQJ/2bAFSfyYkT5Uj2LqdOIbeXudZIdkr
3UdOczfeXbXIfNms39sU0HojWIG/SV3J4/kygbeHH/4w3niWtV1qYH05JuuynlQW4LBQZiCb124n
9piIyFiNiohiN7w2f/rPjOqv8/Km77aFD9k22eIp8WloKVdGOU+0TXtmZFNBtDaFwAJcm0biLnDH
aQi6MCckdqf86EssLneFKCvxHA8Cij2ocgBMPr7ZXWKPVRXHXj6XG8JMnp6SZ6igNUjk4fNkG/UX
wLK/vE87xCOtHFwJ4/VDqoG4GfhIdAKfgzk+Dl/BfAP3ZuDx/WKmbyiZv6y0cZ1Urkp+OsuP2aOB
0CqvmJKPKMK/IrAe7qBl33WZcx7vYUiu8mpulW4D9S77idKmn6pu8v5WW2Swx5z2znJSorA/epNU
pE1Bg/ZubYayFdOpvg4j70yzqkGp2cFlGvuL8+s0p6q9KvixK5n6/ZWROKteFcEisxJp6ph2q+Js
+eJqLmxFCI1CHigskg57mzXcg85vqGVu92GVpHXmiS3Na9FKGk7O5F3ffqS0j5FLiQ+W7yIq3Frh
Dqq8d1sVCw4/Uo/SgvmgfU3/fu2Th78K4ZQNyL/yb6q4Nt/RQq117UEwcJwLl6U2V0mX308EFIRW
dKPTqRddonuEMBJOKWDjGGfg2Cx27chAJKYgDg1lSnwuPSAeiElcRcX6M3PDfR5aMrJgTb9cAik1
Fu7+Akshdo2l9jd0XIfTKZLVIsTorFirM36BZcREuO3ysqfXwW3/u9lC8yY4ZWbjHoLKOIo5dkbY
JeoIR40T1aYL/Zdq0VDVdXwVfyO+fg224znKm9t7RdwUkkjIcw7JztvuEdzTJ84cCH1Ct+12AnGr
o4WWuQo7TIzHa8v/hndb9kbubc+6ivuYx/mZbqHyfj/xxzWC5avCzHHxU7KAnGY0jVIPD1rNNySd
ZuCNsGYXPJl4mRyKD73w9vQfcHOon+iMT6zeL2IN6a+aQKF6r3CCbMSgFkvHrkh1U2CF9kv4wdsY
vrM+wpCFAmziv/5rYun2UpV121uLSKK5p+LtNZP5CU5YT8s5xZyQYJ24zV+h3tXyQqjTPWebHQF/
PFhQR3W2oVbBgUmgtcAPpbi3kQ/aQSoGDlhScMUIcnbPr2fCe5P2LqDBedDgVog+O3QfYAUw2rdH
adBomEc4KxkuJ0hBGVm8aaYWKGC3TBuIhI5wC7pzpjut02aaYwLwmi2ML8EMUD2BnotSDgpOxmpx
3JQGSy6Qvkn6Ulllq2bRRizYd6BVVnR8FLkDBxk4XxLNShSQQ2whgXbk/OhrNevPs/swQ6zEqkep
Iag2TZunu4LZhxv/ctqi7i88SfN9UqFaUn8ziJd7MVz/MNZ0/zohTlu577V7Se/MNwLqEVLI5uq9
RT5ZF+z+5DNKU8545rkzLpGgfTr01MkG5zMnmRjg9KrA4S9QyhazCgtl0prKp2SPC18JI0Xa9MTI
jb0FNuKqE7eQGaVHGQl1weEJ481fW3G07kssBNBadt29nSRFbMS0wVmBidPpaD7BKL9Gavoz32nj
y20CtFxfLKeTgvkyddwwBsGpG/Lc4I2E5OzevWJDlWqUiG0z11D6ohWJwYac47wLdP+jMgwekS+O
zFx+dHu//VWqjNVQaHuwYcw85MeqQDeHkkdVY95OlLUhWIDQw5jdS9OnRVe85HKlxl6FZAvjjbrQ
dvblclAgL5cMLnq7+FGPgJQQuB1hyxGB2tYgq9edHKVxqcpTOhtj4kZk0qGil1iQijoggBTvLub8
JLDkk1wrGNIu/LQYMe4RjkMeFSad7elcPms0ZUTdLeOmejLvj7OmsvcKwktkEic/wmFF2kgHDadA
JyqrGx9J+N/NHy8a030bJ9LcJQnX1b1KfhkBquYIG2U0+ou16c7JM1Hq0tZFfIWArj46KjEL4l0o
3XKRqC4CIXdHWEro1BZ+VekAhZ+2+sqaYeBIQVsB9zqVAosEErXwMTzt5fhcbKuYt/U9f4DFQSZk
0Q1AfhwxzUNJpYQi7BjM9qzzAbEdpdjg4pHWhK8PiSEUQ8WGGjKAOSky9yGzvQvXwKs+ZXNecaCU
1cnf7unYoxdJ2kCmyuGAbhYcdFrYx/USkLwdwzgOonU2jW7FVX/D5vgwSJey3d187rzIbVuT7iKK
aTmaONBmhPAo93Jdf2nSQd2xvijuV6rvYGdbpsdy3UOFW1hKbzV8Zhgbn6GILIXFc1R+qF7CpTmq
0LgSSpL2REN1CuSPjCCIu9vda/9TqhS7fLnjIm1Sjo3lVXeRk2xs0BejcNbUG3hNgAlwOBEXFT+O
f4kBPf+YzNwPLzxxeBuVlG91pX75b4xLFps/11sb9VU0XjFCHFNeZJIAI9Twslb9MjAW5PnZv9Ul
oQMehytkenBUZeqMweOgTt1h3qL0Z5Taxj1EsI75hGal+izEXkSxOZ+C2pHWeqS7EzJ6/dKI8iK9
hCQHxHK4YMWkV5RAot907P7WCe2siJm9i6vwTF27UTabS5MzQiY489dNr0IDxbiHpgKdX23SWSkv
BJ/4nRZqBH4GGBPogFnSUmo1L8VmNAulo7tPArtMma3UKe+3y7dbldPQ2JENiQY2GWdxfVsgmyMX
bgkXvWW10ybl7VnGBaX4cb46NqB3uJIJ9OuydOos+IVRWDdOy4EtJ+d4R1RJzsmd8206iOpqjCWA
fb6WCU7XUCsvdLEa4YmJQm6YA0iVvcor+SPYWLgA3E2J1CdRpXnGk7SJ58dOCJ8G08QrajWW+7de
epQCEjBxkTjVenxXQeDL7h5S3QLBAe+1OnK5B6gfCS0PfkxB6+4aQ2jpdyBx4keKNbbvll/Y7eqy
2bKl18DVjncQ1c9T6V9Ud6aYCXouqDcZpizZRWAxLEi94J8BvdlYn+Gagt9YzaVAfPNMykoSUM48
IV8inzfs2zsXYtbizY0bLkd4osEtc6+KTPCZDRP9iUMwN/ITReik+fKll0qS8ONEr63pkAWhc/NH
aapt2LE20shHpU3fFpv3Mun2RZemeGRMe7gR/n2UKiVP/dNy2/9I8RaUU9UloxC/PLeWy6jc1w6c
M5r3/tmeWFaoXPRlwhVxZ3VB8OrXnI9KwMmt8iQYUUqWd1T0dm7GfvuXeRksU8T5Vu8u8CP3F8/o
A6aq3a7CYP78DT0IwLfuKlsggMQG9VVCAMmqEljN/2rmSSMGUQ4omSKKRzztuuBhq9k3d/LyeQq8
IpgIW8568BfnEckd8s87ITShZwvpG1ULBDNcJaA1lRSyvtJ/1WCcOsAK5R1bnyqdNvi0SZZXbi+H
sjSG+o9abMQXdRNqV0V5HLqfUedFjfwf6NvLe6fJOLPtbK6F9OUEhwEB0bJza2zN831Z2iP5jp0I
ZA3Ud8i03FyDyQZSzfK/otShnDuU2nuMrHvQ44VueNXfBPuWGSguYcrLiRxBh79zP9Iq06eHCBwE
jEFxA3Mv2DSwizrf9g33By1Icxi/mdInpfSrSvarSQEbivlWKIAKhRlUjw7tFFcUE18ibZuuMHjw
xFkWFtySKoaaOSDJtTkVdPUzxgtxS0uZ+fVG7NUSMZhWn9xQbIh0rKUXj1FSnljGXCx3yBpWzzM8
FsQuXxlO/Rabvy9+GbF5MYQmBadb3UPAYzmB+CmOiOnO56cTjMi8jKUZsHoAd6goYC5G7iT1iiK6
e//ZusCrCYjhunt4LZetab/+a32K0hAK9TLB0hgpfid7ROWpne4lVLr1y3bh9F5XdkcBYJdIPjO8
T6CBaP4vgw9kTukjrE4jFbz+kZARBK9kJFE+vNxnNNXbabx/md3E0MofSNgfVU/PVCLtQ0R9mUiV
XRSINva6sduAns/SeSJ/a9faHouUZSWtzwgjTpdopOiJtD0Nk17odF5Kc4OFMvbgRw55QwmRsP1U
8NCTqfXir5Bb1InRsYKjaiy0Ca0e1K2FgcNN2p5Ai8GxWcp3D/J5Wb6XqZPJwPZXt9qDreGluAJA
IIUUWkamdlvK4gY6GaPe9ye7z2r2np1P90LaKPJ8gEUv/NkGI0JECFwZdtOA8JqLou/3b7FD913i
xZOqWyylTzR/8SFhI/O8YrZGgo/PA6vZ3af0EKt9WagCgSl5CVJxnD+hgF8APHoEkSvXBR/Fmz1C
nhTCZ2bbcZyiE0xyXHRzyNTzy3nWdxnCf44Ki8PpXm8/1Cj7kqYp4Fryf7NotpohJjAx58X6beCg
QDKmNqadssdGVx2ImahjP/dhoTNJ8SlMAf8/B5/oGdtx9IDl2tHwZTcUJ8xQZbzFemjILcd8+qNq
jrNiN0UgEPsUWEEO2rA2HQxY5NxyKTSHfe/IRbxz6Tu+3VYY96RQxjNVJyTDO9BaNQChSZs1fSVk
bQTy9BNEuuCFRnBOehuZMeQjjiw3IfPG4GhGk3NbNq2/WQQ6xI8iS/9G/5mo+v91uKsXN815Ixw8
zjNfrHpws6lAgXiqGZmCVpUqKpVtH9wbna/rki81EsRv2TdVNKcLrXVs/r/PmP07Np5wAlFfYhrI
J0XyVlNawJGrjtkI7D9HM549b36x48+3mw1si2cbJWN4e/W2OM3B0FYLUPoLYdhPXsCNOVOUt93I
Q7+nEmQ1q6zuMCpDqrcvKrRpp+S4Y0V7BQ1oHMG6UOs2Dt8PjO/AJpfj5+WpeJmCLcwlZAxLKMA+
t/uA9PJo/alp0ByNwc9pfmh+JFf+t/rVhpHogXFQKxQP25FgO/4zPAEm3XduTAdTxWLivY+A98ii
GiCGKr1kGGAPsA1bOyM7g0C0jcGxh7b4qAFEHwCI8X5GN9vFi/uOAPDBd5gCOID7WWGNn7A7CnWw
2FYWPytA3G79i86jELHUa0bqRYJLw648vQtWv4reRcA+4hpIwSOLqGbqa3iWsCwQ6zoT7MKxmUWy
I8k4sba/QSYTfJ8vYjGEKlooNQ6jYUoCTCR7zOZedPZ5HKjw297rfh0605NF9gGl8Jnlk7kvYCrW
3nn4JtmENH2dz6Z+9R897uL83VqYY4ah43CFYwatP305s9JFOZ+Oj+yM3N1OIPEmrhFrC1EMZDAY
lpiyDCDTwdLHHve7ZIOI8ZZIzHWZb0BRHaiIsYytj+dNp2KJ6KLa26FZ+r9oBQIivEPurCeOAuyO
8fAr6OsItLh1G8gsHCTaooar/Zhv0hcimjD9xa7YVbilosR66GKGgX1n2jVI35oNTamDSsZEsgU7
a9zkhDXTX46Q/vimQMgHYdqhPyUYk56//2Z6drUmpuTQ85MfbcjgGJFRvqmfeHOR7xOuiG/LcJFs
ow4Tm8kWc1iWCnpHWi+8bGyrM3erZy007F79FF8x9rI7wWj31g4mDJBbgvSd30RbgprlifefoQgf
gJuXou131DtTw+CG1tkNCwRsaiV0x8CHWeryIM2029sfdPwGaLU3nY9igBMI93HcfadoJ/0tByja
Ih2ndLlvpxn6ozuEjtkpFPG+ByQOSTwDnjl4SPS+WjKj+wUTacDki7hWXzdjAczjK5IMFABHM0Sa
g/ntJfeDgyiVrkr88UC02/oQF2jHGqgGT8b/cQ7iL6jXMi1yWv9fbBnh1BvMMShJXTOdxQcAgjCE
NG2p0zvh7hVArlE4M52lZ+aMgZnlCJ8lSLw+rGm18jTthvfn5sEh2cC4r6IwySAp95mTePRJQyjJ
WbM+yppvoQjR1rxeQ2Ufq35uZ9tVD+pODORgKUPHMdQymukXRpwSbtIsyBUnz09jl5M9sZWlwXEB
uKWLKZyZeRzFO2zuApWjQJsq4gSY3wImrHhBVKuFJPTmWBTiIyOZmEKf2ZKLjnuqV/dmdOYNCdmq
zsOtcpdA2ZyRLBq/vFqedm1otB/VHxrbtyNNyEV33N0PWDT+c+9uIZ0jvj+Xj5uwOeSPKgFkknTg
Zek+aT/pODRocKOSu0bykxzuPY75mVQW4QJ0pKDNVky1byPpMU6sGCnEPZ7ZDiZtaVt1M/4t6jVs
+F/NBtK7VdRht3C2lGxLuLNzgKPZ6SRkQ0I2vUACFzk1oiF85LVBd7177ExYfTLZw3RxhnK6+GF4
guT+DGMTYNESs94S4yAxOUVk5iVEY/g//kyT+BZZPPGrKMGxNiDSTiU1d9rydJDCo354uMtQNGiN
ds+ovlQk826yxXFALldcVsXNK4bHWawFeidvWEZfX3IBXnFQx+AR287bumTOyjMH72s6lEpEAkEv
Vlr3Le2qU0hY53l4xVU0rCk5XPFKx6TUmyToLlk9DJFzkKJHeNUik3ZvRHS5yFlnZk+0J+arp+wo
t8+7rqCoczwxPPzTrJkjCR+vT47brud852n23aZuoNU6UoVsb060E5bKxGCue9LPw78bdM1YTj1R
LA3DndcRT26pDWiVMhoX8oByEkbJHh2xWpYJe7BbcebsTkc3co1bWmRZp+z2hZUuB/fasgj98S+d
fXEFqA3F119CbMlKAhdWXVbtynuAA0KDCBAWRW6Egs75LVR6dp+ce4b1aQw8t85TcBm3DQM6WQom
tFrhvGmmHmqwkfXWw6g9ORiCprXSK8NrsUhvnnSLW6/ZltIXlb1095Lci/UKX+7Xs0xOgO2G5ZX+
wYi+6+n1ocGBoQWq8aKpvHltT6TOa829aD9AGEhHTHhHg7FTbV0Y219BNMF50GhLvyTdljpkgl6f
wJ4vrl7FKKmh+W1EbVFNeRNeZ2NFpp14/RqWWX+X4BUxKOdlJzHBQE/VXedj6MoXNic8NuuN46eB
WWCaFIvr7kMDiH8bmBjpLbv5fV/R4y+EdMUXljC+q7hKq5O7JHCUU/I/2jT9FuHUMkVJJVmsfN02
rMoyRCTkuGeNwc3DdzzlpFUQ3QEoCxKLJ8nhZWf9XhX2t+wyhRgiXz1VeaalsujI9kzoncN6vBom
1j17uA0wbWmT4D0mzmuTnRkEnb22mwgPT1qOaWZqFQat6Ju5cL7yVvdhXD+kZWuXTELG8ExNU62z
dgxcXIduIjKmlbhAxuSx/gvDwJKcaHILBX0qJa5IXd8/3c9nsTi932WKVRNFwhYx+/2F+XJcL8qK
tVEQ3EQLNMD65vlD4NqQuWwheiVfRhrqfRPlQj9z6ed2IXR9vSXkI3TRS/TWsTy9zwkso/JOwwVy
5J+v1AuB3wqzq+8Bsh/FqLbHG6UJjkuL8iWKAzy1UbljllPML0Wb35pAYJk26dXt381ZcBRpykAP
OG9ei8mAMIADDr7v4b833e4tzOeODTwkXaF3XGU/wdLte3ItEoWWP0fWkl6/zMedh3aUNAwmi5va
U48kcVU3H2ZaUy50wm5O3vCwie6ooFGMkh5qmZODRrTX/lFmC8OfpGAM8gTL1MroB6AvbI84qqW3
dQnGPGjX/NmkAQJcfW7ZJlS7cRK2oEh35C+5qA4quVC4ptQZKiTBeOMt8CR3RxmTDplFFS2Bes2X
MoKxitGMCOT1PrAjDwwOt+9VlUmdVLohGfrYFu4alm2DoWvIPTmox2RR/FAbvXzIH18hL40ndBXK
9KdD7+rFrumNuU/E9LAQPuWt+uX8FxNQiY8eMKkF2xM9Hgj5M2fT0vvUflRor89C8uWmdhhr2iVR
BdlZPcxkZ8bZLOD1TgSJp4OMa6u1bwg4GmPM+TNYtDbWj7fCgR95PYXeNnmVnkt3pr2n3mmkPzMW
hvSz4I8+cY8a3pV9pFPwEBUyztYdb7hziCT0adbAznG2mTadsIbBMCvB6VXMt+Bs3ubELNDFl/Uk
CC/wmj7WbyWUBWhclwtyY21Bi+kYxG5HnSsd21o3nCIYdLyixG0xpgRfk5md37pgDCRSM3tHrjtj
VByunQGQE1dK1uHSEg1wXqeIAOSvoQH5RGG5SDnaXqeqONNs/mHEaWF3a3M6lzcQ++O6zT7o8Z+Q
X2bmuNwnQD1Jb1M2SIex4dkHfvkYpi4g/hqOmNhIAzIH7VqqcL0Mx0ns1VYIDkUyjWqVzkOy70Ly
iKcBP9JBPkU39hEbMhXwo7GspoppkfaI2cPjO774i+renwNbbTVl+QjhE0GMrt4KMJyEJ9ri1mId
3VrZ38w3QLO8kFInVm0jhyP/pOeyxiyBGlIOEm6bZVY99nfD3zD5U5kbaCLu69QSJ4WLa9H9UXX1
zwM/pYuw5rxvEuxD61RSZf/9A88UubdFb5I0z036b4cqcMP7OX0gELkvjux3CsU+Spfz82SQRJUT
R6k7/AZpBWl74BDicIOIuAjFUr5kHwLeCAo+97u8za87I9X759hDpT28DvHXaUS4GBwKoYWAGQs+
EWD0SkXnEarYiA00/o5jwekRfMPka58RdFB58glatj+hGtMv65xGCpvm/NI3j3BD8knrirSN+NjK
xIA7vY4lB8B3oU+6+/gyJ6JDIOF1geAeigXiN3jFy4iBCwFKBl4U4LzKJrFP43fAxdQV+tg0WErK
dKozwTrHY612Ko+mWCDZk2WGuGnmLixTgkS1AHIVb4wYNNjmH/Zny4BHyE71nS4z8+mKe1gyFPrt
eJZg0B2d6FVIy/AAtZylByG0bfu0XonxX/fIysOJtKOa9EFLVC2q4R/ADWB3xnl4myzNvFgz3xm1
e8QIUdsG6btjk6+gjS2Nzck031yqmm6+zOXqwVxDtf/NAg/P+2M0hTr2hwOtgphgYWACRmTV/JQP
Wfy++pgahLYtR6SYvUrSaXN1+q+vRQQ+a/DYEpnfNlaFN7BX3BBcweWJM+9SfyqVeuU7MQC74Gkw
SrzGNVpfouv6PiJiN6LG1ku5px/TBIgo+ZmNILjByc7tMGdtbEUPDyaCd7XKNvEGsp8P8r96yZAS
bTIitNMPDzHv9b9BHTibZvWnaffZHFSqmWvpXg8d1ePMs28uTzvXO+Q6lwU/wfNGi/3VibT4pF9M
CahklHFXmWXJxSd/XmI51InTEmdAoZN7cyXjL3/lXqMZddH36UBdNfl1abGhuK0qP/lvVfCshggt
dPHzzukSxu1lei5qKDpjgsZDPNE/V19RjSx6pkoM0WTJTeDdaWqbdhTXWXsS6qLL8Qrpn9S/RGZ2
X/5xp9Kqjnu8u1/KQ8QR9h2zs9xjASafvFznmkp9t5gmNP//n7mh11GVPRONqImZtOs5+VpDiqmf
hlghUEdL/A1CYRcLx5g2ujJo3zLhN5T6E98/xZzmBxbl3WiGNJtA1yLnPbE4izkXa7lhHm399vkA
jUI9ew0tlZIbGPMF68o0OSfyJkfrv4YkLXxwJovtq8WDoExxA58c94qOilE+xsXiFjAg1gWxJpaE
oBZ8r7AOxFbm3l7VFxyMSkhZL/Uev7LXPLUirNz6F0I8lPaeL6H6tYZ1exKbHCKHBlQvaw1Qv0kM
NcGt1sh/kH3ym8RYWJcyphirx1Wa1Hij9qWgbHhmIP8dL+HO1+1fJkgPxGP0pQ6KD5bs6FRqEsB1
z7UD0pv4494PXjUV0jrV3kHZrDkFaAvrZtQ7ot8C/vAfA0FgVY/qte1eRti/WR8BcNorXCTxn1up
payIWhlhTr+/hc/cCw5YyBJJdZek3s/R7wSKJvU28JclHR5crWoVlUdmMZ9PGBDuGRl44kTXoU1t
2oTGAdY1QrfigMBuplHG1OS0QRtgF4X6CiNz/t30KbDI3RLSfMGTp1jBsdAHNh14celWyoeZnL1C
MLrYPCfU66+hm9r4qI969k7xfYd1+sExe0mtHOnZL+tTfinthccbD5aKQIMz6c4i9tFeTrnkE3tF
AlRJE9bVTz/z/pO62NjIblGT/mFs8tNSZJRtNrUSnaNAp+fnulypWByfzspxGJxktGvFNvOZUSBv
/hDzoeArQMOzBtaVO416u6hk6FiGuyoE8qB68hQKH95n3T0ABy0Wf5++Rk7/MUhEFQ7CoCz54y7F
3ZWPI2YE/HAB5U/WbROd2bhtMVa2Hl7pg7MDUjjzvgYSyVjbIwWlKaWw3minVUA1ZDnOJEg9ZY3Q
/wQGYzwhq/pJqn7OAyVSbpfYTO0kmZLb/YfATBK9PakVxDVZK9gLBorlR4s1If33aqHz5y5XFr+/
M1e6Tq3v/XZK3m4hjCZ4nUXLxGI5fsH/P2c7Ekr4RJLTswBiBAzY/YuZfjF+UZxEXKYvLYao+0RR
NSMrfYrDDpZcHdO8mlGAE72G76BlnEj8KmU2Rc8H9qy8pGi3lXvzaGKdB2h5IWK/ayc0UvvuFdON
GsBkIdEohQ8pDgcsfECAmKUnBosxKV3upvwXbfrPciPfp7bsqaHCDglZBPLQ5jwADsPqFo3NxKE4
8Phbcj3BG26T+AYtEHoZqCtZtbiBwm55/PeCl9QHnP97UfiwlOrmeM+qadRNsCfzixHjNqPeLHcV
3NCXPGRgm3OQzMxIGnGnqgxcc14iuqcenEWQK5m8NVXKrOI88iiRyDxWgsnXmL/se6yke/9XrIIE
HyF2IXz3gaSVXeN/59czzYyvglAnsQYthi92lx6siEAjoa/IsPXKZu0FfUY3dIUvxZINGKbXsNNP
NvuJyHXEMhLL1XmQ5A7DIFU26YfqlGIL7nTVWVq035nPQhIgyOm1dF1kZIkGm6NSoJsPiZyDEfpv
lBdIResPrKlxe5sE1Ex+d/lHdntt7vKDTmCFtML/r6WOnajZkCvnmKdYWayixOpCZ+AVwCx+OQJP
Ege1muysq5QFw579Cx7ehwqlzBXkmKOSkXaW3/5fI/EFiEcmH9eZKGwQMpMo7xV3p8Lvl0L63ovG
ycl3Z+qfcLe/twSNiJzGTLmZO2W/72FB4jHa1HmdIG0mkqOgLrxoJA3Z9Jfic3S6QWJolnNVB/K2
3j9whjCKtmnW4kh9F8HxMwoN3W2+mr66Ud7ms6hz3kypvCC4NpOjKY9qZJPJgvlCuaCcVMYG5buy
i/aW2sLzn6JjriOZC2MS5+Uy9R6Crzrs3IoUmN896apSI2vXf9gv77X/ZuQ2LrQLCeLhier0DLL8
9uUBWSp6Uf05IaXykCg9QOtwGo8qlaPK2Czwy7CNXApr3ebEwof3A9URFVMZ1UGDLDJRAYOBuRym
hPrXLthdaxSv+vlanLlVGFNXVgpABfExUZxB/Ji8merWSXwjskjb265EhdAUogEH+zv0oOoWE6dS
YyHcHXM3+Xx48XbU9iX8B69kcIJvPqD34d6m/bBnlacw3XxrkqaepDQ430OuNyyzuMdJ4cGfTAVB
sZ23Ji1+lC3WT6FWlCq03Fe6yHGksRPl0Cwspe6ULY2QjE+RDQwyR8sq2kbx3TiLCVN+69pMmSwP
2Vi2ImZFthUTK9AR4SxVF7Pk/SQcIAaDF9mMszUUf682ijB6G8nmElgdO6XeKmdf2MBn6d9a2xWp
4r2W/WhphZOHnhOhoS9jc/kzNXaIoxmGbtXzj9VMVOGruSPI+8rPx34H67a8XEukhEZvruYlPOoc
J6CfWT8u70p0yvKzoYiBMw5jx1Hh/aeuQMUa/eNpdmD1BsYMdbij627kuR01RzMzulLKEat2HHTD
zbHWlJ4K3weJMMkAnDfXukrDnBRgFFHW/AOa6/Tmb81Ns1R99rOZIaEpzyxT5yMgn/mzap8D+qi1
oqcIvdWIJyKXVZu3iMFXiFsXg0bNP2xBRb9yyCqPTOPjMQ31ESGJkplMfe/ICl077qj7p23e9cP/
huJGdIoAWmb+9kaI/UDsu/qIe3AnA2EYaQN4q4sQgmk+rvlVpLpxfFBTZdLckitAUQ2uF4KcZ6wh
hbSTSrfZxn7Rb8mCG3v1Ty9DUZ+COusrrsiXTnzcNgjNTj4JgApKipqFb5IOD6rsiaxHjgcHhJJo
CEuNeb8VCLN7qLPVIAMbi+DuGN/sQ0xpRmOHahraPMMkbAlhKkQPfrsPiIxq75rYCi9X0z4+Qg1l
giU5/nupwhUWZ+Vntl3fqoOJBBme9YUWYOgZEzSJtk55cFOnC/ukRMrC5U/z8BST9T1ubFK1DLo4
RFZHu3WM9fE6h0v09MPkYiG3aU4Kr0tDm8bqd5WnPelDu07fLzJ/ULCDjcH9QA6aSePGmHLkcQmD
T1MsNQreDasGkPeT8AmOj+ES58Jzn4JusQkeS229dRQRiCv2m2CWFW72RyH9/0EAEsc/x00OvIwX
djUhBV5dxh5GHx0BeMYGuUygg/qtlIZEHtel1jcL13viySa6iiZbC9WXPRDNFa9DbFBMu/6wPIpG
nJ1jZ1OVKCtcncBq6I/4bw05l5gZTo14BgkTKhGUGju/ig1xYNHF6UbMmbtr3xTHzI5SR8lKi/00
agf8MRHNavh45BivIXz/g2C8RRwMgXbBr8VSILcI+kls9XMX7npxFZgBDdhJc+A3PVeAuNyY84jU
/rZG9lJze+mbv4k+HvIJenSHoH09RC8zZHQF5yyVFsY2MD9x5djDuTlYxTOJ4tbzJyojTMh6L75I
sTQ9paPekqFWtNDqOlFJ/EhOCc+8FE52iwP5uNXzTEBcj8OtezLCmEq+PeB5LDeHIXhGqTafmBkl
DAqj3werhc4BJSgdm3G/rE4e66o4o+c8+HFjqZG/jfiyLvG6slqHS2zdPZ8J4FT20BBqHyJvUfDy
bjhQodfcXFVm1QPQEbDMYQK7eEOLvPXDNlogJy5D2LvFXgiPtal0Er4heB8Bu7qjx3Z+MnUgCW8z
udxwTVgHno83hAyI6gpI6NAR30ntvCpATUtsftWVm8V65lJL4+Un8wbSX8UTCeORUGRJSi6cd7OL
V7WnhIQdTacniEXtF8a13iUfepusl8if0YimJGgIkDV9/TvZudPX3Lv4lzynxa4vIwpqEqXphvZj
VWTTX1DItzwRYRrPoNiAN0Ca5rQEv4kpiuWOm5tqE5MFyTKv1ufNjmp/8OEsaGg/jQZVMW/mjVm8
u31Jg/Ri7iBkQA4O+5Xgar0vBK/fdoTjUxEvkfpKW3LRXUpzg1fz4KCKY2Fu883nPMkc8y3icreC
OUAuiG9YHpROtTGTIhW2z1Jb+XnDurcW2E4n2eoMylxu5mHKhWBJ5ripVqJQcWwRnFE+4IikP0c9
a9Qg8ZYCZ75Au/TlfznhmhuLmb9Be6xkfsgHrnBmpsKyWAeHO45yljrxhlg5e1oJdFJv6l7Zl/cM
yH4x9Hy6u3E+ISZL80C9JtXRWEoBbSPQTZIdi3SCDXC0fdvIt7Rx2L/jPjJQs6kNz5zyfea2ZQh6
zlf5rEw13goen1HjHJxYQrRW98MwrQrYenj6JxE5vDR1DpMfw+YRLGpxnJC3LA4M0Q4Xn3mheVCb
cOkEnqyORPoaRlwqhdSKOhDZ5HZLZ4mFlJHEmcmnMy2vrA2DRq14K+P2Sngyu1bGNufGZhdfeDob
5Uyl7ebnl0wTJlVPFhVa67Q/Z1vz8YjnLI9Tw0t28nZuKE8fic+Hd+CrgdK/fyJKCV0Yc0M18/zU
5QExEXCpgnJ61q9W3mZ5NLk27goeo4Voj4C+2fB9n1xA3ko6b08B5ZjKxb7eKFUqBBfNzyPLNGRi
zndzZvpYZ+h/70hlJmiL2hszOKtS4J8qRnw5vn0kd33ueGeqxg/rSdBVa+86Sba7+jq2WOV+FGlQ
7596T08DbX/JNJ6Pk1iOwT3uvl0WX4zuLGiZa7zFApHQd16OGMXLiuLPW0YuMQK+ok19ejHTxP7p
psiTQUa6DLUyOYJpDTW3ZLEs8nOCJFWaTSoVMm2HDmYabwt7uvawChdIhV0b/Royu21KzBY4YYJW
ddu95T5QpVZIby3r4baexkUH3gs/xl1vGQBr9OjZ074JvN4ER6NNy5UPndTd6tpeOnGZamjIwNFf
/aEHV1so3/yr1FhvVdwJTlBu4++kAbYJM35N5h62vV5wFGuVio65vP3i3HBHGpJq4uUYDSfzcjbp
eFdBNQJoCDKr3cKCdcXpt5RNtG36Oz4LEm7xVSroI+ipyd/EL+6il2z0UDaVYLdNu4bo2P97UJYP
rrZ5KPv3vXqQw0aVrKEJcNg+ak3tOZx3vFWUKXfSyGrWzdHYG91880X4w7njkW1q0I36s9udpHif
cIqB66MQA9bl3aN02UGUZdzQ9FNKHDtsZBmxNM3LrE9HwoVT7T4/dy/8NnM6z699mC5OmqEaHRd7
ZAKfQLinsuoI3U0VqFTml5wk4TIXWq3KYcLhNxFLNo/0bMSOL+RkAvNPj7BMfAdDSAkVBrStAew+
8MqKhbsP+89T1rfYl16OevVz1TDrIqumd5f7aINsi8wuFj7RJA/Qc8dbWlxhIUlBv1tryMJhjuP7
jx4g9QbfLvjg1TP+snYkU2l2aEZuZxu00mBmHn+PTPqZaZFdpFPUl3/OY/X9yPkfwpzwcb1TWz8h
sbYy1VoGEsBZm7P9/qzZQgjhBLU7SVGlXpsW0bDDs6pA2hi3h/22iEJTPsitY7pOu/YU2U2fRNlV
Ye1b/Y03vuX+9wTPhbvJzuJXbVc2Zmwd05YvISBDjq9RHBL8ErSruyzNseSERmLEeXK1X9SO3nFC
TflUsPG5d525ilPm6qKECGNThB42Gu1t3Gh2YvlJkSA0kaUSXA+/7r/nFDaBiGtVLotxy0WGLSfm
DioytXDFpqTywE+2STPLQX+4khfedUaih15fBEWE2ArOcYcyd+d1ul/FjtH/hSR8yxBgnqkdNtVa
Z1oCR548hPuUSVtFFZXoqDETtvL+k3VrXCYMmg00hSzwJ7AdrU/doIlBvHujwRpGEO8D5JplHHC0
Z3p5QMMGZKfT1ElWE0n4aKj4erwCuu+gA++zrPU8lKLJN2rK/2peJqDFpioTmbp4lfDm/eZ8onsI
9eHAlqu/NMCyuuaMtr95ENInA2FGom5x+iMByHK3QQBnkXVJmhqccczarRX5E6n0ySi4PfbMWRCP
dug9kA4tgMevqZupqXl9RMmV+Kd4cdIhRIdF0s/OcRPt+W4X+JDY2YH/ZfSW7GkfEnxFEMqBq4Sw
nSDthFFVfnbP3AeOTPI6RZ7G7J4u/ghg64ibFs5tb+32KhOyKT6eHkOoAjcFMExi4t/QpmS3zMnb
abSqiO0nup7Ro0OKV8n75DgZUar8I3emhZqlfhxNvNSzSRwUZneT0YI4sRGE0P8JPVDgrtpwJ09Z
afPW8Fsq41FScBtkyizYYY+G0Uozld6X3PZHzUos+UDagCZ6Fpk7wzZxJbquvVImeCLr9XnJrz02
5OZXKEgj/aWeyq7oSEFLOEbunjOi1WJ0AF06yFEiCiCldU8PfmKS7BOugBIPcLjmg5ICcpg0VcV/
ButBPKhq44afejrBk5NlTHJtZLc384KHFvn4Ow15slitjCfqooTDvcWq26xMeSIzmv9W2jfOmzld
TCbKL0i0bBrSXDcQ377QnrO3RuRr5HVketKcjb3K5fXuYOz/Z6RnCBGluXDlUf1/ke6qVwhwwh6L
L86YzHPQuPrNJpjU0gyWutKmAqOfI8lw4GiTpPKldtX5wAnITV1+X18wB6KBDdGMoPbr2KVGwzWB
EfwqRmov/mEY1R1YWXGgVflDc6f2V4D1XcucrGO1UX76CwhZihLtS8ABt4pWYDOgLY/p4OyNIfdx
6A0lfI0nur3dXPsbevC/pI5cw3E8XypMzQ0e5OrKtbvFhvsL0RLCHi3aDi/cS565fNZLktbAzZlM
c2pji+89t8CSZxHk+W3azMgNEnLpxWZZf7mTnpyRw5bif3Wz/kJT3Awq2f6gq81+Lx2Hr7zEqyiI
2DIa6OiU4JKkD6+1KyRy6F/+KsQmNvBiKpKqbUYXY4LZ5UZiD4fUMy4gNwneOoyqJ1XYAvMeSqSv
2VB46rtPmWSWCiOSsFdklgib7inGUrJdBTOYniPLR85nMkCfVilCGVMrymHq5rV7OQ4SAcSHzRxT
Ic0P9wJ/gg7zGzrmPk7ky5Ve2oaFjUc4jjAyhh0yLlEBQorzK2Zzp3ops24gUy0Jg9rCVGE0/J2F
ebMqKAblAvTkrdzb67/5uVP6yE8j6r8wh2+3jajjhN+4V2dyGU5wk8o31EilucFUT9d/V48CsFfE
8v4L1C2SzCdiDxZtZAzIj2r7fmIZspZiHXtac44k9q6Vj7sq+qBoJsQvVQPjcqA5cGd0FdRdVZAH
HLKh1lgb/BVRAzq5KeR+VTKbHozjm/VgOGBm7YLgYGOjMNU8mVOwS9JtGBo0yb8jbmt4ueM2fvWB
PDxO7Q7lyM51diYcyqD6ECSNciGb/L0KEIhWJyjun8qCSc1hIWCtaAQKRjka8zglCxws9VpYOpI9
CepOq5ND7qNktBr/4Nu3GjONdVRxj+IP1JB0OaMeFMQco+vTJ3IW5+FJoJBUD2YKCTvhYltX6kyI
94PE5WZsgWsfKSr/7LGVYw6JPDAWW4SDSGCUCTQczYuY4ItRr/FIwOsF9LC4eYbpEFdVv/Rg5diL
Q5U4df1n16l7u9NHey14z71u21olGkfxfnnraXlOGfJYnxT/KVABz2hHXa+c0/fGavBeAboKo5tm
MzHm0LyL2vxrs2Z3fLny0Ds0RaCHCv/lm6cRu8x2lYFxmNN0kjUIFwJ6hyvuEKRd2zczRCzW5nJH
rOU5nF4MWclXt5KM6bIe2S6X9i1iAtENaQ0kLl6R5eaeJX3BRHncYSfmGWzUssHHa1E4NF6vzUKk
1BVsnvSbEnDC+owQxUkqwnqfVWpTiPx+g62zszOe97tS7G+YIskVemGEC79t00Bal0axYHQgMQj+
zH/g7IPyBxOy3xrnKUYBkHXjjPNLgTPmdwCtyn92WQcrN6ml1RQFJt0Msijdxt/7HqorF+a8dXIA
qsvrNo+ra+vpW4h68nShsVw+A7cWQ3YnZrUErGUjBSfkWeH3qnqMKfWmwOMrhFJwH+U/fjjcQRir
hqHznRmuUaJx5hftOYuASwbSkRGDre3lVCDPRnfXNogStubeJIOJ4hfDF7qvXol+0H1LLEWWzEIb
Mo0T7+z/DMzK11BUHgL0Kpz/OKaze4WETbvcwcS4JMCQ4J7SWneoArujnrI9ePxfGqNeW0mBPFi4
ckOGuI9m9sTkSjtbyySPm/VKA4lCapAdPFALNtVzJcCvd8PQCgeT9JCeYoaeZFoUPFrVThcSbI8+
yIVQBzWqPeJyPRa/YDckC2nqyXsItHOXwjN0w7hOOqcysmhT0Fs313xAl4NbCYQ2Tv5V8BlUeu+3
PB2akcLlnpJ/cHf6J7KOwOWXROqZfB77J1eDYoXK1xc18jEyayo713sX+2yKyZZJtYy0P/mu1NVH
vsveuyJDdaFdOoh1kCRPgej1CAAOWP8laBZJbLrlcSian+fNrB5msxjrvT7tMBHmdno//Spe9Lnp
p8AKSNSP8Nc1WH3SfrABXz41dP48oUZEX2MPSe9/8IjNAvP68tH/fdcrS2UijDKeQOxiBVBWYLlS
bA88o7CKR6/4VuWmZoO6P5lH8cBXFQ8BVNjqyoTR62MBV5DdUvnNAFU9MW012RshE7ky4Z0DPuTQ
J/Vb7x72r65CoG4JX69lIQD3XiMRuW264EfhBiXSwD7lx7iG1beY6Bln+dDYECuggr0sGgF9F1tl
IiACfPiKGONTp4rgzVdsLZy1vBYpNeeTQ6z66SOjwaxm560+WzrGr5klKu2rH3fo578/m/GBlmG+
ybZs0X4Vk7S8VOuMSAV4Nd36KVKtS/0oVmD5YtWS1/zhh5uATKSyFG6FcfRYJlrHt8lDNWc8DFKO
laa5SuIV/JQt1WDf+hDO7pJ3BJOPHcjt0ZEYbQXuhhIG0daLcqI8TqA5N37ezVD7GCLXvrBxDI9q
wfVE4/4rmkGK+UEB4KVFdsjli5Xdb1ZXF/ED7GMgeVtFviwKO4AV7EbSTwgpW09eDVa3yfqXy7W6
dQ1HHgE2EpQi9biLELEqS01PskP8Ng2TnbdU1QTan5jeI+GWpH6NjG6jVXBqTUmxUtUSDRuk08/6
vatA4JxNhHkAjFgWvOueK2rJmXVE4f0yYYzkXOnvj7H02mWVuluELoLwtqXnVs5Rz9ZzrvQ56RQX
hc2GOPmJiOd5ad/oL8lG+/OkyDpCteJAdg5/oa5GdNP9HFUsAEVi1LGnTQV8HQKt2MMidHiMffN2
00YkP04gOfWXvWOkB/rFetXeXklQHsmZPPgYlMq1QGbUrIlABE6QMUFjpHgYVBJRK6iUMRV6h5vg
4Ixhs0WtBNJoI//rgnsKYJkUgkFPPX5W1UsngZ10kByEaOUGJLKoVbAOal8xWWlK0apu3IxtbeX7
J+LkOGKVRZTOD2y/7AZlDKdCwRs/pGFz+ehYCTH6kyQU7AAcUm+PlTuIgkXn+yC4k49QLACmnudj
G1s5inyKiwcFKTMGizrwGZ5X0dmWzO3x2Ai3pm8mKpBAwo6K6vSi0lK7jnS63lJP6sKcEW3fQ/vC
6zIZnG3lDAJjOp09RY5U2HBy5h/+js4iRNhpLPuh/XKklC+KlXwyfdP+OoxsdAob989/rgWpMItH
jJHmNpM6m2gZoRATx0Q2BuGChdd0nTIwjHiBBKq3L/LKRK1N+VudutMWyBNh7HZ9ANJffJMrHdnF
+ee4RI+EXFcceOwfXFkw0W5w2VwldipndvZCAyPATx3X2y20qLlvNFvfbnGjkW5PFx7F0JfxxV//
j+eA/uXaUYczY45gJ2WpyWYhOnAEG82JyfQeMZ6V6boixb+q3z85aQVXGIBv5LCbpSkx5nnC4PyK
w5hsnbMFMCRi3rSH9RKrln0XIeGZq8Ov7TVE/Nm8Wu5RHWxfRCfbLOBfWmxsX0NAAJEwQhx00/R/
SO0M9ImILBhRW1fSLSF6xPvNZ5MByj2fXO+yBdimToQRM2Jf6QMuFbHUrzg5fLNIf0ONJ2/1TwDq
MxOMh6gV7ImUztdf2ZRxIJSc+uBRp6qviL9vRCOeo4Pvbi+LVsOUmuuq8awe2HJge3wqA+2tRPSz
Fncz1a+RAo7cmG04xrwPhe3fLfQO5wpDEQCTeKMN1PZe6k+ar+4NaOAWYpvDW7pLMIQtwWIQx6eK
zGBPwzW+xP7qyKrJZQ7uiv3ch/OV2BA2YQ0gYUYMFx6npiHoJRz7pZokJRNeKFkoOxA7LfPSRNJH
ickbZuv0sf7/ig1SIHodHPaGSKP11oiWhLzJKQXgWmIajMw59God0QE6i4TjPuGEGP3LT6nr2aNY
nz5PySXJrg2iB/RNaOc3sLKpWIx8MMk/oQsc9HdrPdlQZ33q9t4vlekB4sSZo9pPwP4z1S0Fpa6m
fbBXDEvF+FOpD5sukXObeS4oHUPCPhcN+spr4BxIR9a6E/NYAoTbie4wACh0MV3kuUgnORKpq++D
V4xstrq68Mo73vEZQGhYxxstx/beLDECr02fcgQ2FxhNEj6Q/MHw/8yEH7okJXmfirMrGN+vYTFe
iaAvsmRn0zuUjTHAJYtJmgGU/VqWOFLT1odvk3ZLJlgfGP32eOTpA90FhJMqj0bD71WlMb9jgL9U
+dMU0wGdVm9NV9soiD4rsNc1nYOJ54J69DZJHwCfPZr/7hqxWBOshy0LWnxGbxzN2P/8y9X2cP41
ot/lvXuhAOp13cf6V6mqzaHtsuYMQJ5qgEYH0mrlm9m7nLOlIA1ztxjDRozfU+KipLCovqg96bAS
BzAcsEaiDtnUGQgN4wRvs72xsm86CNMwHgVyP2x4xKTCQwf2H9z4D+0yKKdcfPp4jo2ggA7KqLr3
esE/JwwO9IXiR/RpU61ujmEynujg20f1TURGYBu2hkMorAC4+gkjrDPETI7LNfNM61lHsdEiUUKS
Q64M7kM9RynYqga/X72/aEj449R/pAxh40CjgkV7r2amLP/BI1F+XjWzUTWsspF8YacZtmo+W1ff
wLAG0BtCZPNNJiQvpCrwIAadLRXKNUCJjg8qVDGug4e3EkGcl9yp3XeLC31nHqJ9WWwW+AKWQN5I
W/L3v6n9oVhHnlvvwhKa+9LSozr0Ikp/Vrk5bMDj7vPuDxolYYzv+J7wqvfWj3v6hQtfJopGzFmm
SW33wEGc4ZEuM7e9n/TSNF6lSYK6JCUeJbkVHgGYDUWc4ydr0hLw765eSn8+cXkXZta9479CVQCa
A0gHPxbaH7W3pwrGbN9a+yCxKup/oA8yCiBiJWAPuP7wUd0Jgl8U78Acy0h0loauAfBPLXVxO9ZL
T2qXtvnCuhRmDE60hZZMEgeiLOf5zCdsSx/pDS4ethsQzW8djMbZNWQGxDJo4E7dcKohkDbnh2B+
pw7ITNAWvM122hVBNt4CsSGmUa3kYga4rtorRfR5pz2uMd+7aBRmCaIGwjVLody0EIPwysEi6vhG
S76BxGYH6lAOQOlQ8NKftL3pIz8UWfxchC8B4U9O5RVutSkRP8xArFqLKVmiWbnEhTNMeR94Kz23
3LKnuCJHfuNnTkcd9aEf+DmN2Y1yiz0h9FQbyqg944lW+fIfLWJfv4w2lcIOsVKaKg7L2xMJYOTp
nCC93rng5T8dyx4gaW8d+f66yv2R7R+auNBmnC1knBJC8Sp8HdAqD10bzDdP4l81DCMMDxVmpD4N
xoQZB9WvV5JE5ggr5Vw7j0Q16UYoM4c+rN2JgJClk5gf8Gckwmwk93ivZ4c9hmsK8msfhFp6oz/R
W0mLrFkHVpuI5PcfQ/zgm58lP7OaUdmswM6ee+v3EOt9aTgE66yvzWKIDBt3vbc1Y+CDccOkFEz7
druaoJmFMiCmfyXzpzh4Oy7wxIQ2/1jcxixh+Lv9riamX8wmAUjwi6kJicPO01qRytJisHLRJHU+
R3SHa+okShaHR0kIKczkZx/koS3jLA86sTpJh0p4d5ZQTCa1q2IIP43+oOQI6NWOarWJ8/CLPiQD
hn3lLUnqz0Lm58GPMB6c6qGnCDiOii34bIO92tKL8ZSWa/QXA0b6rzlKQQsFf1Z//cHsegrIQFHL
PCPu/SAaCxzfE/NXQDhwjLgb8h4tn+fiIy0IdZ8CXfxw8xcum+7lJTVRtjD1/CG9fIfMfjCrnSCJ
VXfMbOf0lXjNrQRVrxe5a9oMK95LAAAnkDq5xnCUp484+skO0Rbk230ET5k2acRnkD+7z+QkQMLw
2IBeP0FIs+QcxzDTqAmpLrh5i3azU9Brw6DV+gXowoDiripznrITzt1izw6wtdpcE1g9MuYaY9Gs
pL5sRbSRkBBWRl9ybNowTZRljZ/g8HJDkC+VGYmC3wo1fGzdCT8WvZ1L/XGgX1kpqVheFQaPrSor
O3MvjfpMqkHrdowXvD0Fsqi/uUZyWh+4bob0VfdtscLbeQX8Nvqt894orjjzv1RnWxEbMdTKuSef
2z+JEukJjE04eXcnD9lIQthChWrHj7vB9lJjBMtVUk5BKMmuGn4UKfyJTiaNHhbkcSf0Vv+7Nkmb
Mwggscc03s2rtaqTVa1J4tLka9mG8g0bhaJvsSCAAN6sQePBsmASEXlJoQgqsWTztl7j2yrv+Il9
Dj27G5gw+QB2fWP3Vt9M1UQ1Csg/BW0ZggJUcbv3KvEKrCQ1YD4E3fPbs4naOoWf5wzFeuuVUbo6
iE4pO7U5pv3Hd90PShr43UiWT6AijPEVqhfVgn+XaifUMEJQjLLqyz09oNk7FhbrDbH92UuR/hIn
oQgmqpHCEN9vUJn2r8O0SJA+CyXXMa95vdzIHO7UzCU9AAHAC4PWERtuxvBC+dA8vvmMHXyUW7eJ
3PeYa8BjUl7v25SJeN6LWuZ9BDbxdIHXZMnE1OyiyPvvLvBGwxEQO+3PdNWy18bql647udyTF9L6
/WsgeGGgaUIHg5rJKGg8UYXWKj27zvkXFy39OJIek/J8N2K8F1yIuBqC0qZiEovU540w7SE7iM+5
X9O6WtrRnXNE/DrOlSJAnz6aF9Uji8+28n9PVOYDuS3ql5D2s269JORTiF201f82xzNTJ8JaAkOc
pCzJilbGYeNzwdwnBSiVwLfZ3JVQwZu2nr0+spQU4it91znLSFm9LDzmaQo13PDXbH+tfjuY9wK6
CthiigCtJ13rx2MGGWvxNki8YXQXF7xUE79+DRt4+t+Y9vlxi+P8uxutrL2pD311lcJ8bl3RR3nJ
EC9iFP29w0X7JFGUGV/8b1oBgFDjn+3ajMsNhwpmKFEo6VxaDlI8WmATHFByyd5gweCXcwXqIxc2
kgg5RaUh/MIn5boSgKtikdmvQxjENQRTXq7rzh3ROhP8wn8gp8wu2EHsIJZ3McO3VD056bl6GCEH
5MeRnrMmNVMXlnMJJIHxoyIyhBqVi8ge/SQCupZDSqu6xt3k7JJIxzHTuZXoyECOf1SuI01X69Ye
j++eqK878UcTitiS917WkKiBL/Sn46A6Qm9gfsLfrQ4gggAU/Fll9VWxDvMpLnSxjiKcgExagdMW
3eGrjasOyGt6LNioBwEupppsLJhht9ElxHsRXRkG4OVQriaYskT13jIhhn2SyeHMVZPqzJlvy/u/
CTJArzBfVTuFds2UeP/KJeYkjUQDTacLCllBbvFwTYWPcWFqVbNZAah/thnnE61XIIEbPZRR0JYI
3P+gEr4ZTFsrQB41GnvAGMKkNccaVDS/RCIC4Yu9ZodBO/E8qInhDogTT3nVmD/8eSeYENBthxj9
O9R3SmG9kmcDraZ8USy2bZkcQEd2/Z24fwLHXx1CeN02ZlcygEFggwJNHsRdEB/EO3iRkmRMwKDI
t8f+ry8LuxzdQBaWABZ46TeXoXcWsR0V+rxH2a8G4XBhgaz9uNQyquLXdKRd3wcHt5SzoYwZ+RmL
bWBdQln+OVUbWFh6eyaQ68TzjgfySC6a8mjokN31L+HeOLE1NhwdSdKGm/GCzKSEqe6Zwwo8Tc/l
qFshojorMYjEGK8QpX5BXR/o5HfhUbe3l2nxJ4Ju98ftvh+1XGLPATOR4UqC8KqETT0eYCp9mISV
7HNtIQvszqSKrK3M7EpScT6jpb8eI6h8/iJdKCvTOibgAghmEWXrJHVnAXwpiSqQu6QXMEYWFEOG
JaQ4KcjGN1NqGdlTHAcFV8zu8ZQF/YvNN6b+N2KxauwZjAA8JnEd2Pk0M6/6uCZkWsn/qi3P0bZf
09+QhMo9md8VPu2wI5ftOGZJDRpsePlDeiuXkM1vfyxrzEuaoaY5ZoHPBIDIpV4DPEIQdT+cM88C
uWRSqoUzM2cs+fQZYcQk9XjR6RAsX0QdvgWlmIcU85WW6QWw/5RwSpXJLjQ8GoYUjGlqoNmDjgsw
GSO4npF8WGhweq9di2dnF1PXiaoFJJRGE8oizEXvacCSUegdjwEj+5qgZPinfp1GpvHo6z4/08tI
CWsP18tEtdY4BqU9wsO2JAVhNV7ifriXJK9p4Stbhv1t9nGDjsH0GDt+edwCJ+GtCeibLBc98Iic
xDdEw+pdcJTFVnpDQcGe6JHv5r/5pCojGibi961VXz5ACvMC0IZ7AJBgtQODDBRF/GNa8/9QclEv
UUmxelAQhOrEk0gDT5a/JDeqTNoWqXI8qo6afIUWxlIt1IQHMyZV1smPBd0skfsYD2alskozZ2Op
8S/SH1MUFHC9s9MceHFX5uRsRTaErfiV/gArCC/FiFcrMZaAKUGz8USo4WWrvEKKo3VXBO7IqgPy
052EeHT8ameSYzTLyFMUR9og2iBa/PXG5dp8x03wxCyKeVMkr+Dn/8PPetkp5erToimulje405VE
j/lEGv9nYKoxxChzDfohTXTSrLS0LH/eSQkOVw6l3rjzqHDPB2Yz6Iz+3sp1wcCKuNtei0ggEYv0
JgLWHJTkxXdWt6lsESRUGV75z4L55X6zq7UsCyT4UFU+B20Uk1q4lhOe5Xlaf/mJ3pcKowA6Bi/L
b6CE9vCyrovJvMkxYj0RMx4VAuAAaNfkPnaHiXyTXbGQiDHrjTZVaoLO6FpRO709Xqj1uB+VQO6y
vMlVynE30RCQitsav8lMejfZlzn9L8GDod5ubPvV8Ovt8nmZ7lMzjICiybrFxtdPvbvnia+8gsED
tBZqcEJPLU5zoZMeHpR8H+7gjpvwm6ZcK+yfpHdhQZxAEWxL+2zkNjmNQG1VLn3XgDnCuGfGATmD
bTMztRoOPGjOH0crZk0chY6Mx/vIngMUvwsQd2ojLUtBh11LDx+Flm7xIgByKCKuQD6BL0F1zP3L
g8FDgZp4v+dsI6rZ5ALajz/gUOmM0bw8XDTy2S1URry4RcHVzWPrk+hqBApyzWN1JrELZIXrS3i3
9rhs1gkI66cXzA4lEYx7owLScxlKhzdTWXg2Vw1hdUFOSFAwnY2JNZWuEFWlzR6HaCbjUKl7aOrd
l2ZXJ6jX5vKT73+hkuO8z7t33XA1gFb4QODr4mF82qcRwlzG2lb+9R090g/6Tp5ZSn0GFRSUPiVb
jFeKLweA8qXj1Q/nczgusbZ7VIbtu82RAbA2Irj/G6N5Ekx3+/u7v+MOULVa58hdmIMxI7x7n0S5
BiCq1YkmUaKAp8TubwjODvu56GyrsWAsfV5zejGZeKs94Qq+9T6fnGPv8MDKxhvwVW4J9rLK0U/i
l2b+ESpgqTIW8BJR1UI8xG3VNG5HGmXoLnBELkxe5EGXUzxZnJRM5/mL55diCAfM1thoomSDu6sl
OeuTrubpDVLunGPA0AkW2HvDWQmsUQiy5ch4C/xzxjspZXYErCYQaCuKGoFdT9V6bIqu+GVLbu05
CRtQbBJizeuCGXbSXEx/eixSjRkBRII74NkOSQD6R6gF+qu5wqRrcJvaZfglP9WrRkEw9HNZsVCI
L5PKxfh+dE+NyasWXQSGdSEAcZ/td1ZT9msjpJsoMNn++m/kofkK7WO+7gIcDlcb1o2xKHClswfh
55tQTdv/f6uJigsnXYY/78lz/zPWYOo5GssQ4yL2bk58WMDCZtt8IBA1htG0vyWnOauHviKbc4kh
qUskdSKm2qiRsJxuOSR/joCTdSEJcaP6TAnDP6LQB3savFJ45nZjW/aCy+jmOdi8nE3DRvJh7Y0A
6GAe8WvUOg3QoRCGmK1hWCrN1C1NeLbs6HbRn3fG+zqeGc5AwBN9bCXKzcWXfc5DRmRHMIbW2r95
ruYeok1W2195GjmX4mqGpov8jExRQzdO1N5cKxzeOYBnAgWtqEKlYY8urchp//bAe+0+x23k7Hth
KVLjFesJjteg4O296E8nmUcZLpW0hPeFmYrqGxJTmnfQxyHfmpnsMVw3W9/uHBRIc5IhWEkNho82
CAcuPkHMWh84qeX8BtEnOV4NzbGrc7R/PpLs7r9Ms+MNkiWNx+0niBf+VVOoGHbs4CjiATcst80M
AahufjXVcwRNXEcVjxa+Vi5Tp4uT9dYRFT87iYVVn78iuSxTnj/f0Yeg4Thw597nxAq4moPX2uSb
CIj0M4bAHH0F9qOEJ9+JgYu+0m8OFTkn7bv90CBkb4yVHSDodEypySHByj50PUPAofzwAtA4yesk
PKbQ+J/KhFWbjuFG7N5NExjWaLnzoErfyM7b2/8Im/ofPz6dyjatdLAoC5QFJzUvkq0OjeBjciDL
j6VmBO8rX69V7YWN2e6gj7zU7Y71hJbwGk1QanZQt4TBsPHqL1LnKMw6mfdr5IlpdL/yfjQYDpiI
pDxJlRlfs+ld9grX2MoV/l5g9eF56nMJ2NI5FraK2jZil8VhNz8j4D/hslgkhXlZAtHF/qhxylRO
PGy5CgtJ1QqRoeB+r0Zzc7TDVR0TZ9aO2Hm63vO9mJzEIMnUcAgL42yhRc7cewnkl+UeNeqdNIL8
IylzhRBLHbLOzj6DQ+O9ccTxT+FoJGU5nSoF8dhWb8wqZzndIfgSqbVf8nWHRgRzzJauv4l5QIbX
85BK5p2u4NYa793Rs7xJQWUXqnJA/JSxDG3PW5lU0xa4N4R07FHskWI0fjzeoEzD0CLG/RW643Tx
fLfIdAdr+7664GUQzdkm+zjL4Xce0ZbLuSwRFjBZFkHwuzGq3GdyuM7pwuFi4JfJPxNH1gDSKWX6
BZcdR2Qz7BnWfF4eNUerRio4U9rbMpNbM/FEHYJnsnfl8qw/SPZf0CbcInVVT8ui3UTkMfSkH0Va
AHDSKnMPSgIO7+KDD2BRlkiYGQj73LAdmw/vWA9obHIssbYfsb1mZdu2aE0f7GFo7svqo63uk8ZC
NquQBh5gkfuq5VrmmPX0fp+vhVjFNj/a7kVJDqzY87R0lmw42UtlXXsqAwmI6Gf1UDqsLVFnI/Fd
JZglvMjXCKaUEOAAIMYxH6RSR5o+XvGeLildbM9j1qCxFj6BU0q/wSqxbEFGdDD4DzdXSTFk71DE
s4DkZ2Erz0G8RmA+Q2zljcG70UojVzqTzFlIyDYJDoHn7heMccO6D93LwtO9rXWkktlO7Qoj1100
gaFVFGJTUW9G4ImhAamb+JAINU0UVlWlsg7WIgbAW160QtRAmCSYR/WA+Ui8qQx+Gd5IHlea1BGw
SVx1R8VUfnOQz7ST2cXXWCJXU/u4xUUKkLoTMbjn6ASv4wcNdGRafNmDLcuXMuvlczIAPDDYGEj3
pkzZXXzW114vTWivF4AmBFy9G44SKiMalCsF8Yl/ihrJwcVfH6wr1QG96LGiayJUgvA1hgha5mT8
wT7PZfM/iy5vlg1ccHDnfORnXEv6v2+Vu+0+X5mMMD1qqP03yzECnnijtiSq486HZlh0crIzA3aF
2JOK9oUPtqW1MncsWNY6kAzVEi/uP7pfcrra+MV/5XZNLNdYohfEnffj1zjJcH+VzUusIdxaf4Qo
VA/VOKsH/yIQLv92xCE2GKUnQR6paMVVrEyD+Z3S73QxsEed/uOEklVeLHi6bjxa54x1Xo7g74Ps
4/yYniVO8fmkLZpz5acZMglfZM7GVhBN3sQ2vf3Gs9ShypgtK2Ln/tIuti54NTrVyAXocpg8JFa/
UUUvAVldlhLaXs2YAsojJ84QhCryWxMUe5tk9NMtN8+e8SFgDOYl7kbqrOCyXICEWnM4YWYuukWU
tBfH+UBlNqbp/AjYf3C09RSj8J72naLeMMhF9Wl8KXgV52jV9PHSv3TC/Mcqr/49brpokAwTp2KU
icDO8Xb6QEwXr5YoPVr5pecACNNr/EB2T+wB4vbRg3ywOQulieEStjd+YV+j7Lx59d0nPbIctuPQ
QBkGqIhTMF+C19i+RvIbFB1OQ7IveWT9YW4+wJ9oTOi9vZspSxhNEnsLx54pKrvXZiGQLl5MJg85
gmC1wqEufDesMLaLtQQDHZhiuqww3b2o6gXmv3/Y5yDUSqKDpWkykN62IN6ggfREi9RPXXyAhXUO
I+nP1n3GMSoRH3WkozIVl2P1jsc18LQxaQxSxmWHFWv3tbIWlGcXX+wMPzonIBUtBdywnbn2yCxh
nZqcmmHvXggRiy/38GWt0IiOsCrRCSVKyRLdHcedkZeikIQdLPCCf6A3BEzreBfG6cR5Ir18+V25
4puNi4U4V1vfzyPlTpZFlswm8C/tHzCd24G97ddHylr8WN68F5BicMaOv5jjKOm6H1ZPhmnXwz0X
KjQPESOkBGEoD9tuJtqaJc9l4M1oqzuTPwUE5l8tdC8wsAhMbUIHipOadsM1QXzHqsXf6p6lskvB
hSSzllGe5rWA9lfEmVYyPF1RlvEsxOR2udPMnkEyUDrcGuCycVw4Ed7DdSVkMa4RDxeFhVeOa84G
waQaCiw+FFKXARQLqQi2STxhm1LcmtL0Sj3Pl8X02Vn0G1RCiqOL7Ikjm1EGCgM6cNkQE4uSJCo7
IaV6SOGt0wUEHBXGmf5h1tw/gnEeJ4yexpQj8SYAh/2ZqQER4LSf+tssBvFJH2FE057MvrXKWxNr
t8npjyvDEkiF1BYozkZrEXwDQyeJg3/txcAm4jZgbylim7KlKis2BVNJYacBj+KXYMHGmsDh4zg9
ZX5cx44558nAdiWNZsOawVJt647h0tJfQfRCGIXYF79MWEuiU7kL/40cS2mH82+148e5DWhQDdRh
iwxKJG9wTJfDbwzxRqBa6Khlm59rO/xFHhO6XEQ8uJ7u003Y9Nxr0SMSIBbElDUGRyDyJ1Dhzocw
+v0rcf1eVAFincrFFOyZdaVSY/+3uTGQDqyszPendHu4Tz4xXHCOg1AZ/pJP/4xlXZ8Zd31cpBG8
b9tjm9WJfzwCmxjHbjMxxTZ8jT1si8qequc+GZqCkf1w9w8iRDVN1kEUnw0CgPJBO7UN3athlTC1
MqxTK4MwcaySAIC3Id5bRnwTe16tsx4PwtujPBv9UQ/09T6nvvMmupqKk8Ai+dwwHPqI6Qvgt0mJ
Izk1DYZeAzgPVipfroSginjeaosvhHcPJSbh6S7hBMtmt5l5L+mQIZ7ZWV5HV3TTQjAdoiG9Audu
yRYa41gjfeHq1lOMaPnkaUl0JpLcf2o0TDTGU2qtJOnC66PmTm0dk8D8SD+7vIaVgY0KQAhyRrCV
KR5gbv5uG8gLso1lg74NjFlpOjzcjuPPhIQyhI/g95N1XZglKH8tPHLcqd92fimtLSjUyBoRORRQ
h3/5J+kNVJSoRkCcLw7tr1eakCs/UZpQxx8B0KGOh+yl6vkmchlPOMF0NudZqQiN8/lyVyci6TQS
yjJ1Mu9RobG0njS8D6ELPEboc8YskzteFksQat7qC5Eg1GutGp+7QMX8yY/2Cnb4LEupOEI/43vH
9ZBfBov6RSUTrvbrzBSqVAoNfeXZ/PIBbuynVkKzHwtjMEFxAiB4NJAURjyTBqf7zi/Kr+LeXcFS
UnK2KmPjyTUEcj8SPhiGC7KHtszDzj8Il1RhmIUZfuYMNM+jqgxLQcgR04nOcFaFNCgyd6c47MG1
DW4A+62kLoDDd/lh/QSmG6dywNlxGJ5bZjgMieXtGGpdj8rXSggGe6EpGifKcT847MQyISx5Wamp
D915kGyaSGcjS5FrKidfPA1xv52dO9rN2zAycMOJW+nCRFyTZ+VanWiINM0kE755NyVMVlnHYnYi
b0VYTZd5eUjtKYplTox+eOS812K9xWrsWYrUavDc6RhRpqtUudk4gTaPjxB2R9KkZC9JN6nWnM6E
skJj1TV182lxG28NgXhz6yImTyy4UOe7RFlOyx6lMVhkt98CvHtTF8QFGN74z0J2ffgk/5Na990t
IcIFD+bIPs06zBtFzseAnkbRO0VR01bIhGQ+f3lxzo0DcKe0N2Srq6KQGQP+5k5al6K8SoE7dihy
9nuwtM1xJfChwVQ2GasrB6a0DmvRd8PABHU0swrEMf9vQZ8oJ6unwpingkipCd24s/UQj0ok8r80
TwIE8IA2uIlsIkcAsEtM4raMi333OR0KplKO8kZoQlr2CWiSdMZA00jp1aReHqiWVEgCep71C8lw
vpz8I6aIZ8Ugpj9z1Ww/sbV/biWnXTQpB8fVPiL85QzAWOdHFomj0PJel+T845k56iutIAaDgu8p
GTxumPTFCxtqXab3FUjr7tdtubEKvsFkMBpRQNOxdvvDFCCglwCRZLOobxfgxmn5NIOXkQ9XDx1Q
/KLkcn37+iLXWaoexQyqF9hVkSm+qnS9quQCm1o1ptjjp3e0EclCkrJPtQPm8Sem0d3+cbQ+HkuA
NMU1CrTEuOSf2jSs0HJR7dwVSRS2K19RXI5FFeD1gH2xaWzDx509YbyjGlqIRxYZ+u4nWawgMbCp
D+FAx/H2toJOhbMUtnStGupekGReBXipgtspy8kz72vVBtyhPzEDcqjAkpULLZiihnS7CYm8Bgt8
eQMqjOGvxmjfLOyZ8d79JAR07PTv9jhegkPT00N1k0vpxR1b8ofN/BKUJ45AvsoTJgemC7t+bhzo
rRS4ZY5GDcaELQlEW8xvIBHmNSc3ZMssfzkgezt3UFUnueIcjeOm1sKWcBZR0s6fvMMuMgy23jP2
reEz9cs2MUhVlR66ZY2Wrau7RaAU0gCVtS2cuPx/h/j8qezmfqc7jTpmNvnA4Zs5jp9CJbC9zgNe
Jfd/fRCrDSox0/jaW2EQoPwBwHHtwAo4PrKO48AGR873lBt0MdqUMM+Kshdd/k6V+aJGz1nKeBBT
tUEgrGcx0vCjdPHh1kIUC+AuxldqYnPNYbBomakRiDMgM9nlevisrGwhKhUanDLnWQraUVC2JuZW
NvGWCEPrGI+yE4r1B00L5B1NfzNw5ROujkqVizVxgzv+EJkiU3ZyrwjfMdY6lR2WGHuztFbOZU8i
DIH9t11v0ifo8TUHE8gTAPYC7A/UzgzLvhxazfGbBcW/eM5j0Gk/TiOeHDAqTPx8z9eq/j0aTbmK
raMtiZh6KCtArNJOGdUTxJAyk+sRaj1AVTqvIUpTL+zRdmyQN81LWJnjx0bBgmYXYa3gsiDN7DXF
IwLGcQp881thzrEIBsaBMrsreTgzyKcU7u326apRFkWyxhSj03Wg/FravUdEnfgJPJl+wxyRcG0q
gBzW/1LT+YLi5IVEeEEyVhMAKsM/NKUUi/HVDYFHy4xGUfHMzvBpPRgotEfNBuRAd9KhVN+RVcwh
YXWznPejm1XQoLfszaErUwG+b762u10kX3rXg2Njn6Bho2Bqby+B67jkKvwJ5uG1pBOZMZlzcj2v
lg5/i7mn8vCTuK0en2fW6L17Mm789GleOX/hNlBaxHOZTRfRDy8k1Gjdkom9LtLtX/HcN7ykpSWc
26fiKiGvkceT2P1S0eNIABELNUMdlAZgU4sKgcpy1/+09YD8SCv+B9uBmmhDGB4etr+SIMJZuqp7
Q3uM6SiLEADm0dFPFnBxUoFdjFGez/0nqiTcKIBfjBZCeLoxYjJXnG6iecxigRg1sHL9vet4Ewxv
VIBuSFkkoXxb8GNu4eF/9HKTJFseoP6xdWAlWEgolj/XJalR0eBIi9Ci8axa4pnyZ5Ww/hL1RBdx
sq1Ew72DHTqxpN4VDl8AH90UK1tc0Ku/5V4w9Dg15pX/Q85UuFA+BVMSMC9Cf+0/oNGdfGzgr4hL
sCaeS1WDQAzJCelWXKm94jl/nTANLxywW9poqx5ki9g4og++SMNnl37M68WCKOGRVS/Rfq7WJb5F
fJPvYWGbkgRO5z0R9TTNxYqJ+Ec/3vI9mo0Xovn99WSjjWo3fCPGBoLAwYQ7tulb/xlOhbYsbv6k
CFYfRcuFnV/ZagleTfLpDXQTcfeQ2YJ0tphTK3ZIRjXFxF51+I6gho0QcBeiQMMyEsX+uf1QZsiP
SRJl8fLIV1Et4QiTfs1X5/+58myhNEDDXmcmkjYYfQzb8sen+SUUzmvcRL/NpEBAJpP3ioPZGqUp
p5TYWHaAybLOKpv01BD/mPnxO5YryDctApZC+zAYKed9xdOsaFnMpWoXBdKVk/uP2hsX76XzoDRU
NMn6/1tMIUHeaUnh2tNUwfNuYV5F8key1mxzY/kFAz8UuMKnC7v1zOEmo0fU595/6lrdLeiM+Btf
BSjFA3M72BjcBb8szOy/R7L0zwWdnruurUMq3/FscQiryXa5CoJIhl2xpAp3dnQklQZBciQ+aLYk
XNQcgUtVX2ojbZceN/aww8nD9vUW7j99gntFiP3Gxpm7rr5L4Zhc77SON+qsxbKtjQvhGlLA8age
Ap5/1J08/KjINtCxNWczIPqWf5i0RflToISwl7yUyN1IXD7oHiXRjmtWGVkofCVlLMG05xesqBat
RgI8UZOyZPDyZ3K12dXZ5dHKtsicuSWV5mpRw7P/1dAHnrijFDHTiopm9qcRm9C6fKVRV0OAJEkE
NjYAXuDKbgRKxvjyy9O/kuXBPIIxyO3wOVi1S7EeqGdVu76p6QgoVzHhYtRnGpL/Fw1d0AHluXSq
drJH95zitgTfTLRArP+UGv+JV0eaxwNKIUR+oUTCjJ03DUu9Syu3jkbShup3eIlmFGuYQo1vXBCF
VagkfwAAU+zLhcp2kqGXvJOY+7/Pc4I3ZiRoso6MxAXtS4zOEw2GCNaQGzXcb4THyvow2ph44z8J
NOHt+b1FbDMA28OjeVJHOdE+6gAu2UQifDzrpT6WaEgCOcdOpa74g0s2E3P5egOslgGauOgIoHwT
N78I7Cf+ytzCrACWbW9RqI+HKgSaHzQYWokiMAY/nCk8lERtqK36ECqYdjIy+jseHLbip56oOiMn
LdJ16oC2OvXV2fphM88Okss9Nk5jNhJ7tqaspCSYe1VqqpPn0ZhEWJp3MunK6WEW2LAU6nqfI72P
I3hm/Dbmj4KCLHr4qPQNnFip/oR/ykcaLLwoDWiSmQ7tIBHa4pNYXsu0tj8rBKNm+aRi5MxfidYr
PmKcp8G4Q2aUTRq0BgEZ84EnQBFgxL+8u7zcoPqiqBdkKG+cPGRH6RR8q4LRwo9Qhf3OAXVTxt2c
Hw5VCFabYuOakpTRTcmkMnl11KVIW4GVsO5ym3enEP9hnCXqnSFoSTVsAUd8VLSo/J/EEqUMH2U4
uVN959Jc5PxJLKyKaFiwnWxFHIzHu1DSKktfu93JKuQnaev41qsiwWQGQlW7tDRjeRhlBvUKLlkT
vNNMDVtVS6qloXDaRVTz9L/6DXlVf4Kb2m84iar0jzakLO8kQdnnAlIItHaFJ1tBwrWlv4Oh1qYd
MWBNH9iE9obebzkOQ8fnHxz4KBCCn0re7jrA3LdcYgK1XW26VSsaFDWCiqrV0daJNZoWeoHwjZb0
6+ap/R383/2oSA5DA0i/J38qsX6SBuY6vdcNMtwxrsGLx1RtJLnjdR9qfU4DsnhctGJYSEbzxulN
x89Nun6VejK7K8MrBSWxTR54iz7TOoukt2VkTm1rc3Av1OFvhYuU8rEHIqgWUYFIjO9IQAY4nKLe
UYmqz11uhwbw101KMRBsmuivC193KMDwgLD2S5OPII8AdC5HTQ1qRQ4B6sLVkyt4V9bS4GJnMTvo
ohnqAPkynSP4kw71yK97jN4iXhrUaG3MOwuYlHd1Grl23kkaU9bNNqg384qT7RMgv2iBSgqXjJgW
V3WjlF91889jWHQAlyxXdR89NMH7hvQ55LsPRSzVMFHtHQEGRwZRQjXx1kUtMnKOlo2pxCVhE2Rz
hJFmYMJUtWSf15Fned63SQsQ+Qc7Xv8+jUu0mCjLDYhG2h9CpCIS3vGXPfNv0u+E5fmO94LSYof1
eJIAq6ybgkmKYYLYE3085O6ePYf80l2iUcdQBiD4JsWpbOdNmXdYNy3BRVQB5DzeAwScZV7TIULn
BMDPI+6V8Ppyh9wMZaogDRxJl46qbGCcQ7DqhxFhG3DgGCsDqf2/nd9k7SuOmPE8mhOj9qDoiNt3
23x+ui3PJcJyFQ9TSZJrCvPuP9HLq3XzWkkpDdHTC/8/2la9V/o87bvcVEb3L8b3dhl3QeLwP2zZ
kZ4iperuua5bCE/0z1nIuisBgADRktpQrFzXl2AsXu+nO0imW95vltWq0vrf2jN7DjHH29w4qU7n
GOeFdII/hRae3xaGWNRsITfRk9PWSeXiByGUcPmLXxGKgXiV9cXolpAz2tL8r1ouEMqu4u79thS0
sPbra6xoqyZdSwvNj9NhgoR6yKIsb6jaGVCpK8EblX/u8/KyMTCDPyh4zjhKhr7Sd0IiBUiXCJBI
m56ldHYzYU8o5Bk6wpZOTl8+rhpasZG1QrVeiMjGWVg38lO9zA5PNavMAFtypujjk4H5ShHoROwu
K68BjLmWKMTrK+DXGAZNh/oI6iYnjYycuJYE5xhIQIvyWLj0pGHfo5ZLFQ9NlBwcVkEDvr3CSJhy
/o1Qjy2Wii5Nv/PwVdWXu3tHwjZBcQ2Aj6UzghCAuOW1cd243hRlW5wnuvQVWMFE/GwthnIgePUL
CE/DhKbWOVZLS7l1MT2VE2rrhsFGsW0Dr5b/OrMIFT2fQ5GmTBk2tEbBrwq58G4kKdHOZDBlkMJo
EDw9Mp+JxsoE/5xgftWYinUVzvM0oULytfcAgge/sWQYdBUfRmkBa+FHgBZ2lubqpMY1gpSYmZTR
J8UOK/0sDHBhK6UbQXCxxWCiyW1fgPJT833WoT0ZvnTi1VilHjNQuc3qJC9HIYQpOg0nIkVEJLhU
vUT6fhGLgGra/ikOlGOqPgrepTBisL6t19G4QHPI5R9A9Xpzqq9kmZ1jb+inT2snLf8z9/122U/d
+rP3gctd1WcsM6QJrpv/lidt/qCM8A7zapYjFOgRDG+nm/eGgesn55m3VOG3zjabGwAHNVDyFIFm
IGyr6+IMjIzBJI8XtIT6QAo2NwNSeiBBRL65PhYpke343qOY8UxCKNVBgsGP2EuF3TgJEjiIJonN
mag23zC0MZoCygl4kpySXKYkw4KW3VkTkvRA8Mczq3I1BSUuZMA97BLxpvF0Ty/Er8aCFlyat4xd
a6xeLDxB9DTrmJOnTEA1j23ZP5LXJTEntH5Wldz5310h+2bfZOYhKOV/ldwL0AR2fsDM+eR1yBWB
k/8cybK+Nc/6YjO+CSvyhx0wimI9CF7tdNnMUc2WHOdM8GFJyaEIxH0WKT5OcJW3Xhr00gbDOHu3
nVrPzZ2Y3IOAKf2d9Ps7MWXu5t8wOCIqt34TG9Gw1rrsuDB+6zF2sHyU4mZ7r+GgXalJJJ+ZhMlF
EIK+qt6Tm8BQa5x4ak1b9n9fSPBlw2a3OxkFchGezN+Fyn4w8BcQfU7zWXepWc6utIrvDZAlYlde
zsoSEEJzE8CpB4bHpXWxa81XpTt4gjPVHeYt4rGOSampCnGgWSFgy243P4ef2gV4aQq5TqJZHhN+
WL1s7MopXwqEztqeQ4Oh6QfUu1fhYc3EI9wwv1qJAR9/CCtaTMLvA/1EZprQvYPAssvYyT8AWdoE
6fGDpUYH+xUnU+gIhX859/6O5/0AAAOjXkQxaSsDno/Kr6vuy0Qy87khxm1SzGBeN1mWeWE1JIa0
l6aS78ks+6RwoQ9gGwXsDz+MBRVbA/c9YN/JkpfSyeDXvOS9r7g7fbbYpIja+eXU+c2CRYmtJFjw
pVt/V+FEhfy4TcC5bzNHiVSWiGv3Ljw/7EUdS0y/KQwvz9lKne0ZYGgTSV+uuj30ZSA8N+kWUj8A
mcCOehO6lpO9zyCTz3itsMScvW1owslFBd9JWSYFThotsq6XZb1mZSwp5gmBVfxdMNNcgsVdgECR
db8fv1TxBgaoMTxIqkJIRAugKOaqoE0afkdyEAQ6gQsX+49RCUEisVokU6+uUm4LlqXI5U+OraR7
dOf3aA6K5JKrB2lhhvIn9vVzL+SBk93/xya873GTZjRhgp1uycN1wk14B7TTRr/9TIQZrYSoO/Mp
Ok2zp/MQ5u0zIQphwPJGTZaDyJ8z2B0gghFgJbxnLLKb0X40rpkf+77mXFqv7lUxDL7CXNMi/9g9
K4cPvsEYTLcaJkQUbXbkKrLxtPHsacLC3GmkjIulhPmrNKyU3qXjh9/+XEGzxMuT1aeTdXCQ+yhz
Ycfo7GjKbsrxc5YEVuqr4FD1JoFeXLI1eVxbJQ/xAysPu+gWItTBImYlSfbBv6Bh340vTsKmx41r
fRZdE4dcP+CsiyTr45dTzxL9IHXFjWOmNyZeWoMFH2AfJydVL9x+gEP7S+TR5eFOA5+Z+7Y1ZvQ0
tVU4fJ2RWhtIUmP0dulQjFzFJ+jB97EnAyAGbCKyF6XlUCFaj8/kOLzN8LSbRJWzj/yBi9Gla8iF
tpFvZff8kTu8eyJqs49N5T6bOHhfPGnokYTq2M4jzGODYlpx9yB18CpZn0Q9lNkY+aYPV1iGjNnM
pcIDssDTe5v30PKpBro8dFMyn1zdlQ2Hqn0M7aUnIVk/GhqO3tlTUnm4WgWhxOjbrhErtSwS5YhA
asAOofrXiVJEk1Dr0TJm9Atyaea5ozCq1k2Umhui6cnZZf4cQzmX3XKq6YNUhNBBfuYlbAGUo/ev
PTVe4hCJN8+0OqLlw9cbNctBE6xcQHv+mIS6kg+reOXZVbMeHIN7kKKjwXbq5EIbj7EQJjHFHgzz
QcyZt9sEc4sYXCwy/COrlpNwfuMMJHTxeBVFybOgwM+l8jBmqCSmTrzdjxiwcmSnJWqlvgzoy8oy
6BVf8xUTgl0zSsI/h8IyM5KjtFJLXZch3B2NK/OurjVUtU3FLBsbCEQ8GjwRJW7HX6OzyMjgAfRC
mhfcfd/rpUoeitSpVg2XJniF3B4DVpE+JV744u3x0l7UsPRui3xA2WTixQINeRgc+Fb/ZIQXV9v/
eXz5OyaEHtouBaxwfpxrLg20sXzvGwt2gamGklHvlMdYogoS083umYSl2stIzMUnHSLQITApCQqS
GJbdHZzzeAVlM3/GXSpLz6WAP7gBSo8fvg/meo+7QYjK7LI2jKGIGIZ1N+un2Etc6gV55fxBYpUG
vvFvTcTIMBt5BgpkwzUpHrPmaQ7SzrLqOb9x3puaXr9XHq2MGjd71Pgea07TY2TdDqSUfs3UT/dR
osApq1v+D3F7eD5VFb3IvJhhE2/yf1YeK4TXVN6c3VHgTn0+WF4EaDWit1mXz+78rD2S5/JVg2dL
+6BA+wAa0JyWXlu7nPgmaQ/vS91v/9/6J07RR5d0z18Vu6MjikPgInL/dqmU+OwVXnbahuO+uSDY
FucZkIm7WB3pdmUOdHEOMIwDOQvavLn+BlUAbT2XtanmTXqv2oE6Nnyktf+PC6B2EKcVLVXkzjdN
r7cNkcGsaWUK418ihhAx5MdCiexC7YCEXNeNOm1s2QenuaHU7RxVOzK9xQjD1r3ITti+EGiUhM2W
P6BeyTEHI0d3Ic6M88OncenxAG9IOIH/mFZRfXTf4dcIt6TV3CemOOk1sYClgF1hlyxiZgcvziew
wmEE6+HdU6FWWo52jqPSeD1QWA2PttfJUOAjgk4tajn2OQ7xoYLC1ctYsl6T4pEMotb0oqmHemQt
EKmC6s7biuknnmqrSMOZddI2Q4dBYl9JfpNDtEsK+h5cmnwS7tZRjtaF5Ia0Vfvio7Arzzz/CnYU
Gac/zlRp6tWMbiQ9KczjVMQvmnymGb32ab6Tkdk2WodyM3wXzlMPZ7GHfIZDSoJ7GTyHnRfwBc6l
0CmpRUuRPT6Xp8UE7st31sx4DvdMJ48gAzz9xFVlIoZcROKbsmZGYEGr+wE5R7rhJAdfS0W0NuM5
kygs5dbOwV9zBDRU8QFgymj+gCXG8cIqBpMLMMBanQt/LsklibJI4EIPX1qEUpPGZCPpINHpQmad
vFOv8U2fdyXISl+KFa17qkSPMulwvlcsZUrCNM1OYiCq8EOokHyBhN5hbRvidr8EWZ9N4oTk/PvZ
ytWtO+y1gNt98/8k+sEccc2QzC1T8I2XS1iRB4oekwHFngf+Fb/NSu0WxRhab7329Df6htu7PSRV
hus8lYt2G9g6urAdBDlDLOeS0eGf8s+EwdkCSQFGPbxfhG+0RocRKsvWPg09S7iPVmHJHMXinulC
3P3t9xFtmzfbKhEnaHgS87apFYd7CNc4JPiMjtI5HUYETWvTKx7KT2EmyzQEc+pgMGc/WYUmaYM1
NV/Rab7Rm6Yg9sS6TV4SJrq6pvgumINbxwQM+mkjwqnHNaVW1ERUU6Pmk+W2DRkNoH36rf26b3f3
a3iH9VXj88Lc83cto4RjDWFWTEKFpPTd1V1P4pAXir/o9JQaRRIDXR8DQH/5VYJNS9T1+RVS2YxN
Nylla9z/ZFVP/IJ+6IvBDcXlIXGdZ3KA88gPszcCETAZz2pK3s3i/dvRJ/6+MoIM/bJEO3ind43Q
iAKXQXXx5fEe5EkwfgA6+kNN3bLZhN+W7Q/XekQ0chJYsmfJha1AerwwspLREmH1JxGbOoOVU5tc
OvWCsfs64xUCIhMlv4qL4ecozwCb3dLT+zwfwJXbNLl+sRbFT7EFV+vHPBHsuuDmBfyeGA3jqnpZ
+L1vGUY5PklhKT8mMN3lxFQlOs8P8TZmah+57/jqPGO20x3zDE7zW2YTORrnTZaShpRkxtzQZUAu
E4VFm+DT8rVSq/oZD5on6OGleEuglmhK4bixI/kchQc1i2QzZv3KvAf27oTDHg5dUoqsr4ykqkYf
w/QC9ZMrPcePfuwQCOCGzwONTCH/junH55+TnwQk1SDkSJrcztTA4bROZGsBNRnmShnuC+/cfVFI
Sb8H2LWW3awTt13CbeErJULTW5NpcsUrH276kY3bA4TlvvqoTt/wYyEvgxYtQFP0pzGrVZw6sKSM
zPjKIAZ47q1OehXk64f27cUc2g0j1PgfMJ02LRioVl1XGwRL1j08mVoDrlQcTXJVX3Thja3WGofd
l4AkGI1X0g/nRW6eu86qXFdhz0lYxQ4GU/FkuGkvTBjEybwbnPGbtS+lfZtf4xEfqfq6Q3GmPZSF
V3sAsjHOt+qr+2XX51ZNUqS9JucL+9LifVOhB/frEUdapC5yRfTCJZFODy92bf9UT9sMYefp4xW3
gnT0onaFw5QkvFmxhHEWzroNcvtuQQc3qgTlxk0r62YDJZRz1LEljAXl2e5vdA11OKbb/sULzeZn
XounCjrkRAy69593NJvDZr8PZ1Jw3erWjskJMz8Z6u0B3P50yqnx/5UX8tGl/0c8NzO4ADcYjtf8
hLvIEoCidstOFUbap23XAPEiENk1cI31wtzl4Rp3t4IAPMTNkyWhUChtDw8QyJkM1sOnqqNh3KpE
lSIwHRJ+O9O5G9INIeg0+BYK56eTNzyuWgGHOvMhm7oubtm3DFfNiCRSMRW7fFTKUV+qFr9ENkNR
cW/BvMrL0f2ozv3h34iLSuqM+0KNZbe9LiNRL6KKlqX0YRUDmzE6qGDq9GYcVCB6HqrPWn4yYrJO
Xq0HydV2LAJNEcHR4jbnfNxg3sXe1MnQRNgIRqNHguAH1iuH2HbMTUp+k9haVc8V1+LwjnOD/6Le
guVv6xUE1z+8nLHoR/HNDWFaKfMn8UXNA85s7SXBTy7gLqA3as4j0akuekc2YgN/1voST2GJIhgA
hiVue6FPTFUATRhj3MBj6ZRTfa5PC9OOFfy+npe/kRjLuH9XtggQnGYGevWOTr5c7rJ4d5ZKYZKI
QILGrKhtMqvHXE8BOILrAZmJegRm4OlBAkdSvpAz/Dv7qHlg0mA0VzREANzrwZYi6YPqw3Fufw95
r55wCIjYed+ZsOAaqMurAz5oIXgOXyTv+jfW2FSdQFxsPG6uM51C7bLd19IWy+7eOrToR0oR+zPR
ne+iIoet3hI9sOWv+A6yGvBwtWOe5ZHeAPNtfI7TCj1dGYBnQwb96nmvLZt5twRBQRDKwvfU343P
+xazqPDg+mybaaTQI3yLWq6UHeBYx2MJwVeeo53Pd5W+Qvyr/tRhJnfa6cwxCykk33l886hLamVp
w15U4LjYOHJRTdVLyp/dQXU7GJk3qbikNBucMsH2DsacDmnsCvNQ9+GqBiAUg/h8RjNRwkR5K4FH
A2uqkEw13oXxy3iOgpTP49NtwOwHJbHqAbdir+br1MN2sM5MCudNJPT/raQ2b5dS7L13ZlGwDUQi
cbHF2IIJjMOu/1Wwk5InC8gTg++76wIwhgfEmsoVo7rxyVOev0kD4ZJmevN1dl7oopK15+0GWJnc
9ERQxF8pjmVkKmCKoh7vI9oVopBh5Lo0Ssu+SzE2/dmwGkKv5g5LHuWOp5gJVYNBDTTu3m/gUgun
DfQod2hjpsaxZWgBzolNO2gDAth5ksbB49Sbun36EhiSHNNHXzokjXRJAGn4pbGjqkpS6Ygq9Vfe
93SaSF2/GD7cMkQW98DCy3edNEsL6vXFXRAuhv/yMcEHU2WXzdop/vFGk1b6WdWiI6ibHifiH9LM
h67RONZlg2EWg2KkdJGoNJ69TC0nKTsv85/lSOeZhsV90aVK748jPXS8i1YTMIPyulVt8WO3dekk
09+3yXxC1U798N+ce7WRfpsHhNMy//3g4NoTqDzaBbrc4xjHIWLtxFqOVTWMhYjwOxC1MiYe1IHH
eJJTfHLQyvr0mvMbmjjphxZks41e06PKzwm1fIzS7D7DNNseyFS3X8ndaSI7EcZmwvRr5AQn/LZ9
R2uzMz0af+qMNpizNMQLlauIDiOGA9BMjleL8PYDI4CwiIkr9gHoS1NHv11PoZ01mvAYzr7NuArG
doSOfwHgALJ5m2nskovSN7pQH2yxH3x+12iVO7X8fzYcUU7+TpuczGePuNtti1Tje1OiXdYz2rs3
+JUBKa4tBa6MjsYSbEr/r4DOk/g+v6s+3MBelk4bdpYH06LOrGXnfdSu+lsQKe3a9PVE2QcAssBb
hVbaXxcpOnMk3dKeDDC02imQdj+4LT6cPdSsv8dsd4SomBXlMSLxgc9HP9UzrYj+HMi1kA3RqINm
bLcXDO2ksTX/ep9qvIUqrjWedaXT6ILOwiynEN8nyCSR9r5MGh1/+rvdOrGBB9cQx2uyO4tAEKNX
8doW6sGv0bflsZz8fEXKOVNutLHAlQIeAMOFoXMTkXYdhGun19LSt4Hd+L5p4IQmzjBruLyeSkCM
gHj9Hlg11A6nigMfkK0Gi9oNa/r6m79uMC4uwYOZCNKFpS35Q7/vx73sS7KL/uH6TzpOW0A77Nxu
fXV7g+Ggt845W+xKHD1/jP3ob7nlLITHTsudQkgUv66GPNuJJN0Xhqwrn3xXWJB7kJYrKlhXKi2j
P8jZvs03n8WlVY1GjMl/KRMzVainml8qKGXcl6yqiTKCv6l00P4i/8PVIHMTqOcssJ1o8UneOCDE
ATlTUyluWtODaK4qiMArXGYuGckQg87uNP1NcaqFttXeYTRjhm4fUIDVm2j6vKta6ntVVYZd0a98
6frClMiIsNYOKzepWFKEejzvW/Kvyab97TGajNF8scdnu0gP2GP21udwLcZ4gE5sHrFJoNz+HBJw
+gBzcc8O8QEOgWUqI6WKyRj46e7k10TgdEjI80welWHYdDx9rS1PDyjhbNgJuCyWwJ4KzyNUEaWk
bNru4mKtzvJuDuf/SOMP51VaXAIueKjrvMbcXKiM8dSAgVI7v8R5YBNQcStKbbLZuGDDoOSZsLP/
lyf1lYOeFHeeB43OQQYcCYQj57l4twlUrwS/n1Ui2BsGSId+3PmlAdamC66ENswzfWociV4JSjqb
uJjwIBal1pgbZie5HQ6eAvFcrziWiTTs4nw+cVC+gp/ASPffvljXZVZsphPb0yXwk0fhg12nBZcp
9SMNXuWflg/lNM8cQa5fULoD/0lTSEnc7goqasVwuZ1y3K1YXKeZTVYNfSJQG0VovRLs6z+y4w60
hnG0oq+bkVTXRPGVGo12sy9RgeauRsIkTacwc9+848X4ckebDtiVVGLed/iHd+x6N4AiwxRHLSqQ
mtxtwfuR9dSNNW7dMGcP9x5/5lDaVAzT8xsclscyspBSYQjRQMCXicilQrH6hAyV8yWbIkyPnVoJ
DYAC71vPMuD6TwN2TOwpq1rMDjgNIxd9ZvO0trpAkxGA+d+Kpb5kW/bC4XVaON/jQxC+Uym7XwqB
CQtBLBRqXGQF8u1+5kUGNopamCVGGamRywaxdIuWSnAMXrQCriWw0jzBGytOIhLT60TMjUf8ovq1
kfK/StwAHyVTBLsa5lFHDIALsHFw6w+JXGpfeVhf+CBSsGokj6kG08gYyDcDI0Qz8eDNfv88Ekw9
QG/hWrG2G3IfDHSapJqmwW04h0NzutMCg277M8JU3SMaA89brCIV89Oo5TPdtvIlgQRr+Orza5rH
t+wYabCAdMfzolLPw6ml/fARoO1/fz01nybMHbQFrJPesXt0Lz9naD/hh4FBlXHRMluYYW06egyO
mn/eqttgGamnPwarMUjk34CV+akjQeZmrSANigDVeFFmI+j9OMrtphzkUSNvUpE8Cfkg6c1iWGhd
AJB8qJjEsL06cnyxvndWklGGr5dRRNLtLYmsR6ENcBKlbv52GXVv3Q1lorXNC2LtM+1wch6BsQoJ
jvjS/yE5a7MB/dPBcnveQ8fBuzTFGE5xwL5cKYRlo2P3NTPmbE1Frhr17S3SYPKqDaq3LoLO/val
ln6hXan+rW6QRuXcAaB/D9ED4N6zOLqepxwuCMZ1N3mr86AYdAegOSDF+CqDR78keqXTB8RLZzTZ
a4yvMcOs7dbNcNEeD07vMxidvgkRIub2dL5ApvY02kkoNV76Jp3yUlij2+vfVjBU+EhfakmqFqjw
nryV042xTofaOcBMOkRadEXVEnLJHkANSTcJbVtxZXgBlpOSgimIQT2PDnJQSRnirVEEHbSALB/W
r0npS0RjKoMvaB9lA7zEKEeMzdAR1m3CpXHhKvb318nd9vDVeV2eaBUQgqaS28hE4JrFlRz5q4cj
5NfAAJwS+F0yxUHFY2vJl2Cf2fOo7xDeb6aDYY9c/O2l21VDHon22F/b2MUe/u25SMGmZ+9dHBIN
QbBnTUxXRndWYbPMo5ZJwFydTJdDun7PnoOmDvhYRY0lBSkHWweLb20qnX9z31AoirwByQCfhjCY
gt5UTIrasxZKgrjdyyTq4mAjZ30uIb/41LahTprZ0y6QODBW7izHWZsooEREkwtIJP3owtIXvw0U
XmQBPHtHf6Glyg+CXrshAhClCNTWwhQdZ3SB6xSl0PhAV7Lm9nQvSIydJIaheHD4MiZTR2EAkcy0
jmJdLLLs7MvGNZ8OZrRxBe5oBRzzC86EkpllF906fBlXqngDBGEzW+a9TLepJeVpYS+msTJwnr4i
Ae15Lbrn9fVqgE2LheEchqlc2AJsy4XImQ3weSsODoJhs8G6tabzet9Akd6zR/rh3IdvjhsyE0Bn
ktzgfcniFTc8nWTpIPSqh1eBEbCvjhhHpQvSHbKK3AhRCkcqZv7J5e8jvjpNx/gRQEq7zEOTY5jS
UfzG/htbGSDWGdv29ehCDipt9fT+fsP/VDyvcpiTNDKh3nz9/Y1QJ10tLgt26V/d0RDbiDlTiExs
HNZwF9h7vQNkWtpdosQOFFcWJKO4ZIJMF6CLkgS41WahOKTvCvOWtrCr6yXg86WGac/eQNjoTBNa
Sayz/KX86VILOxbWW9/KeMjKZsUor9h2HmbNQm3SqU6qNRH9aP4NZ8pl5dEkcBRE2huMNr2xDm1M
PGVWCpCr/Br3e5NfjjX+yNCA7l9N90tWhf7e8j/mGuuA00G0iZiJgYtXWxYu+YapEQyBRYrO83Jw
HJyw5RmnQV1cTONOKfXSkgawiTodEdz6leQluKlP0bv85Ks1OGM+QCIVidxGTVfD2dcMjgBoKJEL
CDWGzk+a2VD3yCJPWTDUKWP0Q06WaCNGMhAAqcRYaMwRu+odsz67jt6Ckj/Gbq8rI2EJQkjZbvn0
77uihsZObK3mkc8fWdFFHrr8l1lAkbKgcJSSMx8B7B9VMro5z7+adpfGGd8DUEVKxQgDTkoV0lSY
G2kH0eq5zVcxjPXJ4YuPmZw6NFqZm9FJor9vDBhw2onrea4SyDFW5oJViixmMG9XCR36RkPVtc9n
eIlZPR+aEUDYTtiqNGULsIMpAWQR1NdRrsHLrgsQzKkSNcVDf/R+rXL19JMv63K8oP1OhF5WJlHB
yplDXdQGdvOgXHyKG1rmglMFpHzmcGUkFjNEYIVBZ4mAb8QUE4QyMdv/9p46md29b5HsY/ZTKAYR
2Un8wvZp/BYA956CnX2LwqnJMh9Bg6H6aJeKL75RN8X7nVggi/PGEPuJAB+lXn3W2bt7w1S7wNmT
Ow8XwmkevCHmITLNbAbCA86KrgZ1DeuVATrC3pAJ/cWiayPxvz8OhCaYm+DPWlDZM1loArHMNxRP
9wOhhKYdZR9OA2bG7gPBwz1yMydA2TvxUXKJTkz6vcjvuZcTXMMG8o1KEuWZlHLH35HZt3Z6lRy2
kl832Y8AtijOJwvSuJKMeUov631oPO9dhWMbSzzDH3npkYm01FLhlHaI/6mbLadJOjJgvpaVIwD/
IU6FqzwBsa/d8bVvbrWTXMwvcbI9AopIun87nBmxwhnafguBLF3PVWHtmd6qbhos4Uyb+zya1aYB
6BIxVIOF/5RzIvfnLrdu41t8nNIqAkFjIKjNaHmLBwgt/L29N7ifhBtkUmoXsGxPh5z7pPXLIYB1
k2JGZhb4itO9M8Pjclw0+VxgPHNntOsFPR9F0/c+VCiiWfEC+FlXICpITXdGnUAG46zayEi7vOza
9Xj2tGaF5naSk4T/CUebmVOzj/Or8oJjO66sk/8qtM7LTflb6HAj4cpNv9yJ4AIC0qQeAX+Mp3Vx
Bd8Uyjs0d2ayOnl/XHzafFPaIFrpxPasmkO80hBxujhzNwvGk1zCTQmBGApNHG/Ef6SzIU18Iu9l
BtUVFn+/FpgFGchX7stmEec4le9ALtk1a29yGoe776shVwmkYQdi/ceC/nGHhxslgSbEMfTBiivl
Ov6IDeVtNN7yoDDiqOF0ORVYCqQCn2OfLG9pJ5aPP0+Uv7FyQBEoGKhMxr58IJUvaiS38MOulmdO
jafdNwHNajPBfUaLuyI3aQxMa832vV3TLqkARJ/2/Wg3dvTbWXVTQbhq7guZdvr+xX43dKfPVM2Q
LLr/69MpQX8KUgekEFji8DgyKgwfqhduvCLgGt6/rxS/3peyX/HjLNoKZICDbjv80M2oYnxN/I8S
adS9auMmZlUnozpYZXQHw/qcX78ZJkbVNmGNs6e1yIWXXH7aoXmxfg4by9XB2OXJiC8d6CwSCDri
tsAIce3J2OqNGTkb+tpeEgIH6l+y2W9WXfbrd1HeAl6kWYDYFXT1/cmt2+zXtwd25un5pzI2DAOz
8NriUXBRz/Gk2WKYDob3t0s9O6UdHpsMrS3FNAnNrPNqoMZVC3AKG9Kl7n5cE0GS/edjhaIljCOl
2ylSelDXo1JWT0QHwcIZTHxhJ6Bu2v8OTOiZllIiuZocF3jf1RqOXiNvQdYcTTyHRuu0AyIrRCCE
jzKBtYa6iAbrxlp1M7ziAvbvTJsQ0wpSvBih8MZ5geut34YPuaw9E3p649qWy9VeCIx+wi5YSdW/
bLiEc/rxpTNvJ0l/FQB2HgcPEkHfjXbXDjvxynoyPYDGopP4MmB9I6iteVW8UBg+WNQse9uW+Kb5
Ny8PpBqVljVXWDivVyu4I+V36jLWX20Pk0EnSVNvm+JeDECnNXCebjz6TIVd8dlCkf5Jn3XWG33U
x/vb1DO9l1I/hRlDVrgR/4TQelP01B4jqywlSrA4miU41T/xsNbqlycrJowLjJPJELIL1nqe2gQo
MZJSJH5X/A1pHXdumOEc4y/zMt6Z+lbSRu47e1p0s+E4zve+msezr2vSDl00joio4aCtENaqXCIn
FBg476LcmJ8w55rZ4cCO9mxLvIhxZC4rzTMzOENegRi7rBzwtu2klOnAqYzvxkF1iUxAs+45kZF6
C+Y8gvo1m7TE9aLnyFG3Qvqh1W8sCrz7kK2gOTSrv3q9yDN4DXUEDkFyTLUIYtJp88uwQZPHr5lP
9kbk9LQui1q84d7A1FrJ0pnp0te5l/8ftqqIualVTDX6VAWT0PALUHh7XbF/+GvFO9zvLmOVpqJe
DtB+3y08zVb0582vUK6AiOeiM+HzzJxsPSaO1P9fyxp2O5EqWBXuoLqP8t3NB8TOOVmxDP+fhRo4
9ImPxFAql+UQF1Wu0eKNNn6fi1L1cuu3dlIjgknz26t+aYXRocvs9k00xl4znIx/MAgoPDeUU2PB
S+CuGhMUSAonMdtf6ph3WRgldgVHy8Q4lqF3Ge82D8/i8R46DaR9eCY2pKYJOVCPcWni6YJ2xTnA
m5mULrT6GaYnScvjtBT91MzxHCQunEQLktuTus49yr+ZSzpjAf33mSc0+S3kqgZQIQYW+cBNdBBQ
w9cK8WNeQzE4BFV3fHmnhiMezP5pALMXM/oyVNIkmJ3FsYf14/a/3j0neBcU6ezbGy2XOULhMfbE
AouSktUxmRNQzKb1rcP28SUlB/QjCex4IaNYGcWv0k3oVwDtlbEiiUhd3gJYHNbjd5usToI4XpkB
u2kzMO+jZ/cBCrsMOzPB0RiE62i+xXqyJaixOGYhAQvY1hkPu9+s9fbPx7WxU3ZrW/TBFt2iB7Tu
S16ZNbJLyIof0Grdpj6edMafcputRIWiadDpTXxnoBFYZ8IATu9FeiV1JYWJ+7t7t3JT3YFwgRBV
kSQ5TmFay1RlN1JzHtL3WrHNGsBvQAdksr0hJIrMh4UcTxiWKRK893W9JM5lVDybGaSt+j4lxH+5
rqCnHfNzMDp8bd+Sh8jGtUbwz2Y09i1Ac3L5DMiIe1y/FWBrQMO7C37eYGAGxqOSha2I+znF7z2i
JSuyo/3Juyl+okoGAsho9K5NLjHvb4IVxwKKAuC7vhQFTuh81og7iZhfFmScZ/Gw5romZLqGC4CO
H+mGqjwILgIU/eqT9qDzpvr/doKg8HheS+1mwT2SBeQjTET4qSCCxBXcbtFQ8BUQafmVHN6cMLB0
hxOPnDEgpz5QjU37r1wClKuFCQkApqKN2WFi3R2mvAhvPzebnkMMzT8IQXKjm2w6ZC6K1hplMihC
m3yXY8qj1Eb/Xeip0azMkP9xyaa/8yI9JKS+wiENRZZ8PhRBfd6wnWnECLdjexXB+J7f9Ss37rEk
YYGDNA2mXHirjBNcnmaORIA+fGIZk+y+AbuVJTcjJ3YnvfZ+Hm+3JzGB4Qqm/qyAj4lPazVhkylb
ZPOljfkbUgQsORKFWo1oJcgoli8TWeShApmjd4NFwgHX2lDgWoFNonAgm/M3QrisUqYUvFjIoO5W
41yoUISxvREWS24o/W9iNr9ja59Z/5Wl931w1APeNpErMU6pcc5BzI4wAWkObLVRdJvFYG0jheIQ
I6eWGR0hHsw9Hu0aHtX/kYpHgAw8Nkf97VW5F8Jw1BeuOGIKufweWTsjigY5Af5LpNAusgjcrw0y
StyedTnWDO39xKk+/7zZ1Fr5Axau74QNF1cIR8ijNqeuBVfluqTmkYg1iQd/vrE/X9qkeF9dtPih
XS4NFkonFkSSM5G2KtJyLP2IxjQ/btOCX5TexD9Pm+xomiyVa1UWiSE/GxZYbx2MLg3Xlujmso94
IxcuUsuAXd8T/KN/PPQhbBf+i5syjrEiT4SA6GiS0vjADouhndBtSEtHg2tdt8yHsSnEHWdsmVef
7+UHPdYSmJ6ngoxpx0jPRBI7hA+UZg1SEzJWEhPyJY4WR23FtsIIgR4iUOJVXZWXtSYy8NvQqeCy
/swUB4P2FnqzUkCgqm/R+Q0PkTLvXsdpgJdxH4wHm2lXzR8NMFX8fITFPP7sY3o+vZ7VBi3D1BEx
0LzzR4heBILTmknaPCX3CBCb9oLJwPBB5DM8ulOFOeJI9EqhvAWuVrnipm5A74Hoaf+IkcQyrUWj
fw0yenf+77rQqrAL2wG32CVCVnagkJo9apnJ+nUFWpe7B+w8Rupszsr5+j7rB9NlP4+Gn0PgN4Rx
t/OgggOgnqQNOYU8Al4r99ssfhquqZMnVZecWiikNv8BcrM8l/3rGy0+wPQWvs2eoUosWqhYfikk
kA4uyPn/K6Kg3nJU4hpUh7ntu+FW2h5UJmRBQACi6fseArUZRVK5gZRG+SVapZ2HLhUeasYqoK3f
7sAllvSLWP3vhELJ9j+jQXju32x+Rhj8W1MDiUd7GhoG4oY93rRQDbyydiml2GK6iEgGxGvVgRJI
aO8Lx/X0KnEd3IjJn+cFK0/cpAitHG40d894bC1MiO7WLNVBEenl/EueU3f4rsN/6Kjc92QBc5ga
K/XngwugnYxKxqqxz1ji+2KTsbXlpdqQprkDm+DJ/+j4XZJaEqn+ACrfoqBJByHa6PaFF8zBJwGD
GdyetD2awoDNT61qUySdZ/DINqF3KVnK+ODK+e+eOVgvb2I8cbRxoyHDen0n+Sv4czzIIm5vRpZm
H2o59pee/QmTN1XYWaz1XFKZvLGGcDhYqSGy7oIdE9uD5yW0gEpz9tGOdfBYYUEqMnqY3gUTKYYX
llTRfr1JNDmSA95WBTbJt5YJ5ELQ212jN/xGQIFXvFSb6lkZ40YSYOc+df7MnJGGRbvXOxT6LX/I
UimXt0CngbDpDR5749lbm7pju8RVChSH1Fl91OpovnFshU0saYOVPGM6nvXq3Zy1aKy4iU9mR5WQ
KxXiD9kdfll0aTk3dn/1V9LhWq2eKiu6iqorVFEyMxXiM4zKT2OznKiV8yjc0v4Hr97PtCuBM+o/
kCb7w/gC0P3B/sWvK/L0WhU7xX3oELBjsyQ5IKm27QBFSThXW3EFeSGkMaMvzjuJ5OKXDNW3ob+u
SdKstkPMugnlJm6ieKJ0wlTXIXQsrX0X4wzit4ez4YmVgOWUyFGF0GUIjhQVxBqzBmdE03cysrWI
AYFDVqUhCvEzwfQ3+CVJjWcodYPkaYUmrfQR1eborhHMyEHGWFLH7SfJbYJ52ctEfWbDAx2eg1lw
agezPBryNt5luItX41gRgbyYAqbnYvSYxSieR0+Mr3FcrKKpWQklWzNo3Sd3O274HUs/ajZEd0vh
IZtj83HBp77E8E9saZqeC6trgOh92+7KYJUsfAvR7XJZGETF55Eg8KkqPqPSfMla3us4EOlCbhDU
STxjS5+yZNdJExYwd/odOEm3DA6nSv1m9b/RHvVRdf8WXdVChGpDuBI+gOwWITP/XafwllmLE3X+
QU/VDP+qhbYrVkVpbFTk6yejBlNbMx6R6Jdr/sbDom3QyFgN0OldskH9lhG898dxqWaHh1Qy8Gen
Ryi9Nfh9BJJbVsoNSgmU8lSBh5My24wMYf2g/DgfS2EN5F3ZTl9CCXRkou78+z7UWVEQBcMrYoeI
Yiutv2ORlSRTiP/lsl4Ulg1TsLtWcfuhgvAYx1+xS70MnsLBoQmMR4DiEhm47jYPomD+HeKEycyo
b4cjoSfiLf5Epw12oMzok/yOi1FmJgTjHc2yOtArbsM/vQ3IuuKefiF5rGLfGWtd/qeaCc6E8TTD
YsELPbXytVa0LyqKoqjmSBk46BRBWq2DCoqz4Iuhgb0KcZbcDqavCgEU0UZxDL/VarQid6TwZgrp
kVMSgEGJqJf1tBlGIYJOfAxoaDOzxIrKCJvYP7C4EfV9G7jvCp+H0KA1XVp/mTj9RGZ8RdoM1qfT
nzLqvWk9hLDp8y0q1iO2G4Z290Li3O448+j9G4PlA4h5oVICUXxc+HC/PSRL5F3KNXETskcWNmwm
gb9K0JkxvBuMsCc46K/NdQkdpWHE06FDdOTqOfqEK1ORvugvG+gD8sTb6JwkOPnWzAvb/bRGjDzm
SI2FZNmm7MbiKUWQgHpyyJxaNNLfBvheQj/Luidehl28aQfN25r3lil+nVwPqo6nY4GV15bJsZJN
15QzaVi2fhBOLihwjYxhGZjCEfzZ6bpGU8fQxE+Yq1rAGjGEtMFiO8RC9eYifPtM+q/Wuem4jvm/
HQrtWgOKOmjPh6ZmJ4bywmuyxEskWc9Y/qyAdAiNKTPQaK/yJToGExQqKqUm+TYCL+tcYG+8DNeO
KiCC7m273A2Owter5u12KwIiX8LNYUE1QKqZkOd/Xf+tphDnkwin/CosyS6l71rSKd7qy+eRv7vX
5X6tFVZEnT3q/1D0tUiVf8WFrg9sOXr8Mm85OSEwR4YI0snFsfue5zgn1fttArsG7NFRH0q/2GJ0
zosNr7bzkE7L7NUebEK4VZf6Zytqh5LLqkfBixbR/frcDG+Lkaz+jZqjvN/HnQEav7FIyUn4iL4d
xlVAsgMY0RlpDeTccX8QHoTK6YLr7o9riTYSXBYWUrs7xEXS6vVirQENHiCp0qMwKB21uYEF7FLx
zIot8vG3+KcDgCcC+WQxe4mQhVIdmGCs1WCun4GcMO+OVIgnW+Z7Qrpbuhb+aMP5ByzActT9CVCS
xeWXazQVMHwUqPh3Pkv0Jhcxgu0XyljwKpH04tWacwK99f9ibdhHE39iJLJGhOsOImEgrsDSm1KD
OzCxPVphCL/e5+zzrCYEtDVHMXK8egKXpurhvPM8V6xY7gc7aE60Bb6mxi0xZxuL9HzaI1AlohCg
8LX69qW1KDjLK0jn9FwB1/HYUJdpgfeMTzDRxP247po2CV32w9Bve3Xc3vQSvAk+8A0jtHr8DnXu
UNlbbWF8jfVRedAVhZdJz6b5CRY5G+mbbjbJSwr4HqpT6J7jbEPKpTDdnqHvYhXhk/cRv8s7mEHX
//mZD9ThL+nmDZGqwgxZbfDLFsuAHwd/+FH5KibL4cipsGxIfEIq71s7CFJQ0dtZ7idc/GYj+GhM
NsXfD09ZhRnOl3F4mSwY0m7Li1b3aXI99a/k5Q5MPDhzkKhc+0kTLQyQBxJHcTLxfTf0lb0IfG4J
lZNLOVeM9h3sSjzsLQ674TA5IyG6HZ7LLKFQyecKx/gMvGJAbtk6gAHGudVypta+ZWIZWyVJAhGW
UzJB5bqYP+u4F5njtHCQzxcvA9jpv2VzDskU2F2T2cMbpzaZC93RMOBF9larGG47i+Z2fi/3vRoH
RBCDkxPa9t5dgwEt7Xm9ar6oNfVfv62jfKVs0E2ILhDox4c33LeTDBybOhmiGvPQqgSjuEIfOyKj
/vSLVU+uaMSXdDReOpQeMjMhnO+LeX/bUVQsmlwYGpPihvMclbk0Ufo0nxhh/Jp3PalY7C2d+3tY
PvXpDTPh4za3HSzqUIOiAGGFofcyJCth9Mbvh9UMXjBCZViBM609r/JmulJgHKjUvDRnkeMIYaGa
pkmZCriH6WyPhV9DywTmykaDL+XaFz/aZRE4VAuFSohZ2MybWNBv88slOpFbDPpgtuw2DmQXXyMF
PFV96sWriN8jP7b+7t/nnzHGounZZMqjwjct9JgHulOnuPI+9z4+19Pn3WL52W5QawKROimnxa7v
kZe0tfpvKYkchRBoncBJDRZ18lIS6wXLuEhjBEN6kKCo2EtQJ12vvHYC3iJibnLqbUtKDak8V3Ox
+FckerACHoomTogBTHHZVQ9W3dCVB8J8ax1lqRedQv3wVKEgwAtC6jv40Fe4ocijlA3jNAZDbx0P
1HV45viPBZcRmg/yI+h5bDh2qLyWVRDUXN/D8L305gkNP8Bjjj6yk9JVOAB3g1sEE1OKVzTHe4En
1Kcbuz9fgmqasdxeeFCosj+/49A5AaBJMIDAQzw+bojCQushVt40B1HQ+m+kKu8IV4HY6lUuUtUq
YFLouYu0PcHD2qdqI75AeiNlSTt7XOwLGJ3xPv/gDCG6eQjL/FreRmi+8apNH+nWNxlvyfBwi/kq
XNETJio1bO4YfIIf87KFyl0TBUtnRkravVANYevC2J2mBHmkoVLWhfoRJBzirMTNKoZ8/mdY0Riy
kDEH/Or0XLkQAberLbpOrxw7zofmIu1Rznes0DBaK0zh/WKqV89axHHj2KhESone1geUnVtgnn8S
MPyhaSp3NhMVd/lfFTNYEk6jJ9dKhQ/0g0ilhlgDoGZCSPEcjhdfm2w1EHgYmFn4+R7C07yKQSMi
ul34JOo2lSi6VdLx8bZWWtycZfDCrpxzSMp/rTICiEZ5JKiFFLaD83n2DWiontA7KB5rYhI2EIu8
8YXVa3j++gjTQdkz7PEF2vPYlWariBRfoholFBTz0l0WoTGOG4WzLgDGtt+rjZQDh/rhWtoLbot9
Ifxvl2aG1RpobEew1n6A4FDHMoIfUKABIko3gb+bTCixOY2nBTb/rd8BL2kIKnNkYpK/NeH9mwqv
Y8GLGVB7al/ViwaU3coghmT4RjmVvZBn3pDcMYCWMyKdbMf5NZHr7+lynzHzhw1LzE1OVp7fWLRf
VzcQPOvz1/dU4+4madsoKYlXO5X2w36A4LH/CBebS5pLPPJ8qpzkAV2Jyb4/IgWb3SWD/83cTCtz
03QroHjEI4c+BnbGCY8I0oNeOXbdI9N59LJElnhQfLMn5ttDfnlJwg3SCd2iIDLclIO4N7Wncnm9
t52j3zHLHO5tN+/W5AFJIwLW2wvifXEgPgyjQvCbnQO8BggHFybAM3EpkkHQya48RxRJFHCxwxng
nfcLjCMPGjwQMXxT/KOJ4zMVjsiCvx/Jqm5f9A9jD6dSBMnFJ7wQHo58GEUchUDqx2jBPyNnuUTj
v0vjvVw5jn7qiTr9AalU5Jb3n7mqGMwIpunTr/i1vF7PG5pg5vRyVtO9husD6/nFTwhAZMoPxP5O
dXaViP/YLHo+5HaPPotqztQSbGxi8vqyIYJ5ukHbmmixsdx/MlTvvxrpBEw0SL6gL1CGep4Q8yMb
cvMzO5l0d+Yd+lB+RhJNSdaIunBYCgsdRFu3aWXGjJJfOvaRyCmL6Gvh60cc8AW9fByuV+iBTVkl
zs27gbAj9qJr9mt05hwfoeYFTZ+t8BcfGWsH08w9yzwWBcnHgAMRqn29QRWJBXDBfbt5AZwjx/o1
mg44a8RPi1VwSDqj730RpwiM49G2rTlZQx/c5yrN5uHvHktq6SwZaqGanBNm6CzXJs1cMuZvpcrq
IR7A3P/PLZZFJ6LJb4ATLt/xR822cgDMK2y0XmKLGSUU6B7ybakEoIid40Bi76kP+bL3P3yOmTiH
zgDOexohkmX7/NDRq7Mjf+wcqKMEoJVIaUV58IkYVyrbNdyGtYsciQEdaheZfKNaqhhyWjeALaC6
TvpYK6NCpXU5p73uNlFfKCgLHUQpY22FSv6s6vfh+YkchafjfelaemFtQtCgRvT6Krg/z/caza+s
zxoStqlKUN/JMR92Mh06590OkdgkT8bw03kwo3pxWlaSOPI5Gmmzk5gktGVaaDC31uEHF3Mvy24L
U+0dFRwigdhmzJKmMzmMIFb4EKgQcBfEiTwpnvV1Hu2CHRuAz37k/FJ+0Q8CAct5xK3CpD/wJdXD
h55/ubmFTxDMnyb8wrMCrVTn0646+USbrlTGZ5M46li/wmkzZhZq5X6ZSxkQ3QcauXZZSZRV+kLc
zTSW0GjasfUZquqaP5psafwW5GYKS0q0DVYEMDFJGIa5nAQsZ6uY+qYsjPdoGJWSaHUKzJ+Haeue
wsKd5UEVgFKaiLWGAE35iNrrFM231fP49oIPKCJJGOhVUUv4XPilZz4MzvgHKhNx+DJY5xj3wAOC
4ux6/jHKzbPupfmuBdE4WM7Be2HFZsoX2Gle5ponjvelOZ4/3/+eDenNg8yBQsZ04gD3MOKASB5p
pv9LtObAVXQBqGKp+VRPp5BiHitaA2RHA6spdwuBsfG3rp9eip6SHFFbv9ux5apoYOL4eFPdgDiL
wBm4VRzqHU6x6B0WmIRsMa4iwo8qLbgJ/9uAVwA33kImpPQqy89m/6EVGSDqO3vYMm5MTgEVCZIb
24qMwvgaf5kXBifwp4S2uM5YemTtpJM8qMaljuURjztCFx219Q3Bt+wnYOCySkvY87UL7yGPzTOb
Tp/uyIRbsiEMiMi/gTGRLuSUKmOsHGAfLTxs1j0UmT8t0TzzEiVtVcw1m0Og7m+lXc+9olbzAbxZ
0kwYrJAHay6x8v/aH25xyJ/pjfVUSTm0VZm9gtxpt3ltafzQwJddmdZFlKFLMXp/XvSSehECWlBL
PhYJKXYF0qyVygtHTsDPSeIOr5HGDTZNHn3OsgF5IqCViIb88YO2/WQmQzE/zLho/t8QAk7WTsIt
VtN5blbCN0bnlSGF3Z90cXs0Wf0dTcgQZNEhvakigItqjqzIVrkTtDbAxbpPU/qE+bCz8F1xCrnr
0ulyEbshC5swmEwtDDQrHExppsSs/JLAOU08L0CtsOp5lJB1DpMCb2NzzGkgurJUc0tHS6B3Q07g
NUcxQqnzqClqOWezIUTB1EHuijAY+dmOES6QBQi+0fnE0cMWcq3keiceYmvYtMCpdNnflJtG5S4/
MIjjEjFy1OY+KMCqlN3OR4TWggHJgM9jdXVyuCK/2fW5/2RtOFA/Ch7fl6OqpUPx/w6VZZFpjRgF
GT6YkMFITUJctYc28dafzQlzoRiHyuyHn4lgT/UdD6gCcTMNZdFQgukd51DHcL669++fuelNo7v7
bENb5oTM7+peFACcFuEoyMkHm0rE7cZt4pKVj8E1HlRGhTLmMdQVqVkhLX7wakkdTpsG2OHTAUVg
p2Jtk58+bYtVnaLNahfzR8U/Bxxc8WmjRoALWwR68TjuJPjS9h+ukra2rKKzb+7yBLlSj251rerm
kkXvgopUamt4Swe1E3XJVn3RPkSKdQopj3J3b0Ckx1t7aKHWl9fYYE/0+q5MU38kweBYJ238QEBR
Ery4F/LVdFfTegoVSYdMqdbr2OrVN8ajeabykVIVZPi4YWAjthkVMXM+TnbHdN9T9lUj9g0bSOSp
xIhsCGhtrAMdK5JYO3F7P3zF74VSi1cXJDkquAEfzkC4npejhvtWQa1DkyzGWgGmg0NVmU2OIbzr
mpdkRl0qZtnK3Wi5UDz08WEIPSWEClOfDfIjg99lOmrF3/yLBSQ7p2xMAT5QELg6vl0IStlTjEJN
brTib9QbO81T14vL0d3e1TXOoLgl8MdEarPe1cG9gskViAYY+/KP9ATCCacz6C2IPJO4oQs85kZm
B94P3o0c9MVhRdiXHrU0inaDiKICLy9GjqNbOepFnHZqCiZiU7h+g0remWoqKPrWj+WkMIjl/7zl
AfU/p7eLw4EuUOx0WagOZ3pg0qLfUYGTb/boHJWxjifu2JWcT3AsJfjHLSEvvYIq3dugZzfO3RuS
YLSF2LnDyC5gY43O7tx4YaBLj+0BGBubNY7B7cfcO+a/JC/wCpKPu2uXFjtrYqYgi1HMhwxk0zlD
BKAU5iYHDzDfhlO0vIvnrN5lTU19HMivLPfd5Oed7B76uCImhYov1Bw9RmyXoai5f+q+JG6FiUTF
JUDEAnoccDpdSp61RWRgH7rzr0K+mqZqyXKXT50j9IejazbB/Dok3zDORp5sPhlW1PUktXxLaJTZ
5Ott/SMujITf3IzFJ6K9x70hM6QD/kjkA4ByIy9xTWkOhWmfGcAqZ2DhsGrzy2PsqQUIrCLCRf6F
FUs3rTTP5koBE65x7ihvFZw5hNd6kKZCy/1FllZc4HbdZz/5rhEGUVSJm5Kx+IgynI7yUfOuWvx8
BpSUkH5wXBJadZDjgrrANQTtJpQVGIYEHI4hkzw90S1vEinbi+0qwEegpzWpM4eAUc+v76w2rVKn
/RvEdesFtmNfArd3apKH3FO017dM452h0YnxvoPpaCOb/84bbD1xR9ps1Uj8hybljo6QgEu2ZwMl
wEgFrmVs7RP/nIkeRLIH1bhbQDNc7hBr1LUQ7+sf0GruRSMbUgAjCcHZMFQngX5n5ZZTXedPYKYm
nFMQMqxgblLQ+MvqcJiP2neuBDTDSHh7a1qZoXNFiiRrs8mP+TCMgZat2IYS/C/C9Xn8JjKVpuqc
XH/GTTUL3Y0FyzgWZQ2MsuCj0CCN80eN0mu/hSgZ4jR7Wkn3CqlQIYreOgPYHCJQrFl5bOPqfF3b
+BPDjydIe34VCPz0VUiDPBgYEhyHn0LON4B5923jfhaXW42QjSqFs4elGPtmXeSP/wDa19TeA7bT
AZzjSoFm8Zej9XmufkdQ66QBjFSeqYggw6Q8WOweKnxiCNpNlrdzAdb411pXw/6q+h4wfPA0MWTr
WjbMaJ7QwNvfPhjFVLSqq8QtYht4KwbW+Q1QxKT5RvjFAZfpLeq+vBWmUclTkVB/bxzcO5gxUJb0
7Gs/T5b/9ooZfba4px/cx+ffnwvYu6492vDyR6C/klL2Mxmbo6WODPcZWqXUPsvayc4qu2eE/1WO
yt5kvgFHz4i+YGzgudFJ7/vcgdY6YF8eV2LE4FpmZRExg8j8HmnH9uf7dk/c1orgZDujCMKrWqCX
TL/okWRUosXNTamAWVVMsoA92RP7ywbYaDlhKjTJ72Sf/PHtcTOyR36q4Q+FN3nVtcpcFa2AD5Qf
ERMR6Q+Ih8pO246k635FX5lBG0VfFxtl8pKxhWWhnLvbZ0JhpI6OHS5emg9wJ0JOf7I64tCvoa1T
YvvNoett+nC52wcIg53ZfZlngslo1UfBYo8zRzcjqkpRd9qHwArCGledmBCufc1LiLIrEv/YVzpz
dM0i67fVk1/8pledb3gF6U8TZdipEtbn89g918kNwo2NWzOl+9bwYYH5OYq4CfK70WHQod6LMGOk
XPbh06ZqflYvGXT4xlRULsfwq2T5d0C9xHrHFxjfFwoth26Q2CJZTpYFFVpelNAhXzyb4KuZSNPV
ZNbgyplR8cESfPoEzFcnkqpn0MS0to5DCz2etg5ppVz1hZobfs8oK25+7U/RMD5brWMqGfSfyei7
gR7Pr92LbzrjSMe5hW5LFomgwvjLWeY86My4h0eqB5jQmyoHu4+e1m4E/k7OU4cYj2u+3PWxdVFe
IfvUq+YGPjBMNzcZD/kKt2YJPPRNryAuYDX1wrtWZ9Pwnt25j+/3x3NevMui3NrBYzyztbAb0Y4P
9CTls098Z4i05gZDqObBH7GfyqJW2phEz4JZ+ML7TMjAzMT6hmLZygGKxXe2rWjkqwEMSSqmSm75
33m4st2onw9j6DLcF3cZH/UazO3kET66k2cmGe5G90D8rJF3DyNiz8FkeDZeZWTxPHs+bEgRxEcB
V4TJNlzTcTKqBjIFz4lFMzZcOkXcwUNbsLAsz2JzxiEmBhz5udwOV3avzkOh9ilP4I7GWQrmeba/
GgssYNCpYTXawY+nmLEUJdwD2DkYgtgiEj7oggGqdyg3Xs1qGWHxerIT3FYc51HLB69iIJKrpw1l
bm1yKSAZo3Q4du01GdZr8T50Y6qGeb6JYqBBjw4PdjDRu0XJNf9dWoVvu7f7T0h49jSmk/NsxXvS
MH8naP7fSaaDt2ZGLieor93JrCCEx/ZPfRcrZ4qcXTbfen50bq/lfsZAXWnJfAC9EpbeoKA4Ka8r
6KxIPKh2RA4KSO79BxkltjVBKugvD7XH6XGe/NKzCsKSFDswzsv5EQK3RoBibGlfi1UJgXSX2DPQ
E5aw6Ospj23IfZ3SoNqx53fSwcpkjnmSDR2/lu4i/r9aujo0SUvbUPIIuSpuw9EjhJw96/VNt2IJ
WYwTxKrOi5wMn6zJG4YyPk1gK6OjgFqp3ZEHP7Z9Hfebd9DAMN+D6xykXazZmWjx2z8aqWBLl0JP
ODz5kUJbNSm3hHKgmYOf14cJwTHU9IRhHaBY+38oN6WLs+1sBTVS9+E0PelxQ8EhfOQo+rVRawUM
285U1ZMSx0iIOUZzSQwgULt4wzGj8UD+nUZns9y8NjY7ES2adW50VQJi36aleZrhDDy0/OKzru1m
x3RSfHBztlYaMZxTIstv3MVfPp7ODS3cHdtzDG+GQBY9LXvcC5oJFrLTaPwTos9MKOTJAUBTPqHl
HkVV9JdCtzWTOekeBxme30D/FvxojHsy04SKpK3a7rwNKJy5VkaQWafO948OpVaDAsjmdRDDvsrZ
B9VBCe1+pmUnRk+6CIEM2Sd/Rp5Tgs3uXOFdRnTwBuce2zu94hKXAU2q9569XEzGhobIy8fR80d/
MB5MFF8XZMASwNbaHzn3ekPuuRe5nHI7oOiV22hK+P97zRa1CXF8cxL4K2IzZXDtm1d9oOYs9dxD
+dbCXsR72foNxZjimUi5swyG772EorMWz2or8JszycQwMzpuZ1EC1kNhwD8l9C2qi1kMrLsjU+iT
TBXfc9cURP+oGSKxqnzdvxumXoZOB5z3F2ahNei2UtwBt9o5ArLyBAxJh37cWlbr4wBIbBlDKbp/
ELWDszSaG0zM7PaSngQ7skintYGFt3USFwKztPUhzdgu/Sqw14MWEwyc/GK53u2RDpTVA1z4uhiC
ij5LWJi6R9FoessuqDbfhCZbDT2PCxCLqzlLazWVRIzUUidDZtlq2e68q6+dCQ3G0awGui5h3Lo3
CLnjhO1ZKM+0vSe4yl9ox1wRHY9g6Iq69lXaoPkh2uWxwWsOq9dpT7hvdqxg1IODJsD0zdw6zip0
v7uOI4FcD9mAptuSFAopzP9QKUBCk3SGXRwKtt0BgxXQiYUwiWoA4x5P297bohveO3TmrVo3Lgli
0xWUsOVLcCWZr3cD5jH6SJq9zDSatYzbDvHo1LrU/GQxb+W32UP840lErKfeYIcCqI9vzfa6Dh8C
/ZSDDuh6sKR/H8pPYL5hulLXi8cw6ChlejbWCdPUixyRxcvLHcPFhHxZeqNLwvzdwpCcZLw1iBvq
ylbgfT+JF75M3Yqjdv1c8IXgU5A/1p9ZBlOYxhrGL209c3AS2vm+Cy/GFXicFniNpZNjYHp7B7Q6
qQudTxbL7xinldfYeMJYfLTNVeOWLr4EMsgwwLGJhwMliMK/2yOwt1FN/uZW+lWnBe/hVkTnjiWD
NzlzNWYBApZmpZ8/LEN3RsZFix1OFQgEJpAChqQYFcC40iMbWK+bx53aqHAXl22DTuYauOKs79ix
RT7dJl4d0x5psIXfgGTfqP0nQHM66zm9kkiJNiR8cEAB+65BxCoCP2RG06yHTOwAg2Zw2k0f44hS
HA1Fat2EFQczlSG2NAj+tknmToL+Fm180JxFl6VGo1zgEG43zA+PlNBRu+FTbFwvcr8BambpjZFd
gEEXooHl0gFQUKpnaR1DtTFFFsbamTyhX+ZBL6oSplnZNASO8Mls/irZEjFFVPd16MS37PSr9kkV
P66VWrp7GXxnO+/6llM5j8JV5OdUKE96m1MtxtaiYvvJxNQaEHe6L5LeYmXLr43NQxn5Kf9ijEBz
ZIAHBfwQ3GudcOAPI6CoPuK+8vTckd4+XZqat+L8VB02YIYNgi4tOyEiE1NCJNhZa37dziDd4yQq
nSbYRAnLhvsdVYjgFBFAuN97r2hm1hpZ+/1P4mN8lEZ3GeAzJ/6uFAX7LZhFIvdgO58c1oT6oQmL
B5+CpVtbv4vfVYwcgL/CZLPFjq6yjUug5w2HtBeBlZTon+PAKMne6ApXKgACroo7vfq6x06b+DcU
n1/MnmcsTou8NvQJew5P7XmnTDc0lWTmu+ZcN0iV4d1S2u1hq08ZQzoH0YcJUCJOMfazp7DECtho
/f2innIM0+yrOZKHxn+EJHqdc2681bY43oFCd5X9bOP1j1P+IbaG6mZB4eZy8TLli/t+8kef5G3x
dPJkXfO9IerdFRHeOtId5ZfdC3oiiE9e/R4F1tMC2oZPtntV21U4Wb+c/o0/vX4ULx62yW5JHsBL
kFKr7Q4IPklXL1ZlLki3RzulAd1Nboml6Np8LfT+lRb8kwFg4gN23lMAdMDhyJ6oT25Xb5RUwcZJ
Wy7dfFMckBsLPO+ekQorx1PB4NHGpCKK9fZoRcwMuvqMOeNLL5L/5556ZS8Ht+58AqrSUbytnMCy
x1Yz23aAqOCmwZEz6mKGWqOhW7+Z6dFW/K9xYOBwebirxsNkMZFBS4u/jXzul8w1hSXghU2jVnpA
U7KjL+3GFD8XXveO4eexQLpznNd6GkjTCVeSk3S+eMLG1fhSgb7lEutVDKMYB+Apr2G28f/zZylB
9ikYf8bVWP3pKZR8lZ2t1oEb2A/8IO6fTXF03Rl2MN4aEpoeZ7sEUaErktINOwkO25WwyLK4R+G8
zGqn+p0b7oBiIdRZC3Ds9G8bQ+sOLycEh2uyPJcRlzjLdi8j9RV0O34HQbU89AWLkRUdoQeupCSo
z90D8tCYnXYpHffYAFfdjMSGUz6HWY2d4VvnEnYJjBp5IKX7zv/yhYe1Hw3NobLxjNEYhrO0wauG
xLSJR68boalFsvgq7ETH+BtIyNJKPg2CI+Tfes3TuBc1b2oBS5u6swTUm5tb/Mdyixgq3LrfCxB1
ku029Lv+vLfAEd6hpBT7iL3UShSewzTpBE2fW1lejzl6OspYfkkzK+L4Q02L6hfi+SP9H5u1ZKEA
yU3nRkg3wsJvo+y58+aRUEWdFKqOJqWJ3if7jhG42q04FBi61JTqzROST8HZFAR7dWv+C13Q3tGG
9a1Yki3W/ZgzeB5bHSeMnn9n1amtNwVEY/5orf85IjIrR6GhGEmHu7bgU8TGXvaXYFHV4zWKYnrU
rFOhVarapd8a+GfAfVVXeqPq8fh7X9caP/DGiLG4mJyXS0+e6A2aH2z+5oM8Fo9ClYeb1Ps8Z0r0
grUYwF2M2zQDBoWyDq2s7rq74I/+YHnizONsPLqqsNm19+eo0cbx6IGz23nVYt2nS9SiSWmh5tbG
/IraS81elhDSPuEuVnn7BkMfLibRdBmt0gFi/G79T/TGFdzTgvff2vrGji1G9b+tTANGlTB8vU0i
laUqpMAxjAnKQ7SZcgk4RRYouep8IcJZ7smQyrgghNHHN9FHbQdyYxbroV9QrF/8lInhsIPEBt67
W5HAlmN4df9QYwUOf/79W/PmI65MBSm0vXCDh7sPLJJetiDQz2tGg1Lh1vl+PHdbqu4rEJa9o1Nt
sH1J0GDlb9LPqkJswRJl/63MUUsS/nX7bTbGZrTksmI8WFH8uEKSypJvIUdJqKheGP6h7KGPcqZJ
HibtGtTZDEHw+XnKHnvfCOnxJ/5/92Vc2KN6YZJQwgOMzLmtkR8/2vrVhydahBxtxO3L/P0XYXgc
RZ3Pcd4uynkMexoAAMpxZOxSUMy+isCesGPrKNoHwnQQjUwXaFie6TM1jtQtGyZnj89opUXHOnoJ
szMQ3S7Mfd5nafu2a0LFaRbVqeWTQ8lSXl4e7CiQnSrPGU4ja1NOOLlxLdx5sy/NcB6v0D9IxI0r
wcPPDUk/IPfwoPrNjnDvdESVt4YSbn3P5dVyTvA5WbJc1FKOHhfPX4CXjmoJ55ipOY15CXp1hCKN
gl175JuGYa3ejKYblKyusgB8hxrGqrDZ9YjF6D4VKxFdlvAH7/eEpXWgjzQ8P7XIW2TG+Ov19irJ
7M/P66OvKm5pb/v8qAaB03EcVqvkNdJfTzAHauGWf2gpemn9yg6aQodrdtjPKlmkxZgnOBMvybN1
xVz+UDwIw0w+7C/nVHNJtL3/Kjs3b1s7/LMHXWnF5sAlE5kC+3mWLclRG7IjJBtIIF3aRHQn/XLp
1l30kgcaWmRrMt8u229LID3gIqDIFwJ0YP4xqIuZlU/x9gDO1hSq3l5MAl6CMB0cqPQivueKjNLY
oAMaamVPFhtnE5/aZ2m9Hf7gh//MWwJ9+owzn654JxoD4X/Y7LRs9gcZsQhhA9kH3ROYIoQd6OPI
Ed0bcKgxpWbA7HMnGFmCc1khDdcJ5GalUT6Dj99KwEJy1shzL/Yc3/KzeKe630wtQRCbZluRlykd
JXeGRtyAE62f0olq86Xi8PN0i/dPMxyXRsCCQLNlP40LcCKqEQqi7Op1Cdi3u2c0k8k4G5NNTkyu
a6J7TrwUUfOqR21nsNP1lTVJJvjH/o4PBrzlIh4qnGF0wFbRowUHxljuPKBuPAdwf3kpf1ek7iOE
oxob442P/qxeB4rfBccg5cWcp0F9fUiYOTCihiQU2Atou9IaHB6gT4owbj25shB3Kx4M0yH38i5F
6iwiu1teBJr7p2JdlSf9Oc/69pN1Z66PEIfLy+0oOv0L+9orc3FmUzglcJgKnIee+22Gb3tiMeVQ
57I8UUhGEwuckSOZWxILGJfAkSrqPChGZZwV3Gl+hHY2jtjPl+TQN4pCZqR0Lg1USqwhMRnc5cDk
SRXUmirlEQT6h1NfWvG7ok8cRAEUApBDXPh2Rdh2BIbwSb2cV02UfBbuUwYFF/o8Sn0H7rNHKAsK
q6p49+F880wo9v+V1AvaBmqEGbsK9uJKqgir629DQs3IPk9LwK7L9vBPAelm3uSSQYcwO51KYfwg
p4gHuS5MN6BWreUJx7OzmaWkWDaZ/tdP+u8Ew4P6UW7bAxnxyOhGLpeNT47USpKPMXgOss5YIlmC
v2F1xchsTR8y3wE3wBQdyz3cJRIiOYCoyOOW/l6fHND8T1vtNc0g4vdlYgtVdaLCbNmSAUy2cSZx
6YWZxnfB5/LZxByKJDXehgSWuZKtNKzXa1GZAgORYDyo+N5wmqNm/I1Cti7uf2WscgtM4buf9zh7
7qcp7hI0CFqgRoXZQ38STWIv9OFpPigkeegIZPtd1Flvy/3BLFaHztplm5Wm+4FYchDwQvpEFU7R
r8A5vMKBDYK/5QjtUG3r4UtMDRhpXQdIAdfIb4Rj0T/aZvubBf3KJAI0LjLUFEjqMTO+Cv1fy8qS
BMNqRjo7kx9qiKzNeHwljVFga5vGHLF3CdnLDvCdGSncCFmt3YYDMC4nuucg7wkcyLsqwZPcwktE
6zLOcObOoFHETNeIDrnmxxzqzzFa4kIIJBpH03Bz5DuR7SKUL8QA5uN6H62BImvlIiNQsWOKQH3G
rB+159GZzZ69/6a75ks8A4j+jKZJ7bhwHgVhShfj9Bc9F5JEigR+dyvHoBhUspJePxKgIEYKNk1f
40rRPTxs7/nNPmZ41F9AQ2cA+aamqdZAbT/gkLOJTuaEHT6zzb17JAMq340o3lr6jWn78wFvU0lW
9XmPXL8LpJNd2LiFwrUx4z92VHOtInN/23YAMwGUFr92EXuK8dKnEvJeqDS+4G6tWTQb+H7acVVK
E/wnOs/B0DQSXcM6cu6Q+xtHf/xB+6dgqM195sR1E9t1BuKoORSZWklxdT4ZI66yqhQ20e8s9AqF
9/kNQwOGx0WQH2JUobGZ2xxvG0MXLFslf00pj2XHGlBftiCIhYjLv2K/SXb5IBRp8u7FZuVPWJh3
qyj5zNLfMg6npyAj3VEpGGxNnxo3YiKM1zhZryXPCRyXSfeThf++WsXRS50s3zvFtly6iZ0epO+p
JV0dIyHa8X+NM0HxQ1heOh9GELxu2scFUuMfaxYpp4rnRg1NmA6aPh9cPRC8paCOTNGr0chDSq/I
xKDyg45ocLhamXc9Mma5eXwn/BZQtCF7Go/7Abb7b9SyhuSqZK22c8PSDU9ICH0X+QKduS5nuwFC
TBUZus6nXm11s8nF6WsrkFbwkC5KeCAbqe+BCTiQZjxE5ogzINjOdFBpygTFdER27o1GEnOHTMrG
mcxnGxiSdJ6maBwaCeN5IkIlhareamfB0RUGlMi1oYhNH/3TbbR8Ra9adcEn/l6Ktt36PaM9+KIR
uf1fyAi1RAyb1xGqt/01uIYfWf4EgUtA2mitnjVQ5cAQzqvFTxd+jRUVRIxo3FOJRHoBwlNeZsu+
+nxA2yXr/4tVvWh2tMgYypDWrYBlUGlx4NoAOhekZYYm360uGp0cz9eWPX7zqMK2u7mnxUzT70jO
hbD9/ecl6dHNLtygFKPEj7C433gvURb4EOgaWttx95PjHcO2YKr4mUMS3SQC+KYnQ1F56ZzSIzLt
5RNrvhqQ0M28sn0WtPsAujsbB1X8/k8YAbWZ+ANFlV3zhh6sukFNuLB3XLYqQ251RxNfsxUOFzK8
U8XONW0wEKyq76EdGgtMAbR6JQ9eIz9E6yXtw8xgUWf5wAkhkBd6eb5HH2tIgUdUMNHv2jnoLU46
uFFYOBGvYD8SR9DyY7I7opI/9AyEeCPoY1xI9L3OcsvUBuXVnWJWo4ljZTsDQSKFAd8uvoFIry2m
YhIdO6HpStlzrGEBShCRpM55qIARS1DNcTFEVAG0FU1r/u/3NWhTP8Be9LJLKzZvsIvuRPEeuxcg
+c8mC9RNK6ImVVg6fL2/KFRzZtZg7MxWG4zlAa3OiG3WjttMkf/BxOJklgawQPVKJK0PcTJVYfVw
fEwyrI2CC7BAhkolgX7IG96G6yDjtvLdhm2xjilUjjobjo8pugD6qBJDHoQNwxuFAIkyra9dpw5A
FhHMKFgkTrctaL0ltuJFjpVXcNXtEFoVok69rxWqozzdDSxXkPo2u71WxaEaXoLV7iay61P9sz2L
fEJVqE8TwXUO6NLQdp3+TiEJE1b8q43J1yF/jBoQxodroduaXREFbLrxHrn0avTARvupbDFdXgEU
kUmGebmjYkv4WBrAA6GVabJFejcYayeZAWFSPRBjvzWA03wXBiX/U5u9R1Ds7+L8NtCm8sZ2kq0G
Czydw6aOONz9mNDr6XHQv1TPqqfWDXOa7MWZj69+KGQhqRDxBfdxXwFfqS0icFG1eoVZ8f6zVJZT
f0igRcbOATyOdxk8tPlToCVSB2/ehAth+mw/b91UFbs93h4zN4oJXazdC9/VT189pMTvYoNDJn7E
2NlVhbnXqhZIZVGCGwbCg3ZEtkczD6WbLCATwaID9SkW1KAmbPrbCcw0rkfaVJper2f0GH52A6Ha
VQeJ3XaiVHg2R8eI1izNbglAnkEeWHp+C+WGS4M6Yk1HiCUH8Z6YhLiuikKsmJu/0+B4cQAmbsoW
+brMAfvUAwJLYaXf5NUBMFV7Yh4Q8I11DC37FFdT+bO4mHbb8Gx7pq8Z6dy1xSfxlgEwpt0HhmwH
3erukvNlGvFhuo+njRVThmsxV/lzBEzSmJ/3a01htCELqe/qEp6j0p40Py/YJr8ZGoeEyYWaBGD3
bWwFoSzVEVOfSvi0/Jcf2w7t87RrxdziNZAwfkTi9f2Tl3ra/FdK/GBrwkG8P0b4vzAtfwi7bB8Q
oLzjTTl96n9GRsYeG5yZrmFb/37iXEvakDXQ4tmi7HkLa7jBQPexcPar0t+gDWQBL+Gq2yTBMdUS
1cr9JbokwPNfKOf6HQkhqhtEAkbvCjIumHyDTQrn9heiy/JtqKVBpolDarO1LpuRhTTJj+UdVXro
2v1/4b/lLnP8TEGnpUVRNE76PkkPVlXKPXskNJcL2kA+vUIlmQibWErqi85rxAWRbjV05IxCcN/L
0REj4k2w6b4P11cRIiIvlBQkAn+ALqAtv7BJe0byo5YWl6YlLIrzWrQ80+Q4gjBRcpye0eqkidZi
6NAPvoXoUw+BqOyRMeuKnfcjTqVmWZlDqCG/sPPZg1EqR7DhZ2Ce0DhqvrN6htxldVvSKCMgJEjx
Ol9Q948qcJsBBKWQ5eZtMQofrIK5jbCcEfirG5mo9qdZZcH4Yjr3b3kT2i/tqILusX2n6bLir0mR
fZ/+UpG+/Z/VFaJqELQl5E9csHWYHkrPiw4AY4hz0FgToF9wzs2orv6r00ZunU4tBSX3SAvyGjWs
RFzJfcM6ZAV1ciRL2iUGjfden44BOPX7Yijc28Tsy7Q6Gas3HcKMDSPf5zb1DYQDSLoNZ9BkG49M
3Ezq5mPLogEImcRDWULXvGObuYZU5c1kdL7yHQaEsKWbAS1fqf6obzAQmCWlWsF2iC4RBHJyaFbV
lpEE9H0LQev2xt5zSCk7BPGjcFY1J+4VW+Av9tUCtmHFhAI7tdbBjvMuKzqkgR3mlsH3dgDG6vqo
pn6jcCsjtAIK68qU5GS6WfW2ui5SfMfueFfVG5MeUFXtANTcKJY006Ga9qg3zFmuxclhGPkvjPZh
eGbPXilkVYyEgxResFInB1Fx23sSZWNpd6yI1ytkBgMNPVzvX6ZviaWSYkVdQHLE4NQ0fBSrVg8r
1nz1+GNlcs3sHe4PF2jzUMh9b9dXTLailZSD6fu/Bjj+o+mO611fn+AGPctIfuJ4Ha939abWs9TZ
IRLO/dgXGjg4YRpw7P+TG5NeQujwhLiFyBiZh0g6DM/bpQlC/NQFuaJPa7DfduC1isxw2NTbuG0S
s4sni3AyZVpNjcYGgJBmJWIr5sZn1NJzVU4vy/FXYVEyCFSRh77oU2LE+hqrr6H/LgeWwsOAlHrZ
CpkIwTb4S2JlFK3HDG1GpW4p9KlAx0Ysi7MKgZRUTyQKfcE28b7okQw4ILOfEJ6duV+CNZQHhdYj
1H6OtEuSKYd8CobREdJWzHZcilzGg6s6wr8fqYTodXCDUK+PK3wvd+wfwFeZNMhXrGCjnZioRyxy
mXLGeYoOITZUYlfLIW+t32YzUR2JLxcaX9OX82XUvMVtbLVBnT+LfOK+aAnSYMh7LQEHAuRfAd3m
AH3xysnn66P7YQGgFRoJMDyWvbTOdU86EGg3BHwLGIOsr5Uv5J0loci/Bl7o1MYg/csc+8kLX/Io
Q8jfwtorvtA0mOjFfF9x4gAZjooSbpVkyPp7CwN46f7RUn1RYl6ymG7WCWP3wXQ1jakKO1R6qMZ0
Uo3NnlMHQAteI3OSX7zwlHuHetNPY9VaoDCa0jMMZOqKbIKTc6SvYEharM26Pijm1Mgh7mEnX5qg
coKBQa2CqjeYLhAE99HjPx68mceGC+ritdzKp1Bf/snTuys+IwjsP9O7Kr7e3XNikSwNx9p6skC4
j25EMMt0lW3czByQu/itpoUF9JVkc3/MH+Rkjn4raknAcJjoXBlKMT+yrr5z8YRd82cIFUMQd3sg
awDTP3Mp1j147sODOZu7lOhQa8BiXlkOWTIgSbkedSWrYdleBlf0vi+5r0trqB52aJOEz8jnRftH
vFZIkAZT3ThVD38acc4euXE9jJMoTo987XJq1z15jFOgpQQVd0Om2pQjESJiyt02LzqKU/TRs4dZ
1qps0KsU9UEIYmmjd3LjPea5qTnlg3G5OcRNIpclVVeqmiod0N/RlVWVK88Svx4wlJtFcqSiqFnh
v1q2ZoW9SwhWO0JOCumhH8oK0DG7f2zrL/BEphoxeqsw3E5PdPegqxmfK5EGGE2zQ4/dgiX+NLTp
kY1hOhuRKqTEQQpGqF9C5+BVi86uBTbks4bpYP3/Rk0d4P8CwBYg7/fWp4dZR5m0Ft570mEe7I7Y
mJnAztJfsdF2oBUIbx16OYCg/qHKQwbs/J39l2ybQGxVHq1P/Bi18XamOtGzzl8dAmMiTGDW92YC
7bmsWNv+K+ks7JOJpP5kDw9P/UA1c5Q6Xe1fxv/vu4utWwBMTA1LnvDdMcsdolaRoUCNli2jRGw9
JMnYqieoWEOxsFvzC17u83dAWGi8DpUjgUfhogbfHeKo0waIKyLWSgVQr2L2ibUKZYTc0D2k+q40
CqNWTEZ+0gx5eu1S8mvg6XxV/WDJsTA8CVKRGa1mDygch6gJDfVfQFZHp1z8ERI7KCkydd22y3P3
FwYro+XhEsYSvizBZ2055KbfzrhuIsK3WB9JfbM6K1B5jzHWvsLhqJaavWOhi6iT1xkWosrNE8ur
QuW7POSxIV4tljG+RQx41uMnYk2TzouzeV/JN2m73Q4c8YgXVxbnF/ljwl1pkQLFK30iYpjYhcN+
U+VK8xKQySodefZDHUgdUycWbA6+cJOnQVOLaXxVxzQue/T+KyBLxZoLssWjAqV+w+0Zhpu8NLpw
jm5rlcBI3nO7ETTLSn6lPpyP9H1msqNE6tUhh5qhmkHCsDxOzPLVJd/poC2V6dmFKJ+3662IJdap
IUov/UX82+55IqiHY4J6i7piV61GOqoDZbrhjPYeL62GDe9oHa0uBKcmAH1uD+fi/VNnKPNFUVqo
zuNDz5CSpDJyRtHzcUihP2EPF2JZj74j5Wp9bR3B4C78gX3wbu8h3gkEXfxZxC/ZROMOVif/2MmT
qrilqEC9+Kt44LhwsdRTKGO8YHfMcHfIHMl3l8CtwZRM/W9kxjqKvprFyFnmltYcW7fzbz0wvq2T
GznHAVKO66xzEdP44br8f9l9N8hlDT+H6nYFG44O8z0bGO2Hi0Mi+3yxYPI5kt4Zk/SV1Ydd/I2Y
c50CXBH/IGRtAqZw1ugHpM3Xkj51ZOz6/gu87sduljnmpq8W2WQNPjEya++Bc2Ul551LLChHl7mK
bo/7KqDuILQpzcRXzU0jUaHRYNASpQJauIc319FIPVEDYNQh/f8rZydORL0cV41Z6JlDrRqQZSYi
hpHRylObXPnqboojQvVvqBl8xyVA52rnw2EJ4rmk3t5LkMuwJoL4AUdr6a9bF4wE8xm0APj6Vv1u
W4mRt+rlWyT7hpy7JxROQOZCf8n4PVTI8E3+Ueoj7ke1u0NaGOFwdf5LNztIdJwj6JIYWlNeXkvU
XdbGqMa0Eu0UknBBUmGaYT4xL6Bzw/O+Fln9xacCrQoLwraO9LINGtl4q80AewWQiLkVHxBPoqb2
7DAIWOLTsU3h0sB0nW8UbMF9lQvc8iCLFtscvtxDYCxNHcrnQ6OSBYTo/hri2XpbS+BmKlBQh5VZ
pc4/1eSzas1LmK3FNBBRb0JJrFUR2cHY58/Hh2vcpkfwwFz+Q6CdoQk0BvAAxCC9j2l7pAs+8nbX
sfDPFv2i0rtJjhoxSSiWkbvtUwK8NX+XPUJReDkxciKaiZ90N2JWE0j8nFXVOoA+uSk6lj3L7PU8
Ttoo4r8QRxy4bPiVedO38Uy+ADm56V7ejV8DMupHfpU3w8Km0wfeZucXX0pgywdfz0wL8x3G3H2s
MT9jNjxfMHQhaqH7syT/EnSL2xIbysRNtej7njr/jaUTUte4P56FCuTpqAisGjSpluXogi/4wmPI
/1u6bm1Z6pIrB4IhbMDFwZj8dL7Sl48ZjdBAagH/Tlp/Z1i95jjqcQbV7DdxPB28VD0vot70SEMM
XyD4N5iG5Clrp/vd2Krs8IaHCFeB5Ghm5vKU/rXI86l3cQsCVoNBluvTZpun4CN9pofu9dJssa3K
ik+oMJL8dTYdUCnhSFe0Ng/4eO4Id+Zgygs5O0NFHTTvrI/9xrbU2mcMZccdctIyDF9inFaGRfUd
yVoUXS8fKACYv93wYVT/8HIREftgjCIBZ6iRt+pZnCWeoGuMPOT5uM5XrZ5Cq3fOrVX3NquQRTBY
1Cjbww/nDxATRdCq2CcVLnO130UM64KUD9s4eg6LLtkFOWkFtseQ3gkJgyvvK50qET68tONwrCEa
qpqT3wAWiO0QG10/k8MlLGDWB6ZAPVt/CW7gFQGSfKsNirikoeMozpEJ3NThgJn6NizEvR4T3xkm
8QypjhXq+YL4XxvaPZQoyomvALhxjhvwlKsWzMO4a/D9L2zse60ZctzG2g+dugv1P7AX96xX3yyk
S1po4QwDMfoWuNcKCKWzrk+/Yy2f3GLtNfyjr837X2lrF2dndakPQMMzssdzD58pzRlmX0wYOEfR
sGiiVLTJbe8mgnk6OX96ZwCp72/5WvLBYqMvOuM0BclWVL9fERNFtRPFv/6E5d8RtqZxpf//pFzd
sUX0ml1tChr08ohymH9gFFfLTsKDECyjfnbk79eHRDaQfykWAFloYTs7uqURBRbxf1rKNqbxcmyy
mvTMrtg2/HA0gDSNkB3pXZyi99rvFuMaqucguwPNJP9a/4OJGRihCDZAznfo9j+FPZBB+U6VbIFy
f5fMTCYvNR3kjzkJE3yuG9NfjrlWnNoLSZ4Q6usZ71EV3O+AIS71T0BKRZsAeMHvpoJ/anw05GpJ
pM3BajS7kTGiO3mk4gT+tBbXvwZ/crq5NbTAgP5fpZnGNw26VZU35cGQ5wpzteAzxEz28jcaeal9
gJbl2SoG3TvH0gJ/rf/tj9FFbtkxbZROQWuTdkeI/JPpqUSFcNhbK8HLIvwlOBNwpGqxqMh+Hp1K
IKKX+FAetYvsPEiACbnF4b6xmG0ozm5Q84knXBitTk+he/rtnh1tOrdjmMUsWRMuJzYAqB2wkpU3
c28fWPn2jULL9YVLDalF99cqz6CAPanVfHOS4H9LMmkfDsCRHjcOJ1uOv6j/+khyllMMj0wWC9nX
rSlfpuHkfXvQ+DCHtjF7IygL+9+tyoo4tJsnV/gxILBgztRfhAhlK44AOgc4dr2CI2sHqp6/+5s8
SqdvIZ5rLe4TK9d79RrA+Yt45UillQzh43jxp1PB6QTtwKbOvjAUMlUGxGdgLfaxAMCJuTiGBwBy
y65zC9c0ca9uQfUQdHnvvcmbU16ZQRtGuogK+gThI9mXGVuPJ/Ahkvu5p6Ql0T56oIKEi6OxEdGt
GzjWtmdPfrwikwVfgU9DbqX+IL42WtGLwT3dRQvyIy7ctKXnygEZl/PgHDucplqRKRER7IQj/PCS
uzwN1JTZG6B0SmjfYRfPkGruskvp+DgOenZpQZ8V+BcESqdyObJyK/l9Kj+KaXqB26wThpf7DJZj
KMhVxM6Ukx0nGILE3sNfP5DGzk5CKsFNcKq/yaeQWPemkJKHHVnt9g0HjkXSr+l71fmdw5UaTmBx
UhL0WIRpU+80ou6H1T2JpDD3w5bsJXRRXMi9pUzHt4sMjc1lhArgPDNYstRhWfoOVmD30F8am8JV
x9eM+QbftTQRizrK2J4YixPc19Z42W4Tg22fVPN14hz88/oS1F9h5aSIv+6tNo20Joyszytfi/Jz
s2hc9WIb+zZ7rcbEmlcDmgLIS6SV/9jjpIF4O0geaJbGfJDrP5Iod9CW0+XH/jP99s1DRtICMuxx
G5IPHP1noA4mWQjV4OnN06NK3ilwXlGrL9cEI74KJJNGVANwIfL9M8USrKdx1aonFi0dK8bjIz3y
ZgQhMVXpB2jNbwKN70dw8HjDGjV8zxWjN2BG7MXb476Kqg3Cc63wXSvELKzUfbqn7gVQTnemXDKT
UhnS8Ca23epuYK25HWxlu/cS0RVXcUFtUCpgZvUSX65x0mirggB7VihkMkG+wmMqBF6YYgEPyiiN
wGVlUNPEdxdfsUf6izNJ21uBYoVv7YFiwQK0RDPo/x4TsI9Tky7pTWkJhqOJ2W73ttEoAVQ7dTKR
5MZhOR/sbMNoLxq7i6m9UMMtJ5RXW2dTSl4R10JUE6btWHFJuXztR13+HFsFzE/LAE1WGH46kUCP
2WLOyoqJZWmM13919+qi9yashX4N8U7rBob8NezSGGNnGhFpu6Ii0dluZgA4cLquGTwEXFFJoik3
jML2CTkrjrRfYhocMKFQeckJK5Vd/Yx4yHHWNjHyeWL1KO/TknE/A7kxLcEnTLhaOjUzgyHnJC/E
dvwDrtXhNeS+rZYD76rFrSBE+NaxatlBWStuD4mHoXJiD/rqEKokGM0nrO2qRqvNx2aX0A5lRlJz
6eLH8WNydlPJIzXS/f5TjszK4jsHqAIQhuxh19ghqrCWBM9YXwV0SXuu1fAiYXu3JcpBlgdC8a4o
6WZfRJwtdG7K1wEGm57Gb37eIQ8+FA72P2ScmsTFfMvvmanqa0feFoKNuCxTzfPW+JhHC0XSL42r
RxUyBhr844tJNP+Cf10v49qeuWVFO6exWb3Pr3d/f82D552n/yhkF4LjlQyfbUERiv5d4DsYOkBx
SMzGpiK+u+MWxrSwB+OoWpD4Vmxi4n7JfJoECcAkNGNwvz1EOEGs/STyiPrCh9J3GNKXWy7v1deh
reByA0iqYLECFPtG4luJ6jaJpIf+NLvzDMH1brwNwh5/0+9xl3dRJHw+QQ+lYoL03ZpVWVtzbUrX
/2y0gRDEXiUDFDToY5Hh95gxHwCH//trMG2Q3XVtnQOBswiK5YIEqRzzb9zsIPY9tIemdxsI+T4o
ajoop+s/of7yjCSM3C1MRvJlheDFs/QblTzmmSVzvrsvRwX5NOCrjIhD8gFiUNaK+M78ifaevM/T
jc8J2lPIGJG8sncgLyAZpX8Yen8m8rZffZwCQH5z30Bp7VfYXJzlZvAYTv9Nhytk332/UjJTMU9z
rQFhV9S91rQ2V48rSLWmaWgGx4vIsSiHLqS4R1m304ebLT8iYyncYeauXvafEDFZ9wDlwf224Aa3
vreA8lfVagJEwAhQb+6ubYGkul4+QGtFtCdUbcabUk9ZuTtdUzWdeqsYnqn2CLYLvBEC4cz04OKR
j3opBMMmLD3tCk88SVYHFmUaNUkOtmH5kBqQGTTDUfQOAzAgl45nEBEONxokQyWEp1NDErm0sUTZ
fAovgGn1t2pn7dYGHTecB3eT5bVna9FxO1Gllum++pApLCYuvOsQNzbpmeqHwuIliCEHRhFwBY1G
kIF3GLfG8bwgm9DUfbr3P6AlbbqDJPRSz68dRTjpHZGhJHHdJ2kRAIb9HmahDMhv6dwDTzK0kp9w
TNINOmeLoIE43Fw4Y8NiR0P1V9upj768WtqtTExKAyJXYNrvK3Smfa7T0F6hGNsBkTLo1mIiURVd
aLGpKmgQlUMBgfkt4/J8g7CsemlMXFDNhx9lYw6p5wKbviA/it2JXh3Gp2sWpgTY75iwSvRAC3Tw
vAmp8mlklGbQducBqAipTYcHktt7kHxtyOCFPvz2BEuasNwppjeEuXZY7MMoVJAaKeQs/6gmBz2H
Y8xzkjoe6QCm+BsIEG93vMTadh31dQJzKyGb2XZORQ7LQbXOSMLj78fDsUZ3yquErseToVoWyBr6
5a7Exut4Zoy5OievFSPyPa2FbV0Rw69Iewoxvn6S5TuClBpYxohNB+w8oo1t0+RM1aEWRDglWA0t
lOTJob9BUIyy+oJWn4bdx+oIjjolSFyIxS//DtsTXy13Pd/+2J1A7Cur6KK+PipjIY/wwebntYTF
4Hr4vv446nL2tx0ZF8p+Lxrolnt1JpwFNgLvjIH9taUnNRDo4XqFzuRR7O3rDC3T0mzia9yJmwPN
1tZRVWIEHwJqQsBXEXRQKLJL3Xt6cF4jSNsBDsywx4aLBgE+psD2lCgJIXueJpWiYZgcyTffrObj
4KmJa7mtAfPXnFokz+w8fsOavsYPfhsO597VfrK1x6XZ8xSk/qt9xWoLAuvfR9N+r2jq+ykD52LG
BXWLPxPYEjQ2UZrfTsOQdOM/FYCfVm55BskWQXQxKNvnEZO+qRUiYApyceQWPpqB0yLPJfX57bl4
62Ii5eoge261VgBBk7bklNgmDdZBRQCaV9iWoTfJ6mcJf/X+mTCCp9y/njFFpbkDbUp2EkimLqdl
Oz0XKkOCqHoQiAXmZmprDC429RpSTSzNhve05BYO30WOg5bQcCC7l90owfcyYW8caySHQ+9A019P
nfLSXZrfy8ZQPDngUSgVZdfYNNNrlUepYXv4Q89PnsHPpiMU/laNZU2EkQpxx8QKggfhaofKgGdh
7O5cxUY0Y9XdGH9BWa7tKg67LNt7QVr281MqB0HoYYqkb8drNYwGHSZWMGPyFdmLWDQROk18vNMI
E+zrnHVbfYKC8PQStCJqobsMx42lFlGNbkXYtWteaO6t10EWQb0uZR2+Vx+XmQ8yxHhnvYC+3R91
1Mg9/vlwEUiBVnxaSh8d6KFeHiMNYSIPiKHzcUVLKVw9l30kFLlzzIO7sPajGNsdShKU2j1a7x/Y
YVtX3aj1xdE9TXHq9kWxg1QMa/kh/y0CI2mxh0G+X/4+FxO75SZftypoSc3aD/C5falBbl29l9p7
0fvckJ9DAuDWK6smjIuHjYaRl7tcdxK/lya0iKFOwtYd3abR+/BW7trC3eP9Y9IduMLDelIcFsok
Li4r/oz925ZftEtZ9knA+m4pfXbcOpq3xL3iB+ZdZmfJ0esxmzyuhwjtn63vY8cx5AkxkWXv2n0b
NBoKircran3E1KtMn72uRG9tB7CF4Wf+bZAqH2rdO+B3OoLq2HO695POf/Tsin5ASLQ2/eL0Ij/o
CunU3IMu+clluaurUPYiGUIHCFmcDXDyLI/1TxfR/nNE5SGqLbJJxfkeneAp1gdgsXQrPW36+gqC
mNQTMQFGjgawQWcIeHNjPUNamDwHByd6INdFTRJWEM+uBeRo6pFT+6HsgOZuvs9/S0fHZjqk4JBN
TQlusxGU0gVxB3S3C5gtsTh/+pcBeyNyFB+63FRSk6EWaWKjytE2hsG+9V+mEd5BdGYo6UI/k0hw
cLnYGnXdHTbscWQi5EH8haXi7ZkfJJD0ZPjNbu7zzKSGqDjJtVUvt2YwAc0lWgI64UEG9b5R8DdM
Pvg9y1l0kY2NwUfGMQIaxSf6hYyQaGFnVezy5rEGvhIqocmsaiMmEC/6tLh8rdVdu5pFSC7dbHMF
6lxNKI4W7FeNEZXQV+nWhcAXoifH+dJ3Oa1kheEAA1pt8R4KeKGar/PQ+t7lutQmSDrqZa6uVNeh
NelKJdc4v/7ambjmf0NSC/au+6reFRt3Rgygyk70WjD+09BwD6iKZcM40wwlB+PqTFPiMsXNAmxo
sW2xaehaEj0SzIC2qCT3FExz+KWoZUJx7HBZ7U7LacgOoM/OoWaGwKGWuPbLk+zt1OYnqawraTqG
lqr12XP8NGzDzskq3wpaN9r7iY6TtP5FzYaJoVlSL82RlSj4MmDQoJkjS/T3l2hA8A6fTV5Blbaz
tZVdjPKsAvsxE4e1gpBj7jJJSsG7rPta7CuaZ0cWFZ79zEaJu2CXSVE94WZTs/u9OzXAy8wxwAJZ
AGC0T7Re5FAtN4Pz8rsVV7nKkSI1MtLC+O/3r+yv0v596ZBhOZEtFChI3vTHFi0cauV3SnSIUFRk
2j1KEcMXjVp+pTy0rtspXsrap2+FF/We4eHouHSZwRBeblnScH6vNis2zqKEiD6g7ER2gCTDZIxO
bfvSOPFeZi2hYpb+CxFVuffZDa3ZjCTCu786AdpdRsVD7ztJQtz4E3iSNgsRsxDkBEv8nMi8Jvnc
cQsr0TulVBFyvI+hcNHnjB02i67qmyR3fg0nvwUm46K9mM7nbjZKQ4PmcQfuvFTgq1/J6AgQ9YrJ
bxyGJ+Ir1Z1r2QZbT5K7IelobcST1Dp3scFI7EvSPq0C3yjEFJD6taAagaRFZ8xHzaaRfLHiJDBK
4XW5QTda9SGPrzvO0egmqWLr/9rSRkXA50yjMCsCzG6GloCbLMdXn4MM8A5O61o4mGYGMIB5xvpO
Kn3Ryv6BHxeKuL+xS5d+iuYqbFumzg9KZR2eDoy3iaVSgE0aBMUmVALo2ARJy9E7R+c9rs6Q9d3i
pIGt3CuvPu4ufvrb1dJOmC7sHl38MmJ7zlxCLuDuX6+6oqZlpI2Q35c+6jClBwB+lcBxZzibZi1v
n+TpjdITI1JuUx3MUoQEoZ4emdIBnwakbDF2xOZAaB751mCaMGVcXJ+P631SN8+paA9GLZYw4FUU
Lx3v7tuKp6PnC/uFEwhid2C7OwjSEyzUroPrDbHwLGTF7CpY0lcWbqSSuKDFNjqo7RgOhgNB6MDe
FiRGK/NN+xP+Ccrw9kSStDackSqsfmI1hW5994XvbUT1CJtAwnxKx9FXCo2tnTWWliETxel2mjVA
BBwB+KUBz9kDbYZav2lMebBHfz6S+DgKZjLie/treAklyFkAT0E/gGos+JimUDHeRU20lnuA4a7a
wO+DGYXNjCnRChrDEKBhdt1z7G66sy47GUz37NIaVG8tF1QCNjvXThma9pmOucmlzOSVGVODnucR
h5dVmK6Nk1wCUH2/tmxQA5dNo61MVS3BFjy2ad2MLixi0fkcwG0fRXQPxvOyvrFmWEz7+K91ypeI
4CknjbUAwmng8VgmFjk7RnJflGt5LBYo6N5So7lTv5Ga3YVdTSrZMx1tmjhgb7iaAfz8+4XFTRxM
/wHpNDWmaxgg2zL/x6+EwFGLL21psggJHezllr+zPW7coES5VNyzsibZhLNyo3Rdte5ioDwrmGu0
bxTbu0++/2n0ZgS8w0hy245LRWIFE3wHpL9iZZ8upxAlwIKIJIWwiiDU1+QJj7YSNqKLSkyysJu1
8sGuQ1ma7A8sd0OsegbU1wPiO5P7vNMG4icc1f6Tr3J99giuvKIc0DqOe+aSOuZaZUzBpKA8zzHF
ThonObDpsPsW30ZIvFQDD35W7+gwZTFj477yDv/xdewxB2UKo85XFWOgoiYPFVTM9aQm+8Zw8Q3q
34Xtu9xqbKFppoiccTmqGiA1ptc8t481ZZRkHU5kRpPdvkTiPgIjuw6qQ87TT6JbV9jjrd+wTDfs
OGCzfv9O9j1phWYvySyPYiWJeeiEy4m3KqcXx49s3Mm35MlmrKnWEc/5LzewGl0hglxLWs2ObGZm
rOM+OCM6lAucqRHWYPVaarlAiwgNJi/1qwqWolcCn5wIeHpqaaoxBmfmrP4qiMOKUANMkHZXKzv6
OQrc4WYaI8+0G/WAkbsd/YUXvo5GxaXVUfCrjU7G3ulcZqxQlllqwjB1jwcQ7OeIM3CUMYqKcMqM
urcAimQMMROW+7jNZa3or7MrcxIxibsusYhwv2yPI8rvFJ5oksVRa1SeIpE9amqXwMzgTbLgWJJ5
1vfMC2Lpdrqyxu9eHoWWdC3GoKtW7zjnn+wnIbuyad9pxtWRN1JNgwF1eCupEigrYm4sTBU1kzRQ
b2ZVVW9z7M+uFC40Jdibk2MVdDMTug9Q05Xe1B+JPTm5ty6gDYIxuc3Jvdihxm+cSGFZcymErr1i
5PyX1mgyreOXGPAoTGSRZhX7L1U15TzONYLqe2GQrC2EQcivTNEz9BP+9el8hA52ihQT49z/xLKC
OIqUcy4r/9Q8/MkppVMXrrE1z9c7uUqPO7q3Y3DsBcTub4zGlG8Z9mtH3vO+F2lq0UxDrBYyIWNm
WMrHU3m0KW/Y+61+R7KNZ9xj6vplJDMVPWTuXsYeQFDhA9LkgZw3DHgKCzrWVylxYHePwJreXjxX
rARA5r0r/m5KJWJPG3H3SeH4NHOQStPZcSysF2KRTgY7Yi/lvWDvutU7ES04s6omMSAjSEYDWP+e
05/E86CyhdzL420Ibm8gbANIEliET8gNir7WKdVUL6O2wZL8n1QfUf41DiTdqBnDQi4SCzHrMqL4
ymnS9234SPxzcPpQrDQedAjM10BDy6YAoYRsqEHqkd4ynRAHPiUn1UZkvaQvawIFbRFDCPRixiwC
wCILMyypsuwCNtwo6KDmHvAoZq2blKKUD/g6jSA5XmNTtD5qVuuISiwCiBGECB5xv3V7MrlmKUXN
qUZ0Edw8T0DEPDXIO+iGh0Y7M3xVcq6vESQ9YzWe5Pfo70Frn2CDBvSxveFdxWpkndeJjg2q4oBJ
Yxb33CSnJBBUDUuDxD+wnljdl0eujphpbUAjEhEP2WG9IabbZC9Zl8zvs28Xz5ANGzfuN66h0Xde
E8JoONNNR1OJ+9hjkwd72Qz120iXVoRzWc3kblXylgbrEusIuHE6Cicp/YBtapIIk3R6opoqZCaK
9Z0N80X3zbrYbwWGM34uvdHM1vopaPDeJfFdclJZSS1ASzdQSm/q+gf26lrw3dKJdKVsuFjF58Ny
fqBaWxeUdhuUN//ANsV01PT+fvoBwpk6lWsx/hACdp3Z8UgnAnvokI/5IhNWsfdBZnc+JZvPJt14
Mr9Arataq1WSa7abECYtVPmFOC6ZMxDAB1e1ihtpVpIB2K4323hMNo4JqHrDtjsX89xYfUOQC8xW
Io1a4Bnb06xhb5TdGZbu9k72BNnLYmO39EtS1FOp9tb3T8eLI4S0dLq+WIBWmtOEyn2VqAkZ/3M7
ilxBUr4EPPU2N5Bb5CZtJWEi21h6lG3OvTIsnRlKMGiOi4odFfUrORLn6/Auy5quw90X7q084COG
kfsqe1l4VavOcgCw9QQYPVybV4JPz27O9jqYLE/pEYMY54tVWchYCQdfcsym5iY07D4j15aSCQLe
Z5j8/6eFkZFiuyoXXjza3/vqCl48v5pgT+QZUTL3TbUFOklg3tV0FoLsQo/vsRB8b6Ska5jTVdea
+HMwpYNtbCnjiNIu2xGmWDDilCrKibhr7RJAtMzJdb0tyZ3F9zZuwDVbH84ltSJBPouRdsn8i8Pv
TYc1Wj1HDVZRxSIn8w0t49RgB4BhelbSIp/C/qkuqIiNWT5sydQkfImMlACSYyv3s9th9E7JaZFW
pDeR4maQi0aAqOas39xdiYzi6Nh4AyDjcHQSoq49A98YBID0I5pEGN9RnSCLHuYX9O/tEQsHy7rG
JtvnUygkfreLGfAK26qRkIGX1tsWgJp0ckdInPEXSOQoDIMg2WiIPijN0V9m1yqDGt2l4GXnWRCg
XWq0MAjUfJOx13F/8VwuoJ6YKgLB1X5jUxuJyT5eASVdkAIecJLLfMoXsKjFg+ztNpwsJEcRF5Iu
082fYatmvUW+pRniKYcR4yoC23330cfCPmhpA9K1agKsqfDU2Dt//IlJ8y1s1+Ea0+E9w01DPX7A
j+tKj1kBb9MLLdMqkVcYqF9o61yYvbVDNurtdrGgazDjKW4t4StMlLViG3MJKRLAmj9iYWxbX3RO
roj2xXZF2aEPVVbGkEGUa4aOaw4nH4DI3C533hE1UucoXmNiwiRdkP7vP2Tw/9MY3ahq+MllJkho
kxkBXLs8B54yZxZipp2MyQP9y6PrOA/4zewzi8LDUoB9nNBylsHpHWcCChbFWxbC/mDeFxfPU2vW
9xyFZIl7gRFoz36YXzEm6+aFksMa3esBw9Ht3f/BMOyWVuCo56lM0LI8sELMMFiXyyOllBduwyDt
xxpnKXwJvagKa07H7fUWITBPpe7zYutbjUkgYuK4yFAdP+gKrCeyiyQWtPhWpIN5Cl61d3ZA/AhD
LplAsnud1e81Yc7fsE25HyfLF1c4dI6woA8rqMvaI5dsk2lBS/msV5Ur99aU91V1Elvs7j82LSZc
7gPbNLGFCqw7oD9oM87NCKjPsoH8dnRrvYHfDr0dhn/0X0ADoU5NDwc5OxsV2JCR730KgBoW7SFx
EDnAGa/wjKxUyyIB3ei+TEcmn1RcOZ1Iu2L50jUUVFgMbx3nZ5ffUW1U2fAMbNPtwGaHRWtckwxJ
7rmLeENLQMOfFFhfOMGkz+WqsX4Qx1MSodjw6tCVA6edER23qoA0mzgJVOiLOoc9zPV7hJlbEJ6p
vpgWkzYGTpBEY1JKKlY3FIpu7JZ5pd/Lv+A+ItM+LPmlkMFexomSqe0oQs1CGICAiWa/UGldWSSm
8emPWtLqWIe4PdIIhmchI8R4mTjeepdX8ONuvdtHjzHWbnaEjcuAPN0hYIBJS+z+xO9EpLz2ZdUJ
qJAJtUAK2hdVVd+gF+PamPNuMx+vnluE7RsFTgCuudcHLlub9NPveLyZQNzd1I2X5hjIyxfBbxxM
VU3aFMLx5nT9aCCHr3avdqPr05kOp+CuK2O8HzA+XyKV2ADB7gMRmCOuGpmG4fPD/pN9fHZ7h2du
xLLYMAOQaT64fJ3zCbqhFxfqjoVhYge1HJr0RLQJctqRGrcBArzIDy4ucFsHIDbJGBTDPGfeDbaS
Es8+l4/rvXOalARQQ1occ34IITm1HG3h+RhQYf63DP242+bmtP1F5vkioms8zt8zmg251aAR6XdR
p5xYcjq+4wBmfOYoo3F5oZRQi/7YM3l0Eml5oYSOjSrgsxMk4igTeB4apGwCEi+lhQDfcmEavBYE
QWAxPalfRMUyXQqVVVj9eMGtmlCxqrSaoyo/vsCi30VpTJtN288wjQ3/MKbJlb6nR7ZD42Zz5PvG
EWhmSNvKI0qOvsxrb5xIZxYzpuAKXUojaf4YKCyogpnS8943PLzl9BboK3V4gs47XQQtfTj/TVWQ
eS1TypnEmRCE8BOaBzkkHKI2+3kfU6mjyLXWWQf5Y1LuIejROop4xiAEObo7Wz/ke5BYvDkJgFpS
xHXDx4pWSFk+Tab3Sd14Vmg9Wt1CI6mqDYpDg/DS76iJPCyLp5BWhItVP3oUDHcRiI1l+mFuYneQ
RDgN57PVVlTVnjRaUqufn94ygv8POVY+rf+/YqYTusnu+UTWja2CmIS05m7A3iqCOX3Gm20sMe92
JPfByMLmn9Vmr+E+ELl2lYn4TJs7hmmK8AwC3ZojtSHl/aezJiV6wW7qsRa6KlPuBuO7B1DCbP0I
BbgCFtuT8lfmUgFIDJHAJZnjjFUtayLOefUHfQR4nGyxtA5pQoe6EQY3yhtWTJLJfHMtcgYnyUtb
B5byz50G6K2HxoFrinnbxRizUIPSKUlXklFCjWJsoJai4nciE5nSPu5J7f25odpeZF36aFzMlOFs
dZQrZIoujqsgOd+xLPcprxERmQN/MiqwEmJtc4nuNHGVZ4Ngr9JYv4X74oX5Q75wyGJzk6aKg6Zq
/EdtwdXEziVqfzP1JfEmoUqMSikrCCXoVFasoDmVx/+dsLHZg3ecVcpue6XVptIfnppSWCH/TQHD
q+gevCj2XuWmpwdw+dTemfPaB4wTh9lU6QVy6U25UyT4s/4QYBYEfueS2BbnApQYTttWGUVoHiot
GyEkF6dwD2mlHo9nMJiusvTDUyVPS5uMjtAVK36envajcU8tHcy2x1CWopmLBBPWeyT3PC5KMoyC
Z22WI0OO6eYLNK9qrwIkolMwsAbXRMXliDdaRaA1SyqJq7AP4jvapMX/56TTMduZFGgy+PB9gAt8
E+vtqzTDlj76frdx8Jz8NEXl9wNUcLIXZsP/7z+5VI8scH2HnWiWxP2iIhhMddTdVMM1qM9qS5Vc
i/zLfx/zrq8VMZOHDz411V7QzGGUEyZarkXUxYx6YoZbjeik8Iv7LJc753c3FxK9NSBb8h8ESSSJ
LRMSN0tTPqmFOODVzo2SUOhRTUYlv7bO+rWltwI7f6Hsmnd/tJOk8XWwwLVSfHSEqBijuH1Cv4WQ
xB1v8GmihIIaumslmKrhI4lLmw3VEEJAqWKssL1yoYANrCpcex55PBUxQfB511ICuSkWxgFhiY/f
VkTZL/36eM4L1ZasJhLrWbd1+ImtNgLr45oOz5kk50gFs5458UQ67X2OZ9ZJ4D25BbQ/ZpX/utan
p+f6bss3cB+ilT5NnKxHfNNUBbUHfP5wsKMazcgCR3zcVWaiTlJ+hIatlhMkIJKP2BhzBjeyyDZN
8/u9rys8F+KNl+qaYC26p2pCN2Ab1LCkssb/Syb+JOmFahA62WtopUlOKlgL2CCcKcrOsW0Wd8PG
FYxZYL/2VgUkCW1nPVlQmfhhIoQv3BE6Km4p95Wabs2soRbaTQq1FBFgJ30h95qrYrQijxbpfTHC
1iV9tap9q0BdpfgoOHGE6TOgj7FW973e6U9FchSD3ODkg/sALZ/+mGwL0B/9mw94aui3jtkbWj5X
60Zgxny4xpMXksJvnkfy10mQT2qzgOzGuRmEj/DkYxqg93hJnZ2tDo6rpZduLx9d6OnRrjjMdbbE
jzPb/mE2VwQ6/onXloMLit25Pyi72S2HlTcgCxZ5JnB6SFyrnWVcpNiHxKB6rMYLSowwrkM2M9+O
YSMYYSlVgwmMXF3RgEqrQWbP2Mu1w5CwhZrdlT86ytmUko/ciyXf9c66RQzpu/Gowezsq62NjWk+
iqkI2RTv3gIEDf/IrSqt/csCS4qMhdrqmB4CVS6ievaMKpZhw4SIf3i1of29ZqrOSCFmeSbrjfUq
M/69FERwBqbISrHPv+XvR1TicXg592pUEVz8UrTxwuGytS2gURJH2uQU16QCOrMc4vgG/dZmKmQn
keKNetJrKFH55e5ZnvGLngjbIHZKBOQp+pxNbGFzfeesSvtTKOUrh7a6AlRT3xqJW/I+UfyvQb8P
s7FFEoy7eL/MpLFT+Z6bqyIyTKPYTMTVuKLqpO3pg+4gpzcK1E7n+HQ+vuX2xLTrk5Lmur8jfUQ0
yjXUqauNmWcOv/eeOhK7JZVZWfA+2bIXadO2AokIJdU8W0Cuf4KP2wIDuhqyk3bOl6PUL0JJKNnb
r5mLjEFMzGFcqGAlARGRS+N0DCUlMplge8xf4JlP/Ywd5OIRbRB0Qxt/F0AfvN7jmlFaDvj9YHjM
c5Z0PWyZbb2SOBmLSyqk4yqU3BfSdpC8UZ8r1iaXui+tJxcnEOVyqD3Gpwj40S+tt6+7y5OUrZV9
N7u9HZk4z3HUx5NeFSpa7++anDTaprOY5Fg+ag38yGJlQZrrwc0bJxH1gfBuxR4ZEMaeQiU27Xdy
lgni0NmuQKQa9MbcMHM0m7y5lp2KvOS+MESICfQl7Gse5AwleAbOZ4usZz+EuLdGdWFFVAUyvCWJ
LyCNV5xWYPS9l6jfisg/GWSnMteWqPDCDYMxiT52rGZeqqVUbGpXfQ6RyjOTeMNqUR7xzvaktuAy
kZZNYVNPOzADsIF/vqXLUje8XavMbkGPbpKZd+9gg9fBsjzmDNEn2X+l/0R3iOQeG55I+W2jDYI2
0pX9YGZdWvk8t4COvT8kNITIHq2atKN1JOoJBDc+fofoYKtoDuFlo86FAGdSzBOVhdNtOtykx737
DENO7jknWE9VLMiGaVCEKMt9OwOdns0HI2xCwg3JXuJ2bXnEEn/IcTs90dFWBzfvPJ0XCUfuefv+
PEk7NYYV2jZ8bb/05KJ8m80GV45p36rENM9n7xtwji4+vU0BjafIrQvzkgh3yDhOpY7+sN3A+nDW
wKLLZKCLtWCasRO1fKsRQVhiOSBtzBSQLjPI0VNZBgg+XK7s/dJBoZGySOPAMi4tIxJyHEY8fds1
mVgWbcAvkepBw5BW4HJ9RWop9q3CO7gTv5iLi9TEvVP/KYEiIDJn2XGEzyljRp+kckXyvxX0jrlA
wGW5airte5LmW0SZnqmX84NoyQQhicl3PLe2ynBQf9HpK4z/m6NWge9KSiLe+GyLORXNkVgfobeK
qHEUyWhmyGEN3/wp+GgDWWtxB8kxw4gUejLikY2UZekmQP7ta161x2oyhwfrm16BFZsYSy9p3mTE
zvdMpMEGTTT7Gqlk12RT3GYjNZEI2hhMk7709oXEAudhZwoS3vRhHR3sAr9mOiSLITezdn7fqtyv
nUmIvORSi2Tpx/dThlTyEjO1VnzaE0tmAo9zNaZ0eeB93OkSDOPDsYbw5JhDgL3c6p2LuCqww0z4
tdL/miDZmnHC3S3jMA0bd3K0JbWYJKx1ohueIauUzXmqXzpmxmmt5Pmu0nO5/K+O5o0vZoe/UGfT
LEkFAByHoV+OyZFQlzAF0q0mVhD1c3g+tw7ny63P6mnzVajtQbHYgy7DsMPN4DiravoFyg6bt6Ag
mMnq3mhJrJP8NXjcuVCNAlR8la/Uun7EI3c6qOCVmoNBDnai8QTjhc5mtdbGnUe34tqMr8QL/Eg8
UxNQoQaJxGBAtAU4nhNKbNv6TvBdOMu8hL1aMfR7iZiMAAoMn4re6sbE0bNiDsN/KsK+xuD3eqRc
PMePS1saXs7+ZrvUU5Uk7f+kI9OYsA3V25zKMOf4XMLl/GF++0WC6+4IgNorgU3qUd08OAPCEm4c
BoD/rk+wy7nigyF0nHPC7thoOCc7iv0hG+eRkXjZZpAiICt8lfwWjDyzz4WQj61VpZXlepbxaqyl
QQibXuGqGL3M0kN3bYE2sMVCcDbqPiZgN313Ux2vIXk4RMmOH3SPJr9XedzBSfQ+/4IuRThBgp/5
W8FP1jvu968pYoHEFPbKJd2IqA8ehRMBA7ErFqZI8uYMPWa7jwvyR7ViqkN0L7Jpa3cA/d4NxrZD
v4qpfWExGxmYjUXlslf2PCprtCb4QE8k1aQlLAVpD3nuNJRksIXV1SaRzIvbfkXcLtf00Sl06BVr
A5jt/TiuV3BObU9dRNgp1JFhCjAUpMKRywrwTwnezgzIaFe4UVzAZc/UXsDDwdrZVQERggV50u+j
dj381rGAJfY2LaGPHH+ZUkPr67HoFyhbL5il0+Y6H6VfkdS05GfLfPQ7AvIiCI9NjxS55eg3ofIO
fC5TklgtSDoUBOHMVzzO2XKNkhQSxHxTVPuM3tSFaYzitnDt+LVHyGMdl9SGwUkN0a6rZd7/MMj1
hJ/y7p4ixRWBd4myrHlc+Qzz0pHHGV/hxUeLEjeF7V56FzvSLnJFYaVXaMp3suKMOJYEdIYjXZK8
HRrKdFuB49cgW3pOhuuilqMAVIn4BnHdBMjSf4cNpdS5L5Fjx0+uQl/pyi+3T3wdCDRCzaa/UP3p
8YToJDguuB47uF4j7f9NtjFAUCcrLpJwLkBF8wLi/224rRobXq/MrPmJ7vumqrIyxjvDfoBZmo2p
pS1yfh4aLfTXyx5dMA9EhSXHYcsIXWLoQTUKAqHW0LdKRH7DbSVuqR08NSGBw7SEjQxnRpkUWsz2
+bd0ijx1vhKJDB6QZYletqjY5/vm2vOPImpHztPycnVApH9Q/IXE/9y98ki/xL+itngJ4iBkw3Rc
sfsUBZbi4a8Ah/NmW/MD2oXtRfseL5tkkUAmTv4aTThuM0t5UiOXs6Dij4GUuI8PtUHFmP5L2cl5
DJw9pcxP2oZYde4Ej0RKNFtRTc0/OURDXA30vKM+BEYLZzGDp/lq+oTPUrjvnvYKTSVWb3PUVumD
vk4Bok4nkGIuzh4vuLN3Nt6Fy420UmiTdSkXnUUWR48A6FrsacmeEEFeZe6DAnbNTaoa0Tg8x9lp
nEniC8w/2vgYvnsubIj/OYj1t6jQciGz8ohAR3wQ4U43NrRPC8yUs1Vn168jJ0OIZDlOp44WFqwr
4nz/DnAipd7EfPSd4NcZaQUm6NZsvmP+pNdtKBF1tlpUqWk4KZW/XZVZ/Nh0YymO+4oHoEHRWJyX
9W6ZFdhtZpvQTEx5QPqnHw2pDvlCA3/qb3IeYgkcvmUJTxuq1ulkqcFEyS+I0hEvm/md59nbpTv9
wxoFZ+bVAAWWrVs0dXJo2TEzDiZGgQGmF1bmhjoM/7Bjky4f8EThc2ltr8iTOrjdJ23usbyIQo8i
h80fXd4pkoHzPrb67ZFCYiwipi7ZB3TZSbxhXCOTg0sZZxuw7aStemYYgmba+DKaiXU9SToKLAGt
P8t17Nd/aCsPzjI5g5kumTsHaNICDoo5KPpz4eKFpu4Elro47ju2tJYuqxFfIstb5/fghZBiqRdK
lT2XW1ZuJh5AyRXe2RYykFZkw0Nq6qXgSPdgdCtROrAa6skcy8oB/uCYBZOY1x8RPek60EARJdwc
6jDIbTNwaMqpZi0lUEAgcGfCHGQeMm3pi5FH1LxsdYazge5P/O5D6iF8MbYD8WvMpEG3k6Ltc8Qb
+F46iry7nPMCsr2skDVEodABLGgY5vthjOoTUGneK8vWTRpV7RFFTysFk5iJjeaI4PBOleCrk8UE
8C7GSV8fsJFymeYye9X/PSdsMdrBa05F4Z8QMuikxRi7NGFqd5RFq20aOCYtEE8s8YD4J+OApUk7
vIV9WgyE5VN/wulhuhaGhdaYs4cPk+z3i/TN/oWCmqwQaSwyxV5NPxKDi4ZjByGQASnXhpIxqfDi
yFLz/fo1GGaahJW3X8S0npHWVa4vpEB09r1uMAlWvMu6VjCmBS2dQO2uSC9SjhUVQTBtfGGtNaJE
TABPpd4oXs7RqveoBi0KGSPK9lfQkvVh87y0vwkE0HZi/hXz7yEHQamoCddYocrAFkQygEgokv7O
mNzbrmubC9QX2lQzNqvIZaDIHcht0wZyOxc9FfGiLj/61NDWDA4j88R2ZsLusHAp8fgtPW043Gth
7BN2PtS9UHwGKzpVVPoEnmqRSWUJ/z0TRcMufPzRAWHIdzQEaDYHY8EEZ/zjBT21d/p7+CezZ//9
T96ZZoMTP2Nb56mwGaArsjl0B29XG3H/XL9KqV8Vdkp9aoJsTMDz82q8nAK1IMOe3Z5Jb6Nnxyop
KYQP479AM3hCNHk2iZvbNQDFaVLyARknwDDK93A5RxTTbYnpUurLxZaT+h8A6JBp+c8/WgeuEBsJ
yenCvGXlsd0lacCmkbhl0nL+FQeGBwJDjdUfw5tXO+LiVwMaaE1H6crYItdC78HKsn6dZJy6Fi2q
2vNy9AQrSEeAWMuoFDAQPmfhk0vmJFBJ0gXoHp1/HgI/sxQJAa+nIxSWQUIdy/loqqvTN3QdwRyU
Gv1JvooexdhnQNEB9/Np6j2tI/h2BR75wIaC4UsvBYiBwsV14wyu4i6fVksSS+YruBxxysHDsxnv
kbKQGcHgU17GvqfhL2rOC0KQF60lr93o0CgmH/++RMRuUyf2ZTAprl+p+w1aa2IuckO8Vmx+QLFS
308w+gV8VDkcYwhf4a7Uze0Fhec7Nd7ZYffFqLJSkr2GuJzh335DaZ/e+NXc9mzvYrY0D+tadZil
EbEoFI+hA2yQ4GtE1uvwLhqN4U9gncWfiBATZGmNeJA2N1mMQiPPgX15P8+y3EDuMyW0de4wdXMY
tUOQ27idVnfkeLOupeju2DdSueAisLNoM1/eCs/KsSp8yVb1K2sqaQD/UPsdeQu2KazOK0ISQ8nT
JY1FSqunCnAU/gv3ecCGhI/TJrMe2q+ti2BbEu/cqTrHAL215zlIu0g4+1O6sLaovNSbG+ajcxt/
sBYjgbzlczBwbmwCjgBO7jWVvy2ZRxwuHfWWtDM4uqTmMzcSw5UU6ZGfQhLeOpQQFgSqlI41EBvO
xGxQtWz2tnC8IC+Kny4MdozRG2e8pQFetDqq1x6gGp9SqMZkkeoTr0X790tra8+zob/ntGARZsu/
g//kI9xc1u0iQI01FjxdZG36KS5DS0rs4xkZdNAEEFKt1LYiQJMMOayPYHej+vN40Dwi9QOuw9Jt
jGPyRiC1cdvyPlbIeXiYQnI7BwNxDaj3vUkwA09PTY86+HCKpbtpqH+NlOJgs+iiIZmzJcopNyA/
Cr4VJs2T5UhLglCW+9rZSabqexQ+TytUCWZwSG/4AxulkzpndTOFCOa+YRIa+C8Ldb8kNTsAHDH8
arfE7mK/0VLERL9DNdxgnN9i9fWbokzHPt/zjncH5JFx0LehskJFVxipAQPqTTnTJbiCkBR/gKzw
UjgO9+f2VJKkWNSb+seTF2PX9GDWUj88Y8GsYyyixKJLkgxnmCKAX2BSTx02i8G8zhwIfvKrMaC1
3s2+aZ3bd7FOAAtBwA/h32Aa0rMmKt+r1KtrMFAlKoBhYArTx3Uun3kzXcVHGLUZKeBN2roOGMI2
/QAQB1bMt5XOLv0OhDdJGpKOHBmzcwLDa2WPcoDbdoFDtnGE1Ofezqxrf8YPhs7nhUw6TA5PAlhj
r86aNva2ChHf/rVTN+xnt9Y/bdhk7qUYQLXVl4N1e5WJZydZZY5LOKbVakszuqw4d+3OeDRgHlee
Mn3RIlqAjETZpeRELchKesMQbsYWd8akDaSmrarfLoGl9Zumx2dKYLF9JJzeu5RVdf4zKtr6oI6p
p4GoWxC+VLZq5HWNjPqV1UCxE9k6QEjrRfX/C8aZe+gXZ8QcaD97EQCzbP2FYJNhVeV8su7COoYz
UDauTyUqZFL74JAYAXrZvQDmeKGO2PwjZtzIWgzrMEUS2kHGp9ODAkAOy0mNXHl1aaNY+wKLgTQk
HmfcubDYCRtio3zrQMvSbrOsQ5qN7XaIHKoH4qtewI264MDwH6XiIOKmxu1lePF/vW1UVCJKOq2j
wkjISPQYZbNiXI9Qms0iIvHmqFHFBOdy9icgubT3Y4QKiJkbeS41Hq9NXoPF8aMpTnCnTNJ6h5yZ
qq9JXXEbMd/Gw6ny5/iPwS0Ivr9tKfrSgVoiV7bvqqhK00j2jvUazc7Djm2PWHvzsqkD2+K7/ITc
vdBrtmycypqoEbYYRfOm2HuMHiOeO3zoPW8tsqBkTUQkEw3h/+aw8X0Ts02rJMLAZ7sWSsL7W/S3
n9ra2yCXefWYlEu8xr/eMsowyb7gAzzopyj6O32N9xvZW8aDjaCRfmw2lJzfHQ8x3ifHdun8Z3LQ
NBaq0a3jAmwUt/zr+Ta/ekJMvoRiEUDJMK0dDCYTdf4htC6SwzYk6gsxTaNrMQNI3pHmorJUAHpJ
ZLL/r0UXedxbuGYphUGl93j+T6hF7Lz3MnioFUyU8z1eFwEdIgUdO0vH2Oa8eEC2qnnCOMBblmBw
L7x4xjxHb+fgr1c2gxoAsuowc8swWVCat+CYKqc6+d7TuKSgp8AF8XUlyTGIOIGVgvmi3Ix8Pes7
RJTgazUpToxA6xjScK1yNQdlIntS0FDTWmf6vAbvhQYrXn6e+tVhw584xu+xezXJ9H6l8S3k3Lv8
ELwU9VGCSBxmAgzHc4GsfKb9pkimmhxVjm5PbAPCw9qs484cwNPfecKZ83HiXrhL+cfCtKz4QZdw
Uf0iP3IY7FMBHLpwbekec9KR7XYJHR/A+oe2stugOSMIvlvHRjzcJ1KQwhkidauyZidTfIA2ruoh
w/JZHq1X3cwzEs8eYOhD5FgvLMne1tVtevBCDCvnwxFE1NNqYHQZOT22o5AtiTUlctVWXU7U1KGz
CCL2uuikJV2BMBAgIVv7gMfHuA0N+A4a/aB6h3L7lyJ/QAagFGkpH93lUszAgZEvikUCI75eiEpW
RdCpIuUfmOAR2/XnJ5x7RFlZAtHOKzBhsOM2VgNdygOjAKRuPe1lPr1KTHcu8l1FHt9EJDz+LCy1
2rWJGeUbJVOplxMr1sPJhfMTv4UazVp9Qiwor2C3Dvfl/sXtfaRAiyjJmhMUP4v4J1TcIgoCKR+l
cNiOQaQnOxSbCbgTjXVMdVy1iHf8K0wSoSr2gHqBtWoCXfcC8xjzh8SpD5Cn41AnUodaSCJS4Y34
Ui6UkwofZvxN0lKC0Ev5GMZ108Ihb1xxr2+t/CPrSMq1Kj3ObpBRihc9ycO0wechkaHrgQqDDvQu
fpBVDSJgjXLhx2KIuyzY5rqcCo0XiTR5zWdwFEfrh3nqVy0qtGlL+3vFByaxjWWM3mXUh2zQEzCv
Dy2Iev2dBT+VWHjWvioj+ObSUgDlYFpfu4RmIz9Z+aHBMP5H83fqwrm6Od+t+/+0NWuW6oKgf1Hw
wAx3zw4vbQPK+onkXUrDhmWedOyq1iaVYhKSrr5qlRjZpU3RksKwR1iCYPy73K8JUI4QEFL2boBc
O4fIBKM5g1rhzvmjaWfkf4PENHsO0m37TCkfH8IBuJdGdquHVjDkjJUejazlUMILOlWcKTcy6j9f
DBKGexkfBDoUUdilOaSjtgFVD7lPsJEUMpfPGXLM0v+zaKGd6jTnH1zI63Cw+VDgBiBpWxhianxl
FoJFl/wrQO0heEi8cXfmd2EXtItFchWcHM+udwvpO2PY3NvSyI5wYAYfVILBXUuiNphDHL9WHHBk
w1L45KfVb7nvzrEgKsBbKaBUiB8jYyoI7i9t2QZXdPjJyiUAXFWrRSnUxai5uqt9/RiWjd6R5K9G
UyfpuUx4xJvkFHCYaMRqdlrObBty8kh26qbuElfeDHl/HpT4sDKoCuOe8CZG5YJvf1qUYsDs6DJ4
P+2vFXI2VCqqC+1puW8G4UuuLJvXlrKXb9lM49Xa3socccaaL8qJrx8ZzkutbTdSH9PqjThSh1Xn
anZiiXYXptgf3ZJShfMkLNs9ZqKAUFjIkP9H33jyzH9ULoPylikTg+8RKluMX3S4BKttmO0LP8+d
yaONHHBfv4eqx26bju0BFnDjx4pCXvsFP3qWuPDy/tmUMlBQtzbKnRthRnMtncXTbeurOv2FuDdc
+fnHaIWuRNlallkL1hizfYG0XaiyZ4s60SHFF9IryoehkxQ9bz3XrUxlF45XrBdvqkEMHHYqx8QQ
COxUp24IPvzjw9aKVTQ+Nw1BjUskQRxhqbG3OdArDU96UN9SGZXaJCHYGqRhSwY6quKsUzC0nqzU
myYYawyfjhptr+DoZKt7PG8Mzoc5VPXBjljUNhmrN+D+I41E6KksBdA5mm+pAXehIl6KoWF4zQgE
DU9HnHfKKpnOqrZayyiUEXiufUfaGvCjiK/w/KtWZJEtZjrjvWKZqiSa8F/mYfz+AZvy60Oj35g/
fZqf6bq34rcNItORn4kx0NycNuGoFtH8ZaShWcy3XiGxxQhKeFQCjlRLjH4f1XdUxY+DMPOI8VTS
fXM5hzRZphaKrndyHCYCq92mfYXgrXI91Jk1myCKC21lWBbGBVX1ocWXR82wrNaBEbgOTB0AzVQx
2mjtZ0fxwV6s+JQesfMpqjh9CpJMQq79bb2gabNGYqY+IQlqq167UNJSozvuNjLofnUSykb3MJkY
JnS15YVNfpwSsQBWOPxGM2suItrGWbb13Kgf94E48EUfx53JcNeyCm/MzvX3LtBacInrVl8SXYFW
mCD0Lq0H4TW+3NF9U0NXCcpioF6BVrYQd1S3QUr+yWZUik8OIXYFsJIjWLVfkuM/1jSrxYsfT/Lr
Kvp2E/xZ0iZGvpvFc5j1stbDg3bwu37Y7ghiciEh0YtyIcWOao9fB0RSFOe4SkWJH2yjJqATkggY
pXxMz6gN4hnA5TPygla8MdUpM56TpJNC3VeYV/kGbcUNjDtul0QzVVp0hKsscxjBPSfvavJ/umkp
ImI5Mq/H3x32WDoKsRs9QOk1F/uPZ+LIaCLtb/NdKBUJsejg4kwmH0CeRyv+ny8aSGUiG7QRzUao
aFO8VahtwM95J06st2p+q1PL45vz8ZqVsuxuQ7FffuI8Ch0qOjnGQyNcMhD3jHa745wI+pttgokQ
GgklV1J/UDy+GouUdQD6OXSSOnS+Mdw0ez1OBCRh81HZploqIwieQg2uQhaaVCTsBcm20NgyxDhR
sp72xLE/yN3IInfvVoNDwT/I2hQ/vRWKRcAuHcwyICDKJxifA61jDO00Vq6qx6BrRbn/GYW9WHi9
Vy0trzaph31c2Sb3766SlOExzFxraBL9XTE8esboVB0vH+EwYeaYD4KGXVdHgCXSZvugor4smh1g
LWiaIYTntwQogjUrZZ9AuvejNkqH0N+IaZpnasx4+awGkuiXmzB9w8SR9AE1iqCzPcxiVMuisQdr
InV/lb3ZTdOgO8JXzk4MasOVpRfp8/gqrxl2GDst0EwTKzFmCE5NDA2ef4/yBoZjRE7ulPFyH15w
pC4vYqP8fu6bD/fs8RgblvdXuo/JImgfLqqlnai6hllMJZ19G5jRUfSq5FS9CFve+zU6Zqp+t8SC
hvi1n5wIysjRHAzRBWJ0XDUIawnqsIwkWBWnTLhNRXZKnttOj3AoKZ4KyiTatNpGm7F0O4Eznw6u
pQTK03M2DSCazjj9cTHA6y3HUVPWtFpmz7jqDUU5MyJPp48zs9DfMRcJ/BDahO84JhmUc/LVuVMQ
7Cp2NRu5jSXUiC2mKYoHA2VjljNxVD+JMvyXK5DnXxPGLB20CL0raNhTkSz859zIJKvA0Toqtrpq
K64UBZpy1WowXOy8tHh23HqGUjILM9QSRgSbNFfUqD6+o6EOIgGTy0EiE0puSXi6Wy/mOH+fGirs
DUj8m01PVYs/FN15FmdbtYBW+FK9LaxOPld4nkUvQS4QPpyF57qXRbyRiPa21qoqOVmWHgKdYa/O
sAXdLFRi1x6CrwkzayVovDmHqWxGvhn5jtI1wFfhq4kbho37J5x50Dn98f4c0D+36IL90447p2bh
7ksh6bCVdZ1Tggia2i0EBzECeMJeogKPMH5vFaNTsv0agiExdm2uUIBSPlGbN5YmXJyysZicDDAw
tDcMzlyB0GEJ/SV43cohYBDWJk/XM2Chbql/buSn/jtDntjk0cENdVYGqXSpyG0Ge5BczNXOPWF+
cyilZaSUXDxGV3asRwG3VtY6hd/FOPQ81nGtFALPwOFYfn14TdSD/LqS6edxY2hw7hfdYDJ8Pmyw
DMwob01nUaXzuQMrwuclX3E7isJeaHApxhd0EBqgxSSqRAQvTVj8Ax8FdbcgcOfoSQmrT1fKR4+/
zbq+f4R0jPUe2w8X5ZMtii42E3SUHaEmZlSlBJUFjXzoIlhREIfeRUl87SpISZJTj3IihNHXbEg9
RQgxhzSB6dbrDurIy431en7KvqzHd7P69HI2KRq1vQtU6Hh+togCBQmVYB583bwMHDwIpj9/37Im
60ZVdceN2iwuG51/X7E44YOjehWbAOHa4Akz6kNt8gNwjoU9f/Cw6IgWeyfJ2efS4pb2AqqrvUt4
qF/smBqAPBuUFUu4EDmuxBEpQFXUD8BnH7iXP24yILfSYbSY1KznX5AobgWbZlU7g1UrxTopgXhv
q4nrttK7GjqTf3ru8M4kVrsyV0Apx+NQ9pBgT8JGEOwibBpvFGW21rXIac6PGlLUVs7Zk4uwZ9GO
k3q9hcUeiDzcR8SrZcMr6vGNqFRQOYLRzSItZf7pj2wJZBZrHyYqy0UiHPP/t1jk7Bqqti1XM1BA
PG2pFG6NOOgD6ShLTaw4L8bas0KloRc2/HQolFOhvKHpsLpW6l8561qVMFUU0OZsGQvUSGFqOIkH
TQeZj1HhEFEF8zEbDDWLdKXji2dOX1Ok8qlrWYEUwc6NmzNfs/b08YnXXf9G44+azRD9lx8R+Ky8
qHktQAxp5RZdMg45xNKZT/SaJApFhTM0yzhv0ILeGrrp0Vhw6iQgOBjhUENusiM5tcJ30ggdBQHu
ziWJ5wuqK3mMXvWd+VZAXfbY3cekIOqjrZnrpQnAtIi8EUMVt0Uq52u2cG/uGLJcEQq1z09Q8FbJ
iap8xUnRFVizA2Ajf2vOL/S9XPYlB1L6UdbW+R3Sg8melbEGzm5P5nSbhMpHeJs6SVcQSmW/ydG1
TEZjPPgKFCfkcOcskOV/J/+MV5OZvWmr+RoJRapfgT0hTxYWOa+sdc3SGBmm8uurjtf6RY12vmca
I4x5BtPWxasWULmcWTNJtvnCGnf4Fa8wFb1iNp1mvU0g60ypoiwv7WKlhmeJ2l63MqLczFO45WgR
MCNqfwX2KO2EtvSkv+sFazsGtqcYipD3+30oAB/2r2mtp5NxzSThitsiuaQM2N5J0PCvDaDtub2d
99+1bvaTrUAOKvIxkXOEt/23gPCTojbiE5JWUq0pbKvVA5AuuMvF4z2PmUewV4lRYVcwcJsycSEG
AdXLGtWNRr3118YXnk8gFlo97bqRp1CYa0x0VZkMjdDqukgxPnt0ciHlEarqd+7qZkybG/qLvLKS
O/2nRLF+LcbCpSiy709pnOTjWIwBTXnwyAvyljWRAsOF9J7mT9TSGwTz7BEcoQVUx+yiOjyJ2ayD
f7UavdYmAsyIp4TB1DIa0OSl9geQDc5uycJQsVXOpcKdnaiW6WHJs34YsnClU5b6MQ4Wc8zkMYcu
NzNd4/BMr/6qwrFRNqNqR5gYMr11JG0RZstzuNvwqqOOkaZfoDz+VbB+ONiOtlPbqxKf6y5Za88D
zS/etxF8/pAibVetYAjuDwSRQG4+u0GhwsafvU228vespJ6juAhJMoSIG+glir1Ru/vhkJYQQfbH
aP6MsAS5LVE92ArZ1wrCW5tiWjMqn77cmoNsyb6hF7w60AXdyn6m5y+reQN/VZsZjbQ4GO4r/AOp
gAFIImPPS90sdOv0BWjBz4bSX5TqvY4XB0MCTmOVh/YkXYI16eoJx+9d6DF7NkPg+BvxMTnEBAgP
8IaYML3hjM4p52/rSo9Iqa986PbPpolTRvv6svwVAseuCHjPtsiRQzsLX3D0s638R70ESLC2Vj+H
GlhOQXoc4AGCsBdQLGrEmFZ1ak2hfalXeXaBeRDqGf7t4oFphG7ZhXnKcE+jYZVFd6RIS4js1nBj
yAucf8PxVwbOVWkuoj8QkU/OcK/8NgaIIzTv69JaqzsH6GnwfRHcKFY0705Sh6r/SgBs8+WlUUmL
y3dOakLAOfCtUPCu9T/0kfShtKBZ3XOjGLCTFQdYgI24hjJ/3zltcUMgzGVvgv6uU65iAijwvYXE
2qfHBddc9Bt6wZN7ZZzAfhLub5MAH6gmT43B1v/+ZLJlPM6zDAPTNUWtw1H/+Zh0LWTL7vLNssUq
oarSzF5Bf+TEmXDwbOOI43uKXM0tuo4D2OPJ146Qoh/HJmX45VEij826+r+lQfZ8Pl8dA38vhelt
sUrD0RKJYIzKECOQXsXrpfksKgF3Osb+befoOPwHnu5zWvFKaiCs+PmiaJtYtRrBzeUb804RWxcK
eh6pYHbpAEpiozqIZnI2r7cDy+N+5kuRPhVCYD08RK/6y98kGXr5kGb9HQsD5nEdSsWzYYDjX2Ba
jEYdCj3rqFiMoD0e9rMQsg8hokngM/HVt2qm9Ln2eRJvq4S0/AXqWb+JO0ODXCetWgiHLA3hj/QM
XinwbO+cSr+9TuTPtNx/UiCYVK46lvf7biJ0/V5j6QC6w7wEgkb0J5QXfFmAfl023T4FfqViiOTN
Zo3ZgoVAJ1AhjRrwhcflG+28auGv5SaewK0M9GNwiFsMkfbzrS1F1NaarrnqooA/L2zflrPN6b0O
o2JMiVY0RTSkONUj9rhxdcuMH9eUoEa+DBUoWAT3eOrPku5KEsoZTrBmROmxfLaw+AcflcVi+Aj9
wfFsXBRw/kKnMj8agqZ4a9bRh1sIigD16aaXxI6h6Gjx3XWGMWHSkxrE5Xuiba9+AJCk/1+cHVTP
HdViDqlolvLiXX3RUKR7ZMAfVCSRWaXaiSK3IfxgWxF4zlyHLBcEcnJNPCjMlTp9f/lemdTL5Tt9
SBCe0y8Vvtj75yhn6jKcacnhKOLInkH3wRyxZy887/iUZVX/jXMoR66L/ivL/7I4YF4uoQ6Wti21
j1y4y2LldNwRzH/rLb0HJwuh2Y3rmyYMxKxTxb3bfuS2S1d8JcFYDhkLSkLBgSt2LRWmOcL5y4nG
J7D8oJ6zxmbzc7iV6QWd28Fdmaut/FaNexLEcsKHlHYlgW2eu9oEHS60kvO3M564w/nfV8AQBYD2
Bjqjjcm+Z2OU2z2k3Li8jp2tYvlJxFjDcro2kMGUMaPTIZD2s2+KzYUpgF2+QBgiJ9xhP1bq3Znr
AczpejP5iNlpzE6Rg2XLAoBiN42TauD8zTIM0M3Wa5BqSn7eQstOGEKFMdeH6/Dq8dm8klHW0Aeg
Ve2/wypkai+kej5Mo/b00CaRxLcwOgJoAmZr6R1Z8ES4IsAAcLcqWUDywaXWzDThdLvPMw0C3Sk1
XncrGBdTRDJ6SUPrvvNV6VQFWALdS/HQQQmUlKyp2SXSpqwsiI/acwTL35CkHKHKKmfvZ+BNq/0o
a7EAzaOkKfomviLnTmIj2i+tng96t16G7uf/lPLZK0i4hxWBVGgc4mGf7DiHfeEgSCnQtLNqxAQw
dZ3jrFkm7FM7sGqC1JJZEd80ScH71Tv/fQYWRRjEqkQqmNfQavGiJXAYuG8YrOsrTDzXZRY/KHvj
x5ey3Z9WQeP1WiOI9P3LHmVufBg/+fbxMJMagYEuyTsMkmAAoN8FCYn/1IeQr3Kkr8xFHKvUhfmP
Ehptrfp2FqRf84LUe25UvuJloyzYwiFNJ5TVK1Ps15bWTTnU23EZ111Rnzmk0rKHd5Il/TgfWz/y
1ORByjagvkUVpzPWMCY93ywnkv69Dt4LPtmaKbdnH1BkSU+pOLCosyQbTH/SpKNJoYABltCNzGRG
YoSDDpm9HW7yvre9Zvh13LJeSHO6Vfh48Zqe3oKU68ZFtNalU6+hpgd2x8O4APGdBbw9kiQfzlRT
Zx+oAkhXP3GfbSEEYtB9PqJFVtQr1Bpnik9x4AEAWVbR+WNbry7b5+TQ6OQpMG2gzg4whFDDm6Kd
ZngVVRxecJKuc0voCc6ztdTFAY/obiSbbUwuguC72irTifvrnj+lDPWMgqStWVi36fX+S2nI3IRp
//WI7LPO82eMuY62BIPebimD+64033+tqLQz8/mDka72Z/iv3uaXS2SJ7qYyEUoT4gWpWaapn/x+
CpeLd398En0Rdt2qXzuECTWVa3LRNCLGNYn37mGUTX8t94v5LA2jszz8WilRXVMJrxl7cI5HXT0f
sf/VSmGQza7OzhSSu3FasHc+BMnMxmlcmipt2azeBEjOfjhkxpt9ojtsOOevx0jJrN9RHfcMchxn
aipeigpBnccpNip9CwCyqc/kc0U1Xk225SD9fGtCD+1woqpfy6s+Hwt3znNVAAayA2puD7CRvVan
iUneNGXMdpaTj7xNEXD9nIRPa+cBnqofDvx+/6Hj2ZtNoX6zl0BGZom6giq/7B4sp/JAcBvmtswB
ohNdpkCsB9xUjT9lY0uaZSXajsENu8iZqX+us+Jkn2KgoB5quFhpCfCS9r2oct1gXRwSk3LDzkMZ
fQWVt3dLY+sgIQ1HYx53XVtO5PPVf7l2iDdF59+8iaWlz5k6BusHo9Kg9BITFFmHKaDgsXwS5FAd
LebG1+UCL1adYenPOXozSIVpDGdgF7kVUUeS8QSfl1esG+1WAjU6GCmazV8cM8DwNKxaMga6G01Y
ImO0Qr8TDsMzFlW/rUZRLxciGk5R9NXJrdjsjeFrZNoEBAx0ZD+YdvoJExeyPdpQkxZyq7YZpyLv
6flc/fp6Et/V1DQDKwTyLeKDOdJCJcLbK4ZS07Hb8Gv+LrPNlR5umxwpAB2UkBjeKCaiQLnw4iUT
YDGpBxd/hM/Xvm62KakesPPaUXWwt5uyJIluPbk0t/Rl4ojeI7Vg18cTHINC5+kQAruP9Ng1VgEe
JXgdkyDlAPJYDiLiJkgHOyqMwKIQ6XWBW15Do93OS/Os1FjRhELuSLDwY9D1q9tdBxFy2c9+7feL
2qG5ZNom0DWJ5cOUM8dh/28mnYpZjPEN1PWX8bMQuMqDA8nJlZufr/WzbGDWrXbC6Dtc6YS3AQIP
fBIfJArpuMpk+ItbmlIoo+xvBhga0plR9fbVVc04O2wxm94U0N/M2t1Nhm+fgdTEwocM6dE2GFFm
aKlJurSkJ8BP8Co+Hog+wM5US9ufU0eBNWOMRNPNUNo22zDn+LOa3Wj8PaIwPeglnJXaVfEzR+mh
yROQ8+NhWsCzGbtF0ZstPzuEfSFYKQUebIKUdbYmOnmqfU2T/Ir42ZVe+knS1hrhemlXw5FKMF2G
KGBao6bwkjIfT8RK9UjRi386X+0QszLpflfQ6cvvB7ZgLJTenDg6IpqtD8Wki0K5jur/hWU2Itzz
78ZY5Unw6OdqK7HixOHgCkZc7CyWJgNQYKlqSB/zKVHLEjbzcGZGsh6+fPdD8PX9cZAXgrNNVckQ
99EurC5RQLIOCrAs4sVe314hHllPMcfpWkdhrZ8SB9E4+BegYHCwN/JvbaQA2Y/7zLwaF/f76FbP
sfyOhuMWcCHj71iENYG/kHOnMgjwvVDnaTcZZmcyvsZaR3rv0WHNG3608ze1R3NLicxKZy5DP17k
6QSUoFj5Lyq951Vy5DbQxVuy7EmY4zDxe/BH3LJQ6eHeqewb/mUYTRjhmC3WN6zq0hVMzJE6cvHP
56zIQeWF5JvSfVSD1wzhEizPjnaT6UcUlJkzmS2uTebvBW/VII0UbVhBuK+J+jSFyY+NriELYova
kRJWVRCGKtMynHlaugTu2YGtjLQ+7JawWiGDn+5SOYipP4IhpHgx1MsefjDLw4EansBRsuq1W1zK
fahsZ5jztEtVtvpE/56EX+DDGapfv7SxgpQODggcWEJvqUm6bVcRk/ZbrFbfN/3dMChA1B+HtK6W
s/5gsLvSsdF5Qd2HmM67b0uHfHCNkUhqzY6JnpImxZbDkNBVsT+QcbeFFQ1mraueQjoApb3I5tax
SuuBImBmuOa+ogsCSEtN/tTiPx2Wn5wEsQA/VCfI6UKMcsqnOOAxN0xYT3TTeU5i1dVfTBIrYlxy
pN0V9nLD2yVvXkpSvY6ID9cLxZNsj5DSEsjQRoAYfWp1xPmgp9tTk3ekaxwlb6pkykK9eMiii/p6
vb2Z41RGgnQju+Q6odvdHZ+Nq3O0E23uNDOdXMu59/5mSbQPcewUSglAZVejbXL2S7bTNwN83OQD
cxMES4flXSvgAMgoPSZXqhIAWH6FuLYneDadbt7a4HVDotR8e3vbSc9CJdbVkdq0dUbNpxfLl8OW
pjQjSji344YMvSUs07/4Haaf4oDEnBxc6rjGU0RTWkLNXWXK6UD4LVKWjCJgEMG/Pyz2/UX2BT05
gjwKPOr3Pk5cAxZCpqXLaXVyP6tN1/5+4ghQ8ieIxRXjrfz2QOrWqxPwXgmQkJAfIih+HzFVScPh
ysct4S8xSgmF/ZAicQM+e5av0Nhd2vrJPioNXwOntscqx8gRlpyE7XWpyC3sq2kcLMkETw1MtyqD
G/MfyiNSCk2h2rOawlNkwSM/D7ERw6bIdSCyYcUB9OUBTZJjwEZOF9szkaLGqHbuSSxVrZt1IML1
jS/L1dgFIFpAw+Pz/9qfsYrPS/0gHD95QUzAQ51bpNVmGJHw52Lot42PKFiD4b46Kz/pbrqg85Qb
ql8xR2px7MQ2fhMCxtMa7fZs5+0rip0bTtNEtdpH4+qoJZngxIoC78HSACLgTDPxjUr2mAcTgBmf
eynfe8a8h3zJj9KkvDPc9wtMXb4n3imhXe9c1WI8hrKoDoBzlK+orgExvTMEMSGVDk+ECfvUTEeA
svQCh3sPReUrvYO67mu3siCMo4FUUy+Y3skW4EOGuH753sNlPLvGNWZsIDEx35Y0lhgyQYD+8OVC
YceJqkuWdqJ/g+FeiFqQhsT926sx9d+DFxzJ5Bb4rqqOcvPv2Z59j176jabWGHdWYIpitRfWtazD
RVT+Uci9ZbQ08iA1EgZvj9DMMx7XksZyOYGmBjwzbgf7YUSFBsVy/Z9NyIFCrYd0WQgABd7FS8cE
eKMQCniith+p6pVqv40tQ4fv2WfQSaMI+Zw2oWL8aAluJ5d8eWv9KTRHVRwxC3l3g8cNnhWLKGwN
AvYkFpSXS2UyRibrI0cprOtl8IqGSU8oeRbOJppQMjTnfO6p/r0WqG2CQAfW072vp65wGyt4tDGo
4z4scsxdIzv9BtpolkTk4vRJmcij6DCXZ4vJvQ+4oBrC3nsFnIg9PIJogjAJ6fXhERqV/983f7ln
wbzbPzDAoXOZxgsx3zFww/AG94f6Czb3svTBjoy2znPPwO5DqZehb1U0M44k1Pwx73yvGBjtD7Cq
IG6sBPsB/wrGsnJ4DV8mAyPH6yO7xVeO5HEDVuP+VoF5tjX88KR/OsaYn9xDYDcw+UelrNjQXZzI
TY9MfQTjVx7Wai+ZJoi1UjI4frx4D2g/LFHyTUrkqcw2mp4LMIodzCtmHfE3uvjhu1pYf01VZu4b
o2gBmlVaYbyEchvXTCp5je3zZhweETGmXH8aEQnZYqL1WRxwiNergT8kwYVXz/PIiDHajj1Kn9Mc
KhnteAu541DAuGnpIYKX1RZCFZD3VQdLtGy5EZ7m73Xz2cMIW6lJTqlsqFgVETTK44W4wkyU+UFF
DqVPuNAcvK+BOuxsZCbsX+Bc63q2UdrqUlCycXWhSl2HlfPhIe1TwMI7bCuhF/+Brqx9Kly/6y9N
/dc+UtUzwwRoZu0CYloyXujP2P4B65xELdTEQz+cWSVwpAJEobxpsW62FkzOLm3Gus/f5SCGOovF
2cKT7m3OcVqvHvWItYrDaC8R5ZxScsmSxWVfg9pRCB5DquqXaMfKSQpQ3Ou3p4gexV7O0pbxq4E+
FO22Jxl6dklo9K4kbq611NQc60bg6+fLA1sWpi3uscoweJIiS72U6w5dzAvUa4yhzqIXRnPHyJov
bhSWMPAJwhIDaJDrZZmkiaArz65zYcbPSGSLV5nLwBbsYggYzefwE/ogxoXWla+/RuwtCyNl02CS
oYwFDKUXEajjhtvcuAfyNX0Zp5vyPSrqCPiq7KI+1JeEBaATzsgGF1Wo4N2q57v3O1KwLVHVEkBz
MAl1tlRe7AL5tqBfdgxHjaM62Iree2XTEMB7pCIiGOtiwxF2yjyskOIRxj5ELljVwpnHDYO9C5i6
yxK+rGFunOhZ5ud/k59tr09Vjnn1Gco7GTyeK75guJQKvecHr5Hcrd+wFeI4hQCMTeDXoPwid3x/
eZLJcfAmrkxQ9ThaMc7xcHJ1gQYybW+/Ei1tGLo2aj00aiobtTgPVBKNYtOO6XA+LMHE+Hozx6/F
MZ3DcMIizm7ASBc2qzGqILHZSavZCMSQXdZJ4MWl1HNZse2zeklVMqRIkJvxYdufT0Wi80+T89eK
aMKKbkf/o8ggGlan4AOq846EjlA8eX+dMzkT76CNmWeminHW3JosEPjgASvgGkFCHOIqFu4volzT
IyMTl8W9VFIOaKww9RzG7F9THXIUeKznwe81bXD/c/fFPClJ5bFeXCdr69dNJGQkm18SPnHUBJN4
r5kFc1xb5ooCFmt2yrCHF2PZOV6eUanm7VyEfL+fdJXEzOmY0bjgsRhrTCPwVYjQP40sYSscnltm
ZZgKOf7l5tWss3TdJ2jSMsYHGaoHoT2EQS0QAiGs99KVy2iFS/Wwts7byG4hizQVzfHNynxeHcFH
9zPcBWEyDRjn0UYH37v5MUEQBQ5I75z8iLBTPRkOppcPOOosSQxLR1QNheY/VrzJW/NWk3B8MS5N
uIw1LXouBmmNoeb9M4d52w49QK5ziqihNh3WeQ5iiCikhE37VUSWtLwaQhsPAruZ91zx62mn3LfL
P8HDNyNxNjGtohd6BKVA6W+BcM9jnUO+FwtjhU5gr4+n2HCXzqaKtA+DwhuolqskUCD8ExCeNqhA
iloHJKJW6Zluj9MJ72jGYT7L/GSq2B9Bgd2nTminZK5N7ahIQvuX2mI3fP30BkTHViHDq6sLWyfw
0HTobYMCeuy1DIu/OCPDfRLdHk4FZp+DL3VoodKNqUrM75m20M48/k1EgSocCUtZIcTkIcm6OlAk
+6w1gYiR2I0ljYLOGp/vB+rlIZM+cd3qOoTTMyfLrYvsKQHD4ILzjnS0APD9PtUp7r1ZbKp6QfdV
Al7AU3P6wkWF2BH9Sipflzo4jDzQoqah45Gb0Jl7VbVeQiMC2cL5i62YoAFwNDhT2+cHJlLYuKQZ
P2UA8NImiZHJ36ZQ/y/LhpWvSgQP3NKGqPp2OkH6mLNPmVTxJAH6ETJC4ouo+G+qZYkKxNFMIYFQ
0MVy2J+vFvdSxT6rKtS18ltujBSd1JKBDjH9uwtWpQqHQcqE8iVqhutvIqDd2WjIkOVXseIOSsZG
Y3m2MmDerCQL2RqWEwBaytjUmUV77KBTCS3JJSwseFSW40PjjcyrHOCIXSLfOKn2XvtH1KB/NBcM
IkvbsVpVu3TjHdybVEvvnqub0fMTSTdw6+9G0xxy2S4qdhAQH+4khALEUYlKPEboRIkpQpFpHhra
a+qTQeiYTt/0/YYkC4p34LbgCBi7ikIXfBlUNFR7H2XtZjGtTZRrHOlsEAezGjkyNwOo51R8hGRu
8q4vJoQ7PtJX+/99Oc0GcExD3Hl0knLDYI8QUlXwifrwcgZpV1lkESPSVT8muDv1oLx8hbGc/+J2
gFYNPoJ+l7rLgn6wsUinD2spCj4Rad6XHciy+YCFDmqgrwtQK9WzllAK/dQWr5AqOeGaayfnMYsY
D7F7oS54vg/tlJ0lgWqtctKVptNGjc9BHnKDJMZapJUmFsdveXOuPGoksh+LWde2dGHzhZX9IOIS
mM+2V6gpUuY7pXiSDeF/UfMfMZzeZ/pubLBu8E26iN7d1KpwGE+kg+lRju84FIWRxMX0jGlQerz2
sa307AqWZ3XpGTamu1dY4qSiAd5b1U2UZ+VxB75+2edawRIwNo84Z5OxRWO/GMjUaUNkQsPmaDJ6
O7ZQW+2qiV424Obyn+OEz+kfiVx6V873FAi2JmhBxZk61CvtIZrly4DC8NCqhCyS+va1+XwpO/Iw
+cF3iBPesroCvXEtobTOooS4pj23rDtbCHsK+6sWk4ADWr6IMIq7sxYVQub+DmNC5g+vZ3ZgWysO
+28iRjxgobylnTMWiwbE4X+wPQ/3lALjO3Wx9GxCGVOqRz9vgEQW6vLmDT3dSk4YHux2hjkL0UGe
zGu3bvV0XUFQveCg4SulUeLfpoAraGaA61xkjHBm1XKLfPk+p96cJDlADuAYQPDcQyNikFGSSHxt
UeGDAEfxhBWxXnnJySmUIqFqq7GIlkdlsQda4sx8bIMkRK6TiEAzhm/neecsl1F/6c9JnNjRW/EU
k5piGX4lzNyWVrVp99SPyse/hXO4CNrvgp+hioOsl1s7NAsGsXWdqdP+gJuvIxnvQ5p+BHqsIpWJ
91qyXf2acPXUkGkxrKvLvZrYaEMKcgM7qZGPITz8pxzU1LqQAM/0Ko4ZNAFsGvjXrp1OdQYmMTEc
6Q7+7OC3TwmchPCNMJG7zhQj6pBaV3WK3WrpDL208H8MifcYwjVu4PqI0i5j7TgUCJw24RgrbjTk
AWOMtxxQO0iOUJmsNY8BG4ONOAoSe9vjFC1DtDlkPHXpGaeHb6V1VLQZVXA63nPnE+e9r/9XQQFb
6H/lpnS8F8t349NGO7JbkF7RmiFoZ4x/KmvRQ8d9n/Wm2DJEZJ8Ilo8AcRmwQTHjByPBhtq9PGkt
zcspsOcPjz64DqQRTMk4wx8LhQ5M+MgKZCVpDzHPgXqOjkF+k1FIxKxg9IONGxFp+lPTYxU1Dwks
3k6QaXHLdlTUxhkGfVpY06QhFl+B7WuokW1Se6lVObKIFv5oD2v0HCbe/9d0wGs6gtPr5EZxCR++
xDPJiAtClrP7rkjeHPu1FCq5gkD3jSJlUxJg5HYR2viv72RbKbAgs+fjs8ntp3KGCF+KSbkA1EJT
rakQEWoR4pPWZvXniXtk3ZDBHle4/OJCA+ZqIrGYJOo5sg88ijBRGUotDfrlHj6IF+DQANrQl4Ky
O3EYWFeY0k1aJdNeKlCjy/EAvuvB0Prl+GbK90XNXZi0GcBuxXX77qHfOmQZ5vCX3J8AXSNVym9o
k32vHUjKs7IJZInZBPjUC8oM8uTaK1vK6JJCjUKKnpHGFlKZrUnGCfQSWIM5q/HW963+fi4fsLxN
DBl58A1yuoBQFsAnxl8GGzZdkpOVF+1slTjYtvYunsivM0F3Et1MXyPwkhfC+qUwi+GBP2fyhZQU
LkH4nIPbpOa57Zko00S3t1CnQvywGzbD35nd03NTPsNdDatxoNgFP0TuO3oJBaL3LefaF2cME82D
rdQgZ6jzE7OFtJtCALvt3CPBNAk6yDPQy71hUitK4aPav3fMbAC5eh/iII/qwrSpYk6LdlTBwfgJ
tQWpEaDdrLEQlDKMQVK85Hd5ttsY7Cx/AQDzq7cp/71mVukmTQhDq/g386Wq9dFcEjkusUsgaNF8
LCsi+5MOu1E/fjA62fUSXRc98uhrnf5dHeuUnzBf11/LW0dF5iUr4fju+2vCyaUvM0LfBvVC/pbY
GjAXXZKm0nq9O1mHiXqRKVZahud9qxqEj8Z1l6jG8G21hMVxWSeM9myITo9AMxraYEv0i3sxZdhw
9Hvf1+xifMxvVdoiAXmPtc7QgOgFXxF9DwlrPMCwDGQlhspyV9sCj3G+laNATXtoW80l/8lrx62I
wamwgQhU+ArpIupdteZK8AbVN8kRnCsCsv5laV2QjQvsstPi9PZ6yffWSCQfp3aJRwEqXUi+6Hu3
ts2agTYAzkIoV4Gi0yBDQWmOtMwhnbHTvYhcrjr2yfjN1TLQm9yJRaP2nrdMXVEsV46mMBbtcmtg
1V9Dw2xrE3PnUbyHBbKFc8jh2PjMi8uLjiALBf6zGophW+rmYwia2XoYOL+JNZIUv9IKenvVerG0
YwTlLMa1mNcgYs6eKuq88xunVDlvtNTC7k8+gGtjvvOBA9LrK/zxcHfYb7FReDvTV4mm0LS/lskY
V2eN19ORiKG+mRojTfhx7FssIX9RQXlgJiFPJA8C1giLvtOCKE8bcUx9t4/Jsuk/8av0KnhJfm0L
wtg3JzAphHt8iyG1RcvGm3sVh91JYrkw4jBRkFHU1Th2OQ2+Up9NCXOMJHX9erQFnmGsTt6/0k/N
zt2U0QYRo5gMJAcBZWrcaYv1v63b/LDep6PkcjAJH/tnLocwVsVX2XXh5x742/I15F+IFHyua6Vg
BQwoWGofhbQt6S7wO9QG2XRydzEPjtZUmh8I4bi9OQMNeF9YG3FQimW3O1aQpcLD4LDYcLQvhp4h
XBkDSsA4YH/gMfJcTOFgM3lSRDHNKC5iDFKm8xfo2M7DsRsrjjkcQ3qX58PCk+I+IGUYwxmYKK6y
PF6nNZGQxmIYyx+Fvy3REh6InkuS8371VKU5+4BMxnhLnQHAsq/hfcrDGYLOPfH47kPfQhw4Nf1m
N3Z7dGSF0b51udFv5pM3zyTpc61KU6/VFJOWzmKcKPXV7M9YORfqIX6tOT0v3DIuQa6Q4QgpL4Oi
rB7D1ODH7COAmZmO9fMHSGxTPApqIwSWLIpRF80tmtSC/rKmqK2DibGbl2S/adzjhvh3arQYxe/1
T1hq0h4tdsoZpOKJ6uamfKbOQzg8ttKZgulsUqEjPtnqixDa3KfwYk6/wDWdO0qJ0lC4jQxyMCaL
DRqyqlPHa3be9jgU7ibn9aBCuvi3RCRNNuF40YKaBgEHyA03vUj87sIsvf+qn9XZrDefy3o/i48N
CXfnfv0zuzf4wz2cLccApZhDQMDIaKejnKPAOo+qcQU1LrDykM78zfMnfLsaoFUi756ASQAiUXYM
PzTyoDnfKxM7yxVtqu4DY0vi+57eZlriKm0eEH+lcHA7X5YInb+HTUnAYf7/FBZImVvgndfHNwGG
BAfMcWb3onyoyCRO4BMJ15k3B6neLNXEfHOvYbxROGOw09YhQd7ghnpyC4+pMggIKQVKNX4hsQ03
QwqPPJftLISbqNsXIjxjQEDUDzUkc1Q5zEVttEgwbHrQ+qRxGqH7oIDea9gviOM5wWj4xse2SAA2
7ctNgHXhfwnXzkelvf9HotTOu1Puy5Gl4GMeJr+maGhn4IHy3R+E2uu3U1CFoAKT/h2u/eU6C9bI
tulzk9UpCEHzUNpuDrlxZEZF9X6DPwgKbxIN+gjQQNdHr6vM5HQhCF3pedbSL8WywkatpoR/OlX6
ajH41ISd1WQGH99cSycGwk+UoAOnfRJkzaVt2aulv0vp6t0pdnEyu18FNKBaYWsL4wXyAFXZplHD
gDM5LTTGIJFyfmKD60bfxE1bbZdDUi8NA6R9rmrZ++RqFCKxeWRyLDoyGIzjaB84mG5tFNeFNfw4
afZKHSFAgeQoE+hRFfkuyAj+oriwELe+NOocDNEoBOT8oTkDZ4dkI7qQ5l4wbmJ7ko4ziwU08KKU
w0szgUfl2y/CtSFdC/Ae78OIDWeUid3wx86sUJgd933wtU3dSZnmopstOzYnxhsFacGuwFHv+DIS
uxTyEDoYuvRuw+/YV1VZ/BvAV747VkcBaJiUjuY4i+mLja8ecxl+HfqeaOtYPHhvL18BkfYIfhdH
A5be9s/5VXSl1V+IrJHMj7UOsdL4v9kMKnND6sdhiNuK4j1pd2DwWCpsGvupBBt8yf8f41mkYmf6
7V589o4UzUEB5YHQ+WIChKQvZl479KSpGqJbKF8Hj1AjlxHcj3NYuD+6ulUGyqHxg9RnoSOC4RRx
lBstVQmBteXzo0y8XQQglbf2KSH0wqOxHYL2zZL5EIcWRcpuLLfnrBFPsW7nZ3/G1jAKBNlX82/8
GL5ZJldTkLBZUCPGa0lrqMytbXaavqwDpwY9acN4SlWC4u1UYS3RjdfWZ0ozZUdwq4rk/8+sO+gX
cENCav6TB4Jtyo/2I97z8jvxboQbLx5RJ38aX5HkwKe45MrXfIsMswnmjKl2Q88GndKu0QbDJGhD
Xren9xZeDEYQP0jBsrR2uxGmg+cmv/qWkFgSX2Wef5IxP87WfS2ZX2SCeKHriztOcHS+DCtUxs3e
6QnvFkAnvlbxCmgVhuOZd0FEKxctZ6YZ/HzxvEEPBBuuWWxCh9CjLEeM4eV4w+7Qq0FxTLQAZu20
sU0Ca1r4s1bWahcOqqkma6Ma2x6qPZpAJuSNNIzuZndO7FrYbl9OCfI+NnF1D23eb3Tl6PygesyR
U32TxPM6vQqwBEuDyXMTX+SdHUl14q5r7bthB8bGMee6Tyn3AH2Ht2YrH7bJmGI3cjeUEt1uFfT8
6ZwpzvOHmXwwP1aNqGkQYzxcbag2x7XiBSO8YBiUmqbpY3VBLHb/FKgJGBpbKTFdxZAPPoDwPOP1
Q9FlWYmLM9JDXhHbXtt82hwz0aNsTBJCQVJQrh9+cc+CNV19yE9s6k3Dp6QTQfT08g3V+KA9J77D
0/hoBnLxTosO/iXphPfK/3x4XTeAM07O2Uu8Q5OCjFu6DEFObbI7ovEAv1l+PyXZ17ARQPqUrZZf
kmuKvHatHumgAQ5PSzs7MFoJjY+6w6UOHGqY4MI9GMvYuse+AGipDWEW1C5STsitxXEi1vmNQhKj
eRihYhkT81PH7X3jC/4FiBjtyz47of/MYJfI8ppjMnAJ+f7tAwagweGb5dllNFk6oAFm8XKwmS15
5KNdN3XIJAPP27dAQ8+f9YMUj7cgaAq9ipanordM9isjZdVwAbCHN7HcXgzQtlzzqQa1GV8w5mVz
nc+bdHb+WsWtrn/y0maMkvblpiPlMfMPuUX8JSaeyYuVtUldgKWiGas//Os8wY1Y6QGCV0Bw1jXS
oY7uCDYCXU2G+pFZTcy2n0t/SpaBU9yKuHEx3vMXbiomA0oUQ5Plud+4aZLPY2dWTGVKOQzmj2nE
+D66NSz0+e1CT5oHKCgbPvlggeFQ/j2swnvkJyO/4MMN3MmNJ3rBx6FfR4GJcqoIca0eXNXRRsHK
Sw+nUPyFCmu+3l6Wor6Ndc4+jk/dO6jzzi9PsT2UdFqjO0bSTyTFNaFU08t7zuu1yyNFrz4t/Xpc
0JnqbNTv1qFR+RDWhPAWmfpbfCqm/hVdi2oVnTxa/DNju248ZsJEXNmpeIsn7hUylzm0zPJvH05f
Vi1Dr0LtIUM+uHDZkh76dnDkcdlVOUgH98GCcd4kgTLKRO+dq8BlEwwg9d2nkNQsrf1vq6fB3/WD
vWRJ6R7sZa6x8ISTay6feD8FvcKPlwYyuGetwqYVTJTGZi3ccnctcc744UPiqU0/e4JPAbSvbjOd
YL0q7xt2pkWTNqQPOUXlGdFa1b+6P9cO2zNVYMY3DLm1rXp57fv4j1oE8O3x63NsEItxSXTtlieb
7bYlX8kFf3+H+srrBfXn4RULQ4lbpHLNPZdKvl0wOLeKYTn21wvYbj/3kXytxsxQYV/jxHIoX4Zk
ozBwMJkN5ofMHuWZJKn3rWir00wGmHY45RBexfmhkW4u6p6DbD/MEz0+zAwQQyCFR5x0v0XoxTTK
MED8xDgeTBGXkPMf5gxBRKs8BTSXq6bhewaY0l9I+kxRUGj8a2gbY4Aby4PE0WAHh7+6RQqlz7HE
Xkg7qMYcacFLLcJndFv3hyajJnypbTzj1311/EFGEMGh9hmCgXCQY5ORi2v/WTzXCz17cCoalYAE
yTHtsVBGPc53JlZIkIPPbjlIcWWJrRhVpWNXpLGaKzLD11Z3PRkGhouGM3QrDi6HRccrRC3o1dWV
oKDAcu338bU+/aYovLXdIVagpGwn5bNSaj8JeSarOtjjJq9QHiycbUZLWeR9QlDFNFKMvA+CzXl7
/1i/4+hnpwUssNIhMbbvYI0DxHQED4GuIp8FXKIE7qqBOz/fbENiiw+JJEAOsUk+znyPmhNrhMp6
M48lQk27HjY3tW5arDANB5/62J2L8wK/HsEGCm9oVoGHq9RIdRcuXMtafw6fYCi7IoiO1bddjiDY
XKHqxknsPFLjEnBKjzhTji9kbuKWDJePItzn4ohicCy5rCeclntPfOyL+tiKTsHlHmFnWJTnhtGW
PViQcoIZ4u9d3yyAAhM4VX71XfJVMj/OmL7rFBBkLllr4Am3BHTwx/VF+VBkWGLD/EwmJmlq20nY
TdRGCU/VFhQDpkMH4DUzLXJkq/v3Ih6yC6K1wA1eSAhbJe96dXo9/8t3NpQN/XOUVpgZ353GNmB/
/gwQyu2RbM8fNOaBAgsnbwzv0TEfxDyakVxpCjSU/DG4uQjfQui9QSZtpfGYsfBK+4qtP+oIbNPb
620yTIOtUleePgmb29R69Pk6WZfeTHTs76J1hFgDxbPGzM1l23iulQlCKZv9qlXypc4LRI6UzMk+
AlLwNJY+D53cjG57siVaed8q4ODD6aSbXhCBD/mbv2Q82D19LdJ54N4byg1plCt+JOui009DEGpz
NQP4+a9vdVjWFES4pA2+YMgmq+xuo2QsyRkQvhmxq15LHGoUbP0eBTxI+kd6IXUTwted/yAQtMe1
fGoAraxhR5s4OcjJuKXccDiHXOWPDgu1huTh/XXSt+DbV/Idbki2aCLRxAGH8tSP22lNmRY2+t6d
Zuy7BpcBf2P91Ok0wRr+PgCKrQ8rlDM7Zba7vuwUtzMe+59jOu75b3tPREfoSHITvokJTAoODwPe
M/9tD3mTPMQA6Tll8ju75c/I0bfK9SjmEKiUrgMvRCjJeidb9Az5L2eoE1PINKVMlxe3+E2gEolp
MIqOnhDLKShb/kRO3waXiwcD6fCyroftP5TiPesneFocJ2eFVHkJl9zN9aApuatUuiJ08+67c1Rn
u9Nwuk9LXa15TENQXWLu4IHcgcFmafm7TnUSVW6R4OuQuy/0ALTKuApJSMa0mrZx7yNAQb8y/otS
WS7HqTtvLjjQT1DT7G0FK363iCsI5lgt6yIiIjSbRpO3JGBABit4JSJfczLJh0InyQGSPquIHsfw
e7/obzV5h++gcy+5QjZ356b7TijoVHZLUBwYeDSUGAGY9NBMjTFraKIwob+sn7KgqQC9/dzD57L/
5VDRKgMSHLNDfRIXxVc5uWzNrysz4t34vFC7KYhKAlFW0RoiY6USyxJwJyA4ZDeGNrlcEzDPwtA/
9fupW3Z6fd3Z0SUeoOvWmrlc7nGFk7aQ4h0jqyJIH4tYIO0FKBA28zRyXrxnbEPyv1zH6q9GTjuH
8B1c10aeCZ1ElAZxM39n9k4Z9rATvDRT3TTUyO6RXSzZpQdF1eYP5t6WgVvVg1QRlljSbnw0nAK4
zCl87YSGajlJt/V/vqmE9rqaGVXZMVHnh1/XMqx2NPshrgahHdDBQmJaMPmX0GMu91NSokwRFFit
xXo30cF205UaV3gEmspc3XStgGdlph9HBoNCJuLebgYoJ5evJ4uT3xEE1jEHejAaL63Ye7aieQT3
1wERjhfO0sTh6W36ICrE9I0LtavwbzRk9uKkaHs/1Fgoo/Na599LRLKOIyAkW/ahe7+turEx8M0z
LBIDTyrtAFcbW58NMNbZDqfDEVvjjRuBstZxrSKCLdc3VyzYe6HQn5LI02skSzFL85cdNwuNvwVM
IEK9B0z6cAxeFHnGmFRqifrQdeMMbXvO0MXMPbdgHQ4WAFhBLdIUTr4R6HJToupFhBJAAM3qKkfj
t1lPtzfNgAf2dIEQ6hy/T4R8pdsS3kSi8jPtQFdYE8qRtiq2M2W+L6W+wRC4KVmNA1YlxueVt1LU
buOoD+rGJwtfI1t3dxOeqke8XKUqkWePOn+mjsfmo57MSyVLxh8HB/dtAJAJIqsZ3VRC34CIP88+
pDmhwFeJoNTOIw+5E4ST0U7z+eVbKKOO/lpM+CaC/DXJTFHhXLKvv3kudV7U3Ek2UjptGk0htpqF
poSTwF8RSHOyfO1anYITSkjobzRcgZPvvK5K5TsN8O6l+hsWzZM0aLsqRtLWrpcq1QfiO0im0F9P
mZP3sIqIeBrl9sEjWfR9SL9W2UhI1XLfTu46qt5qx7UziWGp9r8Pthc87XXyWql/pwuR85xHyyQY
QoSTdDBQ/xB1fQbFbsEiGxRnHO+4umReldLduJI/4loQM5gxbgXTLoS+THukmaJVCfa26/iTmAWu
/AcBWqKG6yfvXpxAtOxhXh3NgwpOb6bKHIACX/mgAFiwnCiAadmEZF8mk1CHo4SEeglbhGTRj93/
ebrZS8pb0QYEV2oGA283RDTptOmLz8RDt9YLN9B2it/uNhQtf8crgu2gSktxtAa3qGzo54kS9AEo
udB8TGMAcTeJW8VICWy/S3rspc0zg85gpUVnFqHuhWSlECif482hngxLOKVRefhbTSs7Gz6Ynx1Y
wqIONKG+C+xjMuwcuFfwLyKDdPJnYUhL+x0r7BdvmLMjAqipICERx7z4T1+4ttm9D91l8iswuVxn
IBtqmiaxQHk81j4azq5A4rotT4wP8lwsNdRXvcbm3QqM0IQhjpEOdgcZuVrY2KyX6Fd0QIk/uKm9
Ma93QmHqOycLJH6X01AV45GGy8fpuU1/MwkBMiXxtZWhQ95+dr9l3dC5k74i44ws73+7I6WIx8L1
WWWIU/EdGjPo8Jp2B7aV2yw+WnFQ/Vizka6w+wP8s8sRdYVgwY7pI60o8El8852Jyw763C29eUpX
QI5V1m8gbOU6ZGumRGD7x91gTYQV/piNur/MIM9+Gxx/NuPvGpWtQbe3LwmhOhnvOnpZmlmR/Vv5
eOMnTywCvssCswLDcHS7swjmIAW4dGOSRiBRHZTaLWNzPsct5tudZyeFSxuwDFrKTC+twbYKhI1x
/4iZBZg7f//lKTsa63UvEtA2aOj8ouFbzna5z92H/YLzVQEd6vq+6X8VyTz9HzvAkqcXb6Er4ilO
O/Qg4VnvVW5DWZJAtcX224PvsffZQQ0G4kYFSDhcylxUmWXcCiCXnD7C06yADVP9i9sIW+8LWHZa
uXT7s7yadnBsmbDc04ZF1mfdjW83eXHpJkhwE2zac0DFR9rew5sRjKru1uRM63VFEbvZ7soXrs0O
d7DSg9GVFTX6kPP5mBedzOm2DhGI3bDQUJd1wmAxZdb3daJy0RMq2yVjI1WWgU8ES3HvJvxK/ufx
OD1y+mEECR9V/fihCg6GZWwDy9/i973+vkk+ay45nu6udl/s0pb9WQMrJWBmuLBOj3G+bCURjSlp
z2I+EcRwtDZ3eq/TremskE4MafBUQl17Wy6Jg0JVHJuALH/g1rkPEgU+313xSTPGb6tonk7SFYfo
JTcH48QjE9rRGtQJlrRRAHmGBXJpndvgXvl5GrZPE+fQwaaRmjfgv8vqnZSbXi07o9MYDmOJevtS
XeMoIW+enaOSTyAqPtfqJuuNmwb8nkd3joMLH6/LXd0kjNrxUm0o+Naubue7veiCk0rn54zT4zJC
CM/BuI4nijnPOnC13i1oRI897Px32x5dDbYSZWrV3ALDxR+bpEF8M6I7mF3O8M8+5C2cKi+EOJ/I
AakuOG9TaQI2xgREdHblKUnYtaYVlrcKOX4XfdkVgPRUxahpT5GOPfsBhxJdmafpzjj7zExPskSh
tzBt6j7LfmL+MaZato7ep9KzSOlHuZ9mF4wavnq48HfO7PJR1+19MfTDOsmyHehRtlHPJpvl059M
MhnU674kwofFexZaaROu87vkzzOvfuxja7m3G8bQpLNx8gvVhzS1Ce43hxDGJoflqhUL6r6NIPiD
f+owZXAnAtCg2nDZFEIRMSkyrP7Wryx2BBKA5VY7zB20d7J3/3VQjvfdleYh1NEDhGM1FhZIlVJr
k2RZH6ECHw1/9lEExhjSPPecNIWynF9/v3ed9N/sGcthuFxyIc1TrMhvwams2N0KM6BGWjLZqAxb
Qm1MxkxCqV4k3q2jz7Rr73xkrZ4dCRfH6qDolyG46aIXqRUoABQVBfS6HL64GkJOHZRvLeRHbr/W
f6jWghWpG/HJBZsQdHVe9LfKP66mN3UtGkbcvGaGShkOD8tPKfO7jVk4xLzqWPHFtxLAPLX3OKBP
Z8FLJKYK53fj1Zmq2sw/WfqlR++U7EpHMPxHRpwVK6tDrTLGpJiooOv0xVZiKQksrw50TRxPCHze
AySL5KYYyAJ+WU1rR2Vc9zLq57rdcUSUB3wQp8EbvPQKI847Hly9Se1gSmDup0JNACoI9PCUkBrT
18Ylp+UI1vwbxCVTTVJpxiBXcUIX/fnP3Upfe7TTZl/2gEygCFAcCDxNpG/YJStjdbe63oMECUZo
hGoTl0ug4kqRHSicIQ+mFlRyg07VSRWgu/dJdDgJJfl1TUWHsdBxpO0SLcWwT1okrw9JU6Cf5kVa
IJwNLbCbv33keV8i0g9n+tlIhPysLwHYc5Gtv0gizo2qvNyoaI6xBMw3InJuLyDqnn2yBlSLwvc2
0AOJSHc4RYCvrwwmOC6eG8t1L3oyiXYjShSRMH+DE8E4986Gj8CcQvS8JV0+6wuWf1Qx8+MRQxKJ
V/8GoLad9qSyqp+GupOaQEaXIwzjb1oDRS/CXZ8v5UNO6Tst2YCfITMfw+x1fUW+ulYABWu+6O49
YAKD5Xg3OqECuwCTPXZhRydJ7FxAPxCZUJIvffESZ8czdk4UhNSuuzdvjKJoyRV0MXLI7VbX6K4F
+UxmgMKROdh5SydzB7NGLr4GjC4CPcXiBljivpdGOoxW/BSfn5KblhmQQLH2aBZv4PH4gvLJtGZs
URe95P0PnbOcynZQiQyecmPJ7e34rQGDj3ILc1yFLptfYaurVMGPO4T8Z2UOHkNpH8eCYBz6RoND
4tWD0GhNe1NBfW1RUE6XYA/VJvGFX1U0wqZg4BiYScxzbJcjX63gO1745evP91v27KHmL3Lx4M3I
d/ysdSHgsW7r8nNTeFM3hBmSmQtaHKJD7YbyLOq3S8r27x8IGxFOu/l3yFN80vZ1hvFDTmnPhq1w
omx2pTy/WThVHkW4/3LtAI8Pv5rHksNH/VPaUutEYUdNxR4o8bSnk34DQEwvc1EHMZ9hhmTLujHj
2U6HU3uEcL1zWoPoasETQxaD4gB/7dXwf7HRNSjIEWkwoEat4EuveOgpPKDMhDcHFiV0xPhHZwq7
hfzu6SowSxxJL5jvVpGNXud6M+VGKqEsrVCHmrd0hXCr73/TvrYsBEevTuti16K34yNfJCFVQDLI
1YrN0EnhXKjp/BApY/Da9pcaBkyY9GCgkz5cbNee9yWgErKy7rJzLXtieaXPLBcdMZL73CmxkBMe
qtCdAg577JGyMHid1DYVFrE15etAKvnp8z9BKL75tNNw2uvLp/GMEVDS2PB19TDyfnleecCqtND2
yaTG+BHJWRzoiVmSz9Gs0+L4GmPPmXkM8IzjkJiJuY3K500/egIg9VAAehq5zSeY7z7xMcpVrvmE
m99XAf3gctByyYXSlKXcHlYd0M8YT9tMScafsVwwuLlqprlI45QWWQrBGou/761xOKgKVUkof8Jm
BZod4fjEAboojarRygSBthRw9TSLd2fDK9ZNhyvHofS5Gn506OpUJPpGbBPEstFltnSzSrvM7F19
C3UQeS5poqYBqXP8znch5TDgda93Ixky9N+cv07HU972BZOxRgkNel6Un5j6aSe1VeFGP8aSAR0M
puabc1WXdkP4Fh1JLmqkWwWzMvcDxjR8dddsgYngxTiN+XBCf1oQH8Zfrlm0DiiYVU7mWCCa+nmp
GbylEFJAC0tzI/Z2a4IFjpQJgWySlYb8bCjDCXO+XrXcKKFCZvlyHHb1io0Q4Ib3TL72kV3EFNE8
abaTxkMLuFagn0g0I0pR0dcsrpjrvPiwLyBHUZl7PKyYwi563VKPWppV0tOgrpPRhORS2Ol6nvu2
MeR/OaapdKjWYUFWABw26ffLXx0KZY97KCA+Zy42UfUfNjs1YU3YUin3UCRmmKf+trWhrIHNN95Q
l/pcPMKYsclJSudnKE3yk8olbaBaiXJa/lGjMROlpd8s0NCcc1tCyoWT3lhAhTONYcRWnEpnyP4b
hZs3cN4BgXJuCRjEB7/gnINB6wg8n1/EGQWEcwgNdnOZlX2zRBA1qxcFKYz6+kkCdWqhals3OC9R
UtER5EA1HkGF5TwiHWgeAmD0l/DhsCFSfp4phjIpXfXyzZiBo62f73yE0KxlWGHGxreruqYRScfI
JQMh6JEN86rVoI1kaHD6fXDqZbflgG0EsbyHWznflN/dJINYkb78AJY+M0BzmQC8mPzKYfr4GVVO
Xxr/WEPTsBGa/epRC9yV77loKZNM4OHc+kmsTYJSTKa2eRWztyfzovEME8u+HfPsCS52oGDnoFd5
Lx8jQTzsTWhWvNOoG81XfVz7qag6CMxaf8VKyWbUAOafjYsq4D4WAqH+lkZto45jIugCweBrBqUA
B6xtSUEKOnCkvAFpivO4LmSerN0bTYXcpDNr9Ml11VIzftPPxc84fVibzepvTrlOxqYFOUI0CVxE
9HmhAaw9yvqcSDlXJbI7uAo1X2PGRJ+eTMf5I4Fpix7+BJOYsovTPR1D9OmhCzuxyG9pmdovuNsP
5M5oln3RvehmNnmWPWG+Yqh7g88kUo570BRy9zxB2pTaW/76A9A/LPcKLMaU3dW3f1Q2X+is7EEU
P5gyAIoIdx0OKhJ9EM0bj4nhLOBK1nNESvrHHD/UVn3QxghFU6ThJIB5Oc8WE6dTwgOYCDKQSIES
kLPIkgpgBARRTgDBGXjFk23lTDzMLMGlkAoI0BQDHpiEPJLdMXFmOpnjjPfSn5OPd2W4Kmxv17dP
y8FVXjrv8DK7ASalw+JwhfpxhuHmBYdVpEidEKEzMn5R8Y7r0KukDs6HoDQCqnAbep0HWkbO23l0
vYDcEIiNm6hocP4zPa09AM/HB5zDBAmaApivsqcU5B5U9XRKdgLCE8Y6Y8G5wJjQ0MCOjOUviXMP
m1fq7W0NGBuHzsSRtg/omM4edkfzqT2VZqhvWRjc2dtOL6nleYaT65vLfjFZLCPJewIaNkpJcxEQ
yInCLWq2kUmwjCogdRuyAEQAe1hVLZuMRQxviXHFJA8P6wZkT8FCSTft8RjKHCGECcg9ZSgeqHsU
a+gJVHc/l8T2C0MkE/Rt2sj/pNyO5m+aRjartk3PeKGILu1+rhW/T8sOB8sV2LMuyyV35h2yc+Az
t2muh7UmE+GXDohRX6FDoE2wZ8ykyK5jV6wZdU+C5mrhjHizCTs5jSrvWc/XtY3lshDMrz2GiFar
BhWiPW5jmT3iq8oHQEfBqewmfmTH5VAnsqC1TAm+2eCeFdQ9E3egJsqtG8ID+3LSFtVJQFwhFGvu
1rOJBC0pFwXU9S21iqyidKW8U/SI1bhsJXgnzB/HNkLJUdJId0WkSjFLDd9JS+B4mRPJ9jGZgYqf
7jK7Um3Kpg2yNGdkQ9Lbb78JeaB2LvqVSU/vzsYElRnbuKhLDYefg876LDF4YbLUSFUuPDXH4Xg4
xAlQFosKWaJMWLLL5SqB/Zu7whxb3cgXtL+Ae9/+Z/AAp97jLcjYAqkyathB+ihtdz7dansHaBEO
5wPJ4r0VK5Yr+hUowBkn6LDL82acri1E0LcN7OaBCVAM8KmVB/OfdolT/LpDFiOLEFo71ptXG9+W
eBnzsq0mP6mipyL1YzRAEKAJoJmbwUVFfzzCXU57gIdubiAtmK9U7+2SQD28KFY7YIntB8u7lB1/
BmxssFeuz7zB7SsDZgkzPU8UT35SvqDaw4SDyndh/rh2MI0JzzMAE7y9ALFchvZUOGzw4qcH4LBo
K8a/KXpVkVaZuYx1NYIwJl3+zO3PxUgGPOu8oF/zJJNFHnHkqZn2odo1viT7cJKTy0eK8/40C9ca
KxElr8nkn7oZSj0Oe3KOmIJH/kMEgdvwXDP+X6GLTHkSYDooszb3lYzIsnVlSuVSHnzXQ62EHPsI
ZIPbQAS7zX51SdpTL22igavNsilq1HrtJRek5vhY7JNLMKV2kvRkrsIMKXmHGK2eIv6lQoFD9i8l
p96zS87138OLnqI3d8WtRUq3heB57yihs/dn4EOUgu9ngmVs0gsaLwEMDAu2TY6cqMSjBViM1IOp
Y7No0L/XqPIah9DuHwWyrg9S9JjaUkKLz2cQg33yYdVRDl2KJlDCmPtOuCL+o5jyNNaVF42YG5P4
gF/lAuOlwqqKvu+/bsnEQFJbOE/+HXmI7jsvjq9eb2108Yr2vzLc15ccVKAMG99FhkCjST2R3RsO
ROqJBlov0Nbn9CpZgCrxEB0aJ/wcFEbzLJSga1vOSbAJLV+aFB+uY4oIjcQMX9WJheCigDLV1y70
ouQCfcFM/ADutf7zMyeSUpudA7DHHYCVP9FMaSYXC+cw3mvC1ccg6w9qg9LSnWUmIG1L/Ji2FyKd
KsMFxzc3y6Tu99jWKyaYIzPK+Y6kZViRuTpuP4pZh56jg5N7y9blXQAFQeWgZC91hzx36T1IGePo
mNJsR8eKd2l6Ax8tNEBlzvkkM8ouJY6qVGiu2Frgh10g4zZlq59tdp5mlls6w42IZsms4m9L1rvA
mWD48mTluj2sYZsGH1V8T5oTTaulKfHcfMK8D852tfG3yuI27qqVGrUwT2WIgbFjH2lEABaUs6/3
aHLzBfeqgsvec2qkf3VJNMG9byZl6EdHJSYI1Fu910XgstEg/CIAGRQTI4XWuEn/TGX1xYQy3WY8
l7KwA2jZjHNrnqg5xRpIR5SFnRDS0A+ObUuzmF6QuR1+dNnqQF89rXfPkBV3rGvfnfsrCyg6ZXva
oTOrq6sJLd/8wWrJij2/kI9JZ+X6zTWsgrJ/CTOME5v7yx2CWhE+CjBnw5h04+j1Q82zlZ8lftIS
M38PztD3kA7T60NRwEr8oScVkLSeLaUdn07OSYov9P7JxiZeCbx/fBFgBYzZzb7IkbvQJ0RM2/S+
Fu4nrqTXeh5DBXPuVnhgFUvUMdQnOy6ZNbivwyBWpgXYNrYodrwiZxqyz3ie43ZgA/cW/yTb45nZ
6O2zmzjjXfws8g3zHMsVhYbijlHgw5d7+PCEDx6C6rUVEQ234hpGn5uOU8Tz6dsTcTI6BvOPLZe6
jmXv9NSovitsxAp0Swq779BUsmlGEN3G7rtnoMlIom8WcnJonYzwm0770WBcdpBVBAS6V6TstuMk
rohk9zNnu20X5B+ccT7p4pVr8GgzXUFFn9UzFmAGn1yH+oTr6WqosEfxdMv5gsSrhCPInzpOD1Qy
l/iH/RiXcNdyybWhEPK+hdJluDJNqTeZD8QO/zW/63cwhV6ShhvewHIO9IQQTO5zRu6x6jqcZdoY
lZMj7KQg9juPdFAeiR0iz3uy8UM2k1KCZ056FL2Mtg62jISsfcx6MCIrIuvaunw6teK/qK5BPl5S
/thOuiDaHYUqv7B1ztj7ftvPNQoiHJ3emJYlu38BAFa/w6Bn7elH6zksi+RezdmKhBrQNyt2ENXB
JUA45MynTEzWHuL8HLDw81SslYvp/6l4T2/7jnGMFtatzBLiB0x4RgKq0whXxpYErmQzJB4o+YHW
8kXsjESNsAKlwoTZZM72FPA9VQTUi618dc05Jwzt8a5hOad3ThOWMbrId6TbhnVlaLUuE+xSrdyS
OOPMnYEb16XBOFroZuUQ8k6YP6ucF0a1v9+abTUK3q79sMnX4NjaVAY9inOFAx9pXJKwriQdFs4i
wQHxSW3m75tB5mFo0FXEWmB7iIdemzaEagy9DrxirW86HEiOMPu/aiTtaWApV8ReCteygOkk1b2E
mTP3sQaq6Fr50+7b49HaH7ftx5rahUjW0XYuz+eJvlljgJcLRWQAFbSqV8d2Xn6Qxy3mypBF3+ds
a8QvrgdbMUX+VeINjHwsTDyx2YNw5dUhCeFza8zac4eSp1rhp0PUESNb0ae2pnQagu8SRKvWOshC
n8yehk6s1X14wwqeY8c+nUH6BZB3+YyICUwzYLY+6dGFqLMKeK2vklCBdC4r8Aj6m+lS4ixeNA9S
toihwRl5MvKVBcJBCxAEZtecAR2ctXA6PkaXqx3x6xS+37kRL1vrVSpPjmsrZ4oIfTrh9UvvPfHR
uIVCJoCTTJVb0cD1Vmn7mPgzew96uIA48fGmhd7WMOQCkU8PWIGdLLxr1tMaFOKLhbh1QQ+qAUPz
XLxZ2soJqSpowYTOVMZ2TWmrhmVv5yqDm4OW1BGoa1KF6LeOzMyMNHdVfxrbEjADZBi/rlsuUd4m
apig5SyPoSIvQwdSPzQssi+yo2J/HA6hS78RTarSkW9anPSuB7UYL3KJQmVilbIZ6RXU6McVW+GH
q1IRYQltw18oDiJRJrRxW4nzEfXZcpgzpkWRz9ie/67j836YysM9bUI8zh9U4N+3RpngKw4Jb7cZ
pSGB7Tsk5AoSSelitP+N0h5rPJ+tkAjIdJYheTyFsF2T6/FmdRFmwxCzIEifuPZE//YMSAXiSM9K
FjWXEQHn15XXlZnwo2icDwytgGlOH7hoT0BrJszqX3ZwnA1L6isbFZYqabqkb5cdK+gnXpyHzHdh
OMIEy2lN7OrCH5eEwVgMsQV4WPBbLAfRi5lG937ie7qetgEkfOOcbfyIxBusHTA6MbxcBMidvTwe
F7n0w28fEdg+SnATDLM7MRIvbxtB1j366FjJZaMk39dPsusaCnF9rrkC3GGC89JS5CNEFLGKv/8/
ds95mkOEFLQ3VslkCfjb0/pQ5D/VzefVch8d+fR6kUyiN6VF3cZyWGuz3CfYuGcjFyWL1CQypYWR
bnvvvun2NJ/QSTKDwyGDmoPnijOgsXjf8LV6VHDURivGk6ip2fMTmvFRK1uPkZqvL/R22CRV1ORN
gCbXrL96yheRMamKkt6ZSTDMgWZXxKR0xl3C0U0jqBX9bQjlt3pjz9hWHAPOJX1DQPqZCJwoLGJd
gZ9SeNLuB5dJH4/zTS4qldavnWNgsmaUSK2gRzjLjH5a9ZbhQBQrZMt0eYHYJKvw79V6l4tmnyg5
3m/Q6VeSg9GJ/G3m//BEWyUFajOPlGztBiFgTykisbIAWhCXBHtBaJfSiPTJIkKZ5ufsF5l4GLm1
raZc1Tg9am3xfhkDs78RcHR2HOrPt9+6Dnyz7JkjZdFU7AvF8HjVPoIrr5ZVG6XxlCk2GSrzLTwp
owwGfIFbt8M7lZ3mH2dzXq+o+QprmhH60nOuxMlLTborVkO4C1p2HUeNdQIbx9s/FXvV/o31883/
kdRZFnpqSPMZHhYEUlMpnqq287kLNvh9RtSfFtjudKsfm9/t0IW2aeA8dP/Le1pUMut5j1OLxSO7
2Tw1evJ3GaqPf/of1/vcxKOtOajImCCR0ARzrDHxm+jghDumqxG75XKen6Xkt3V5t+bprdHQg312
S7y+eciiu0MWw2Wj2Usu5nxyDMJ7rJTRJeIUXwqNfHBM+PX2y4RLbBVGYmr2KfkFN/+fJcEmzWsi
fYHvrz7TNj4C16bCla2bYqLqd+1+NQU7UtQq7p2soM9HWjhbzVHUNxloTpz6gc0Zr5GMw56byi9E
+eshu0uo4qx4edcPPyel9DjTxkzQKt5dCpU0tP/yBPIMcAAMT5xERvv6mlICSQlvMObKwfY0ek6m
cepuDPRvK92qk9d1WKHv9YUUPmbZeTLY6F9Nle63y2gXBvoSFza8w4d5tZV+AppPCxUR0gBUqttR
U26UNIiVdibftEhIcNb4TEf3enx5c/M5qjo54geNv0/W7My789/lTlt0cCdXBpITLFTec5C+2VkP
E2lLJT1voqGFjqwh3jg6qgF2MXf9ui5mMMyf//j7KcCdxG1YMBILWweQ9SohJfl5UWZS0Bfbzqqw
BCRqDnup8UvU0Gtm2dQ5BOvCjYIi7bVZ6LXplW0fxZyem8V9NWadMTqjjAafNvUKf7JQFEm97lyy
BL9X83m35aE6MwvLgdwM//Bmo2eA/8BOB4mB3sXdd1zHGPFwYCo/gCA8wuzl9/p6PmZ5DgWhx0pX
gI3NgYsb1dJRwD7wgBGCiE8T4X79zneRzfjGGDZwe+Zf7Aq11tmy1eX4h0LzhmPBDKJvKnRDDrKg
rzXuL6gIlf8KXiecaowyRba/Df0FYXk+YWMAnRX5h3FoqAH5DTpJxHdWBZz8OUSUpAL7Cn1PDd06
9TmFq2zi83n+MPoYQU+YPTWtDWEJz/POmRz9GxKOVcSlZfIMDZ/AFEKYoG1QsZNVJECasT0zD6ur
WcfaYLXnrnuA8zu/xAQq2CQmjnBIqE6K3g/KcwD+j9cb2VF7SBlakbFgYHzTyjF7fZyYZVL+hZOq
UJAnh4vjt/hNm8Ux+MaNY+fB/kuGR0xkHj2ruxFTJ5trcMTMDhVbgvme4tJnX1VFZPn/coivsIGz
5yKIYaVGBVslRyr9AHr6WK7cqd95kpDS6rJIj9gxZoY6Fi/lheun+2FEUsLIDJzifzlJtktjqqS0
v93hWlhhNDZTNK9ACRSxmR2xJTD7Z+JW6yMBIJMujlAtNSfVuH/sN71s3KFGdjuQHX9Sua0YGYCp
+mnnPZAfQrVObPhaJEx9bPgIn0/1J31poGiyiCa6wc0Nxp5CEPqyO9QNyQEWVT/9Jr+R1nXvH15h
7peLEdnUS19aYK4MGumn+hDRHq28ZirWr7xrUoKhZqC+Q/cqhR7qsN291w+smAKAbS7wVIbma3zF
DMS4AroaHgwP9vBTFefFL6nXKQE/bGycR4b5mwimQi1wyjR+scfXKd80oFm3BArGd84INva4o6rs
ZFOqF2ANK+gFsXs3uPRAwmrO2YMcp0Kpp9rVTY53M7ypDrKYFfRSNkvnrAcqNgJw2lFkYvS+MuO1
MUbDzvQiHEfiU6jpBOOogNrzdcflN1OfJKZba7TIpasVL6ObzHuj4GUfyLZIdHH+kTQ1kIn7mVJU
mEBap4aO5Z/gbCBwCUSIhgbST+L58mcPcPY1yGAURTl0Egb8hhVWIaJx5mdSDCX0fktRcow6SDXL
uB6uU42rKZClFAmzrf3fKBch/laQgbEX+NAnMNzHbVWBXhDaQnBhtZ3oY3pCI6dZ+D2+V5Rn5pDw
DUJ/j8fX3zv5zOclChgree8LcUgiKkSKnIKLHZasibXYZYZ9O2YCEpipWG8UP6UuiOhhNqfDc1tO
40QO9siFlBUbsoZKsoOXgIcnIML9ISRTaZbNxQYJr5dLKfCPDUHG7bs9UAeDjJ/FityYONK6jjB6
FhZcySm0oKdth1DM0e4Cb45R6ptnAlCduFmQsfkQcV8xPEDImujnVRdb0Bv0rNB/NpRqd95r2TQC
aVW0/Ny2tSYFGSxVEQrScVP5d+XMOfv6mCpZCo2T8R5MW4nrwKP8Dy09H33moB6qlj56TyRWuaI2
jR42iMAQeCAEYjholdDL+bsNKhVIUaC/AEWM+WJX5j96M79WiKhJ4kuS/qEwH2PbYsLGi1n+sNHC
pkzQXJS6w9tEQb9GzRGcdEaNjbEvPPmXAvU86utSBgv5bMpHivrbRwrdER6+H6Onne/LOCZM6t4i
W8UX8VUi5U1bvLxmZRK8p4V2xPBBdyTohxO3zSZ58ckX2qID0u3d2YrmpoBiQIByKVEs6+OQCJZl
KPK/UNNKKHOwgebz820I8SmS20jErV4W/HEE6QJkcKSJHEUVCZ3EdroJ1HezZEJ5pGfHethI4C5H
WAmm06s/C9k5eeTlDJMCbz+PIO8++kL2h19pDODuuRw8Inz5Z+XmQ+1wmvlHgUffT/efkaiA8ECH
/M8c7LDtPpTGqW1uE0tf0lu0kGNT4L9tmFKKfvTPz9n4fjoKCh4CNFCLnTG1qOv00KEbbCI57XzK
9sfea9Cbxqyx7qzjKzD+52fsnSAB9AvIJXpTL3j5V7zcgP4vU9b7iWY6EXP1hUgxNBDGPUqXye0K
q4LBrRQnRpRS8tcZUVngb8ocfGJSu/UqcJ74T6SdjWqYFf2eWPS5VIs5Jq/SBB7oR7NaGc5CRu6T
iwmF37J395Rtmn2iW6GUQ3kwVhNOhlJy4NXxXX5jTvDze9vbPbzRNftUwridyBm8wOES5OkJcEe4
jIePd/AbAJPlsssVam6zyslxBd/6vm4xqF/helfBwnT8tcK9LUOUzCoeQcR0gFcwY/PNFkWKrar5
vj0pJdxjrtYJlUPRn9M/UtNHTG3X6imBoGHPLz0n3hyovrrULu1dEyRg1UMP/vvli/97YSAXBz+N
7jlMbBA7UAv1bNirAbPXqaBrP+a3VkOs2j5+nTPYzI9ECo9NikgG5+p8cfTdu0VtJlu8A0Gl52xH
vpIho47CeEAOBKVChJ7JGGnoCAzonMSh3yEAEU9TmedqVJwvtYJZ946H2ihA9HmdZtlYMpy8yE/8
tEToS5ni4QxEHaXdyTCqDCOsdouaG6f98hK6Rr6f8AcnUL0/L+f+98WCutAG+3arK6mY824lYQVX
ivspqvSe89SZAujn6RprkI1knwIv4UTit8tE63Imolewp+K86AYRmfCRZRGqYARWgsUHcBgbbzbw
9VhF7fUaAKk35638A902+Pj+oFOaQ2vJig3HPtQr9A3q1wZKbZb+xwSv52OaiDkBJQZC0Gl/SKyb
XbEEbbiJoPVcnZIFadpxCEWY7KzWX5t7XNoXTA8rwrC30LdtnvSW8pEvoUekhCSWWkC8NIEuHsGe
TrFdww96NHRgE3H4Yq5/1jeV8BxMWY2qSjwBUd4mZbAWnGaGu71XVghZCKTWUym2oNho7C67T7WQ
V3uzykFBtqJn8xb3ECSyfYOUJNlYVNxWGJr1B8LJtAIe2rY1ap7dsRm+BmpnqEezc74OhYiAAL93
5uFbDfitbzETB4DRuw+8aH1S66k6qEcFOzvPCCRoTq8IcbK8D6e5WSxsiwDxwt4DoVUFBh7bUqaK
khb3RhGz5GaEO5EjrYaR3tg5LtIOthyY5ZitBledVbyh6Y9laVu4Scp6l+beb9nMdafBvMeRtIK6
yf8IU4oBHjmW9APCPxcFQuTYNIMUF2Z9Kim/8P4YjbpBytWjNzXstVWPUmIgYrkfjztFvEgZJdRX
bMaFSQV9bwlz3EFtu51KhYVE/E4BuNgcz+xYkKwIZDj9lWwhzu69eLZVtx1EDxw1UqyfKITFWrNM
GM/kiufA+BvVDc9QvCEOHRPpId7UkZRRpVr+9tYpvkP+OOIcX3t01FczIdQUzLe3YbitsShFFmK7
hC3HCaS5bUBJPBmxxu2pfHd9THErtzuv0w3UtDYG6hdEURFRWsbx4tB3uFNuyXDsEqpk0FyRx37N
yRzBdiKAhQhNHFrRn4p0oyh5VE+7wc6YKNa1lqrI+K7QVzqgthynVE3UejNjvU9nB1MkLXJP6ey6
yqnfaPomYj46Bhzn5s9RKMY2vt4yHOeEu4q1CdbE+LjK8pJxYz0DZHCKe8/AEXpM6wbAS2ixIsjK
IW9LDR+Gv+UuiyfJfoIQlPnemYskidgsFK/xGHTxr8nFdwmD+BBSZhzy9VqdGxkPjLiOU2b7RMeQ
TtyXuacJsZwvU1C1swDi55lrYO0Sjkk+5eR/qVQ6UVN+X1vyv+raS9V1XrITYbHYFnDUpAQ8zIQb
c7eds+GrM5nZwLNLXqwt+5kwm5dbtOJo/S072ntLe15xSkeNmLbwCVAlPqGFuCAk/fjClIMA/+/n
3dpFccwAYsOgh/oGAYtYsaAb+IIh3YlRX8h5T/kYEuRYZZuK4EAXfjs6q/3+d0MGdGxPzDZMicKZ
P5OrWuhzBX5f3IeZQEriWSFHmh5aW6DHQ05Kyfw7F14DZNRC/yQ2OePE7onuhobVdjsHIAJCWfEp
rndUIF3L7II1gKec0WcYVwHohTqEIlb33VbL1Nv/yO0MlXV3H8EWCP/K+6FoMXAqsRAR9QnZUUPx
8wOvly6Dbkt3FJB8UTEqaI52OE/h68hK+FYZEH3K7g59O9KDxq2aa4SV5mqcbIqRmpnSu/z5ylJb
uWRtZCqf/DIsr0eGDF5VruWYOIJOIl9tr0ov673gn+4fLEl6EtXghH1wBwxCIJtMVWRz/1QaPyI0
iFsz8VFbksJGqIHDXJLX+5ZuoyoklLwQGj4iQQaZYjA8ckw2sSNjrjerWo9CM+8p9z3x6BKqm1aU
+p3Plk3ZoNYeeI9/9NRhC+z8x29dDL2KVjJ1BnO12G8vjTrq8P2W7fG+nLRGlpXuuosTsxv5FbEl
Izp2LJp1BBESV77LEIlF9we9TlYAJ32Hwbg5hLydC1B3MaBRtODR15tjnFfqYpG4sOvIjv5RYd+D
1cDflRc1/Pug7NEU4TONuc8kqJbVaXt5DZwcAO0DXPGejviMFz1e6YOtJz2V2XXBzAFwLStFFXah
lk87oQPs8HWozub8EjvnIk13J6V9VysE4qYQvodKDPgMSdQpNgMW3we/+hSbxmMceyuSEXxOmIXp
vxBIlb7j0fLaWEyOPxMbxa9RQ1KbiKZwPxXGq4k3ye9/C9XJfO79lLz7JH19VynjWdHKDKOe1S4Q
Oqip6GDmHq3apoNRu3r/z8gmegv34QvmDMLdXg1Lhhyu9qDcDvaWn+ASYKnENBajKGlqwBOcBGZ3
kjPVhi/tztQ/mGw4MpXbL4RIH24c0O8cet1HKSKFOClcsLm1ZwUn4EcOcfOAA7uCPWMfwMJ9iDRC
xv1+LWYWMM4a5MC3Zh/O5551w8NHKyaDbi2onprjlfUaJF0qdya99hwty21WY51ZQARI5t4UyXLn
pyzVvBy0104bpKCexqn59kcvAmxNOPQ80281tZdnwV7QK91PLTM4wx403ivJr+wvxFteO5mUo+Nt
uT7Ag/sT7GV1aHogWYI13J38UDZ4xTflaluR678eHt9qyqHYVVutXd3q4/4hah845a3UmtCchWHw
v1cn0JpdiZlqq98sXURINJxE4iq06GLQYY2keLNxx7uHQnHzMCLPn5SE8ufWE1sfkxAKVKMCHu1o
LyH5esf/RX7neshvmb0l4eaYesKNIVy2UcQNilryLIZg4KWWjhxfMxt+ueeDm94VT4Um6rrqf2Uc
22gQek8A+OVlPSgZFIamOZmQpDgChxvZdQX9B96UY8QMqDs1cpmg65krolhxuTVvFJhk2CESMhBF
PD6cqFpHJa70XThOHlC4dgIcTbC/kE+z212hPTtbjo4Rv57Neb0m+bBNDgKydrQWSbToaTpPbMD7
H0Z4kC+MneRCGejkb7BE2ngUiXYkEPUNShqSS9Zi2Gg3L5LNiMdbPC8TneV6sqnsCqI8t6JbpuxZ
wvo9oaYww/+01ekmERuJsMoLEZRKphHIB/F0LqGCRgYv7Wjme0/U+i15nsYtBlGyJ+7Ph0bz/Ont
hFD+NZeeQs3FG7w7kZwTyxpr4+laf6Xywu8OHFo6eAurcjB94ap7wzo5PNHSGj4nUDsaq2MESAOA
3rkh11tFrIbonglKko9p63S6PneE5gArpyVqngeiQCdF+h7oONue0MJ/TAzJczoggJcsbi6zH8e6
cUeN6xjv6DIr1JgoIY0pdSHBKoN0TaOtV9WIR7Y0SWmlPZRz+B7oj0ALagGe7G3LUb9erg1zlFHz
A1AgvlhKKbZCmgTMzR9msH+X1hwy+zo3bOiVXG+iZH5hO+LQRVzgjBe0XQkrevpPMDNopphTiusz
ZLjUC6kDj1kUiidoLJKryqS8P1+ckcRP5Nn7F1ZLXHo+WgwssrPhNKQ6xkkfuPS8MkjGcWlULtIo
2BvuPLhxNUjWb+++J5JJWZCiwuuTKRTwSmUgtY8qsYhmuGKTjAq6TUPdY30p4IxD7hvbAhMtbrkK
yLjtGOrhOCmbVtecmlavr9rX3HdLzPs7fNO1J1H5BTab/JZhpzWYBcaxeVKFUooZTBtYavIf9ktO
cttSBAeavddsvpVqOGZab1u5nAJOT+2FsnGrbLZPq+0hwes2gyQwVaKOb097SKU3PXkgGWqs39bv
oTDGw8H3DsAN4Id2fhj1+v+PelFjaa+rJKoz5hCJ256XOLoWhP54yywEiVfEHseN3jp7KHAxHOWn
/Y05iKmRdxWFsZPT/EyRitZd1IERtj54ebUgomva5bGZBzg/d6r0E6EleSuk0XHgqA2Tff8VfAly
c1c4zDXLZHcZAa1cYwsDIcn0nGKRCRMwqvhD4u9VtrEBhbHqHEa/Yt1a+1z2J+KTJXobOSD2G/Dd
FpuWERl5xPkexgRXU942jZanDRZ54VzY87p5USLzBSGDn4ZGMWICQIooGEs4Fk4qpowEWCul/HkG
4LzjSOjkySoSQ2xX/Z1C934Dwhv+WTAkQb3iV03HIfWjbmvSzoHow8Yh223S2FcWFhaNZv2HxuqC
CdbXbkZjZleyJAemf+A9qU+P8vCDII33maxVgVsX0rWVjHT3MIwLx8wUF3tfeVbigMA036n/k7gR
v78IBK/XHWKa/79ecb5s9MELULZGDtv4bGxmR+Fy5GTTXHwIF2euAloQunrqVZbJ0UQJuS6CpKnr
uCrl+ZqGjKS92L8g4xC7X4MJm+YfmZ218pE1NPMLKaxsCUV2er0TteiiRlciw8aP+fHKYCmlVNSx
6S0d40ms6B7ykrIsiQx6NZAdbl9JfQNbY8QJMcckrNHDScmSP2Pn5k+PYim5MHIAd6dS2QBa0Apg
OzRHpweT9HXKT3CaVuBcbuMGBbVo8LjXcSUbMf5mEzh8cb43J8iaS7D1ffrDmhEGIzeXqw/7MSWp
N6BmwkhvD/H+NaiE08CHWQ+OGeG7ZawXSJ9tLOlfiyin6zat6ZPJwc3dMfMHIdGlSHTqcm5BZP+w
dpZgwbqYnDvRez6EbaoRxJilqsC4N0ir/iK7/CSJpRpHDpETsa2KPrs2Oi0yMWLBVbAlAXSuSmmD
KfGLA49Ph1nj9lhXfd9oLxNblnp2f3il55xJGTIJWG1uZ4TVCLgNSEbB63ePVgcYnPKAvYj6SHY2
4A+2Vla1L6hbRWXLQ78VoWkhog1VnsbDYH1+QIye1zeGIrIvFQI9s+txHTiubTF725xfFCieYEpu
VgHxQKD00deQK9Qn5JmpCG5c7eL10sTqkzGh+JeiZoxFgiQ5lE6PBjnf4uyLM7+0/4S14Kqkiu2p
ZdOnma8l290dt2NChi7MoEMebf1vmNZvJNWcdI9mIitqZ0aJcNjf2HHQLR0xp7Mok9LEHDGhE14O
MWzT5G9JKYneaOVn+NDt1OBkB+3hAk0ol3hcnMBbdXiYM7yqgQLaoaTfuqw/fxZcBJFCT6bzFGo0
xkVSxma6iXjpEcS4Qigt0OC2gvudz3Z/7VL3WkiFqEILzHHguEEpKV6mMM1gLNvMU49aolrSRUE4
vVM9fEPmhNiZWSls6pX8CZuzfuKf0x27sOjQR8p7/EOr9fBiU4IgMYL9Ijw0w4rKwKxB6o23B+kN
j25PwJLlVnPzK6YXNR6qGNmZYJeVCNZTPR6IX8uBsbtzm9L8Oog8M6UU6fMufR6nf19ePBFSzjhb
d6b1NpmVWV8I+6dGC6oyc8WeQhqhdOEOQdpcYqhhTIUuw0Pjxf3KzVHOcB/P44Ddwv7IpSFkEY44
k2lZHIo0Sq/qJixh3/uLF6QQcN9mCPjHDb8O4sY84vw2IMZi0CdZ+8zGhYJ4wP4ALcLbPo2gJlqp
vBx87itLrJngUrfXuhm9DhZJxqDRZGrTZii9bSuk8TeazymgcyvCqZcYPixXqa3qCFB/KHR7A8AW
F+lT+hzIVmYK6/PgSHE+ZuuRsOoqpUsZ0l9RgRzaLopK7JVNZyX3nYW9DThJ17fcfFQaP7L5C+Du
bP3gU8OOsa/mrlOl3+ULqxLBZvDZeGnvXcSyOEdbNq4IcUXffKLWPzo9OnUgDxTM/aqeP7YtIw9i
FtVysyDBMet9guxmU71GagzwjW3P1ABEdm/yjLL6WJllxCeWQABuWMePjzgIj32mT/Je24naxcVZ
eu2Gmv1sAHFuQQXjjFOfraceMINcP90yDW8CyZnmgaigA2M0Ghr1qXu4IeScj3qJeqJvP7cV+NGx
S7sIuHIQDMc2bA2UAAoEzX0x5+W/UbU6pPTTioI+mn4qJfejdXUysbPvq5O6HvzRtpt6rumWLz81
R6uGXhml/t0NHJE0kBXxMXy7i7X+albnFq/BCH4brSslc4dOJrmYO6PAprRdpaI+TJJ/OOLEAqyw
pno5+XAXh2n0MT8IuWKxBrTvBksPH5u75/rR+jhQe8113GOrkjHcKdAvgB4p231YamriPsy+roA9
0tLYcFD8DdFtzkjK+3xixbpNHw/idU8MA7ylzbXbg9LYAEPMVuZgzGYqR8hEEbGdy+T4ZcmaQ0XR
olxKynMpUn/x4Decm+4UjC+t5sfxYrB8Py+UZZvHnu0wpTDUG/pA6/H48EUmxK6+hZiSSTI4m9dH
9OCl9sDFdz3a5DfEIBwC6TcTTAWbzyH4a9gRNMyxqTS5C4uBVR1iyaEhQHq8fn5tgfZk6X4XEwhG
ARgb9Un6tym/XHZDCpbuF2/gRltDkuT/CVmakYo4nulFcECxV6K33g5PzWj4z7lPlOMTCM4PvFS9
rCyqo/L0qYLrnY6okXiOcwkSoofC8xRPuNe1cIOwLcoI/xy+JkKyGuNdThd1pVm/SYzcyZRyFLbU
5EZ5CMAhLYENvVfQmHX0BKXwFXDK7uV6zBdLva6FJlk9l7kPRgPCF1RTWd+sPKPcmPd766YGKLqB
g9taJoxyBuhiRXYnWYQKidR3ofB+DyY/CQrCk1DhCyxcLpuDN3TrfHQj64F9CrCox0c1UUhyjNSE
/hs9wmwqxI6gbdgMESfjXJam42ZsehiaSi4yJHVXUlUPIL936CCpvO2QtoOu9nvzbgeF9NSGCdH6
BPWgnfRe8T1XpkD+ui5G5Wc+WxhA0Ca8B+4iCGt3S5IMel3MI5kItfGyx9ZwxewQpQ0vZFva2MlO
YybqtfL2I1bPf/IDGAeHYacFnSHFPhx0skkzvfmXaELjUyGYTSB24M4S/4Gd95F3D71Q+F39AM5w
LHPfL5iu9cQLAPSGYgSlNvPih5s6XH2W3OpjhQAqeLsGL2NSk82lDZlFaBlha73aVO7kkNSDczWE
F2I490rZROFT+eQWEiJ5Qbj1mayIg8MxZZR8dELBKGEaWjKMq5O6ddvvjLMLETPS7b/uxoxGsvD9
K4yx3ADJSi2oeI9jwjDl8x5fQ49ivUwQhOfQUhApO4xJtL6sTwcgVF8R5tDF1iypVAvL9anCfqPA
SDs7Ge0pqJuJ4ZjD9L62yJ//hjRMolJndi93hMFYDtzKSN6CtQrQnhLhDWZUXzyiD2FaB7N8ip2p
JjcV81d8gxdhD/8PwgBiQAIWeBRoxQlmlbWX/M86XsojR03ZubjnpT4zjB0yofoqS2B7/ghNgMds
Yzs3adb7ksloxHDoFkk6RwnBf/DEL2cAK4CXvp2+JGFilw0ibBHRKAF4B5JIfvrOsIwcp+2xGqGE
wmK7qpUmV6c2sBYUFx5pOTSNeVHHnAvHnewPM6d+icyvrzbgp7muDePctfz2NjEzitINVf96WgLb
PnBwuWcrXRWJJ8ryi0OlkcjroA1ESF3fstsFoj37SHDYjLyB7tr2JOTsqlxqBCzSBn15NFQAPGXR
zWhzzmeI16m78ezJaBAyj2muQsgqefDaVDFwKtWTayNesIlbxHfMcwybJ2/iok3BzvLSmNsKQPpu
uwZJoyvaUKDlR0eGqgdBGwHnJn9qN1Sph6DwJS0SBiM88T6zj4Lht/WWCuqsTWoe0YYc93yMqD61
pB4os3aWwUgjpbzPpk2fPtECFLszms7W9TYLZIy/rE2JNBkZQN0iaDuks2r2UTrfUubc0tm8fUqH
S42Z/GneawEnhcqWVa5F/JyRVTc//vVd60RGFsOAGqPn4Dv1xmrSB1olvlQqx5reROcuMU1oKOSp
U5EXyy8VcnT0CNfM9mrumiCRWyq/LKPN1V5+ImKw3sRvZVzAjH5NysQUOO9TT4M+JziSfsQsBSLz
SpUn9UqsBajmTzoRDVYrQ9wDc+VHj+ic0PENHwkbs++z9hliX3ciLCMsJKzR9elUFxwwHFWoF5Ow
hkFSIaUWznyMhLt6+wHxU8d5uPkoOP+NShTnTM4QBd0+6wkYO6D02MNtM98xtXHv68eTRXksb2vD
Vrwr+2T9MiNN/Wsbn3BEFxFs+txNQvKwN5BwNlmEJ8/m1UTvPjPmtMk1NEQJoH+hHyA/gbR0UU+M
cQeUP/igjLTHbscZ6FJQLaLUgSpsDx/1ok7QSrNVV79vJ00X5YGJJeFq5oLtYIUA/p4t18dgP/cl
q6ihGOCfEK1+lBFsfFRmsAhxE6bF4NmS/8By5SPwPis5bZokrou9WQ9IFBoTTD7InW8XYaMs/qoG
z/Rrlzs9mILue0me1EhKyIMM7T6rqmGgQ2FSg7RDi5Lac413QczN5ba7EGs/ihH/IMpgsf3LL+6g
+bozoyC64Q1wdj9rS5HVFXoDJQvC4bc9wjrBL/4xO5XwLjsm+z8RyBBsbIVZzSqGOIFJJabjSfDO
ShhU500xDh4i05uLHAen0ZpWTYST57Vj5pa34HEE0oe/qiXPp7ypHANiuOxJmzh7zCgc6ztt42qw
HXCjr1nJAYN3MWKbS2sKmKJifSs+VhQVTem5SEfwwUA7L3MhwY6aYNUyWRiLeFWXdR5WTjXZm854
pu3gSW5sytT3rCkwCQbn8YoaWhhTkTtv0zRNiqnywySqbJIEbYZ6j8TZR4D4DVl0foL9AOifWOqP
a1zmkzmse+Jv90v8HwM/WHADUCN/Z2rWjZBFl2usk5ImkRINHykdyNDxA5KP4ylatl7+StYE0Jnr
bBNqlGy3PeeSZwvkHXPiztHW3zysfalfWxQFMmQRKyuGkNGqh3Tw2jCS0VaKbjXmPARqJZoHeH6V
QxCRMFlRG8dwCfHm78VXhKjtZsSDy1AUyI8tXYB8HmW4PiThoYdYomJUICq6Ur7NN8Okca4X1FKw
Z5DTXkK0IkGU8C2xX7TZV0S6lFeEei9yn/uZJfh1cRpoYKLuKACsvfwOyY2hCLaYSgbCwZFuFFjO
SOUAFQe4jTZ1TTs64b6ru4dLM1Iof0AUHyCW4OVKotR+u9XabRp25hg9Erw3SBSATVTk8NyahxiO
tyde3naAPGrLhKJm7F/XzoPYlylBt8xAPh/lypk6kCr+AxPzAshF+IKNGVthb/ZWBtBzVMQ5jHKx
+/prWxm77qOX7cUBh02FihEENSCCX3f3NraUzBzmfSy7vP27zBF+FF9GH4as3azHmblVJSMAc+Nu
qOrwXWx/lZu0c3kt9IgOygWgob3LMoJEcsMGlUQLjt4/qXRvJqsmGURmT9RDTdhHDGF6eTR5hPoQ
rpZUyDp1vsH628tygYqtJuB1NrTyIhfMEmNU2s3fsOSUQlYnQKnMP4VXh6Uejf8hf/73SBat6gkT
nRcOdUDuRB1TTttV99mr5vLd4aQDI4qUs037PyyErgIr7CsgWEaw0EkIhzZQzWV4CKFpR2h0xSOs
hzCrdtpEpoBSxbB7aAfl2zRXv34CLh4g/dq4qjjFXgnv01aM9e+e2e55oyAB08u5R5g1wfUb3/Tk
7zPHkipBTTH6TmGKn3+opJ1/JzN/txLFtQIbrVz/ut50UUYVmTdRR0uGzStXbQffyEGrMgrDIQTi
J/OXs7RJU7qrl6Lac6HftLb9bclIsAq1z5SjZVjBsKriQ7pQ+bsoAbhKLhTMJDd3NTqnu7QVJzWT
yG69bi3C9rq0pFmq1eH2zAjARRCJd4vLjsDMXz/kES4AQ6Ja2RduUBrp9Qcrgsj7fUof3btcsWUB
hXxA00OXhdA0aj0ypyorm1wPOsRLuZYjWoCq9cMosEzcbEStjDwR0QrBMjZ+BpM/YrCdGrKKPuL2
PrJEhR5OnmHEzwlgxtlYWH+T1j/K4HjdeHgY+f+6NB6K99lGdrAxghroVvbE/H4x5MJFYy2H6Jq/
zg30iFqSVh7yL4CFjrF9RDeJMCDrF2gvUfIAUYEXBZWBdv0eyuClX0m7D8JqMWYAlwkM++yLwesb
StHucdC4SAyngg6NbAEcn3D+HGevFN2xVabFCq9sSDDbsqiw7RgLKPFSoHF5gOXgCMEh/f3JGlcG
pqMoDZ9PzkFMsihyoTXyFqJkHkPr4zeaGKFIcsvIhgEmzl39sbi/3z7do0rh18V21HdokDzFGzmz
h8Mlei2SIgfzKusQWWjSf0J9DjCuhSQm8ChN+nQky8qwLak1a81LneE8+tp0B4eUyQ5y8GQV7pmg
Md9y0dthTJTfWFoIzAQct/TEB8gQUQFDHGSj8rnDBNowxjp2cWL74g3PVD/1Z1+p8J3ZdRFBDa7w
NAyyc4efP1nKXhb37dylcWllE0x+I9E+miRS4jtu82KSCcsgcHrnzlZdaXMTa9hKVUENWJWK+FJI
NOtluu7ZG7M+DJNDelNHQK/+hpZJLmYOStc6bg3jOVEcuQ//OzSvMhM3jg7252UVAvVB/4QYglq3
I6X+Kg12dTFifWwzYWY1DuRcvU4HyOLvkm//JMHAmvBG4vI9WwwRR9gHqfvKd2h4iuoIIN2HQUu1
0BhZ2rZn8687XIZroDUtYcG1w5TlprcGrs2CLyy7KwY48r7/jRyjS6UEruPqfT31vrcURX7oz+n0
pHcvgYYu+JhSJjr4wnUqeYpJwb79P9r77YEnQ7Fg0swM9RUtfnnIG2xQRKmLPR6a82n8BHbRLlX2
cLON5XRj09yJNs0Z2JCQ1W59NLivkiMVUH9NQN9L+iouJwWGCjcrZ/mbD/PyFjLtQhhrxv5Iejv3
obGw+H7u2jr5HnVq2fFyrZnWxBsRgTi/JQyg8sCuwZMgSY2OEWrTkMCPtB7aMed/OKNR5dOFyERJ
t+tw/3PzrQaRl04vFZlCDoGtBrFIq8OwsjMzNi3bhryPxtQxZVZAt0vkKp8gFUqMD02qJwlCsibb
V6fJQ9pHAPMH19ClJ6fQtASNnNmdS1rGr9HTVNuH5VRQ8d0+bDLXgd1gvRPORb689hjtSk3XYyh7
qsdzRbt4KImXScBT0E3AwgfRYPDk1I8/+VNHEXZT1EDSIxBGtIadEm6Q9ttjozIGl/J2ki9XzZXZ
tPYVj0jPyjcG8flmfHTgJqn5CamRnNKmo4IBtuDQqp2YoBItivJTvR6hF48TetKZ7/pA4GGY3/gg
V6YeBYrgMTA3EDRb4jo2cTqZmSKUGPx182ZNigxtMBh8zdebW189oPMIaFkD4iuRNWYw0yD1mDMo
XSdv1Z7GS0AhyOmS0RVNBoinW1pH+Ymcin4q8QrrSsedeqfMERKFexAxIGndIOoN6OKVfePUWlqA
auX4Hxw8Qkw6kZyKrTz8iERZS2v+y6mI4OQtt2MLWpqIM6/nYfyFRK3Pvr9gk/+gsLV+CpSXGU2h
XpJGx4S6LWkK6VBs/HcwDN/26X1wFAit/sV4VSPADvYM0yH7zB8OjNPZr10IK7bZxuCCRp9PPRiP
CM0vI4aNMZTFOZwQaDw85Kw/1br9+MbasAJ1j133PuEra9CYSnsI6ENoFCF0nPqktfsL9w9cgYzd
ubQmcs+JoRfCM18O9ZhG84uCjSm7KRTGjV8VvW0ClEY2FlbdmEUWZzV6IWJ4kqbU7gafXVwesCE6
LiVBLyMJmfQpYolhbaQM3YYoWw0PCpcXV6zCXCC8JxRB21CmtKR3rWyFfriX9TnEBPfWdKTgXHF3
hZGY8odTx0+rvxUHFIzprOCEPjUA0kXjx3ucYcgBshP0mAzA7Bsmd5pR1IgOM/EqAZSc+QpbAadk
aJ7zie4Ogm5Q9cuvv7vhNSvOgTrcxIMvP8asWlw2g7gnCqGDsk/rPYj+ZLghmO57csC4cP+jzD+I
+Dv3UDd5bPxl5YHGnf/1vHDklJ+qPy7cuXHLLQ9wKmDKx6bAAY8NX8aDNLfR6h9ota7/GPY0yc9Q
c0vMaQXU5EhHgvL+7wpJJZs/qt8SQ7bhnyknW8ZLtsv8PM4I2NhfBbhNegPELb4nYfoNgr3Vw8Ow
dxgZFdBzyqN3JFVPZcnZb8M626dYKFYHmvshWssrihR6GkGquJkgqb42yWdYMbZbYR7/C+G3TtKZ
O3yoZ2xnbJ9w+4g8xRZJ1oT+sXWzMxkTXY2j/ZY9AQ0u1AzS6YIbpKK3W2UNhPdW7tot1m43WBrD
pOVlqIwOZI34Su0i3Xdz8Iw3LL885y4tkFQIBihP0Z/GuLbwGpBpjj8pCIddt1EgRIIxns+p9jON
aAiAdwluXj1om6uPs/h/2Tf5uVGNoePsR1TiW7wKJQWSpb82WEzF/l3JaTk5h2Z3vR2VFK2Ljcsb
zoInbhD7+VyI9KsDc4goqMC4XU0nkoqdVfj5ApKZ+yUDtw6Qe3Z/TOtlbR2WkOvhETYNqrRZqFDn
CkqJoRg0wpXghWMGHvbyvmOEwuyXEE2lH5lSDu/4bFCHztyZu1Cav9aJYBj+1jZTWWodeqjW8I0Z
/3XDEwdz43073qJGw6SjmPRmDVVzZBN/uHaojXrDCd5fE10j7A/ss8ejlB006Lu1y+IP81CcjEJw
WUDLYjgdr1NTnNDy2IG89qTRh7Cx+ZTXy3TKmNocHOyTZNiWW0EW9gtwo6/hUcp+74U3ksbfrCKK
QvuTID5Ux6wb4czJTzOTLNj/sKnUgXUEfRHRF29wR7glkZ9efE5vcf8JCNmalhdAVq1LB9PTx8ts
u4CpbKC0g2cHqWNqAQDW8eqszdqujpyTVmEOzSuDBIVCx7OV0A+xmZ27tMH+ci7/1HuafmvckBwQ
83dfDqDda37RZ5tHk5hAvd1oEuyHjQnWJZ4ta/XCgC8DV7gJ+KG5PNdnFv0HX8Qp6exvh7VwHPPI
lR1o5g2m4NoZZzEd3IGTQA459AcA3gsLV8hUIfflYOrV8W1bjr+XPKRd1NGoD4FVcRoXATyxf1dm
m/m1ho4HXB2Hndf1iOrqyq2ifAr1LEVeZSsO96/qKiCt8YJT0Ovu/8IoK2Qmlc0ApyglbN4h8eb9
CsGux7VqShaZvVQg/XHcA2l9hhyV8z/I3kTuZKztRPwB/8zV8qA5iQHL6z4suJbvOsdegqsYmQnD
i4T5hHi5nMMsTHfllUH8XSrd08RmGRzhNuXk5U+8CHhXIop6jy9UwiauAWRjsxM4paPc25cwrsWx
CYwOz5c2eWhTMRoXnNJnkwDd7MFdeje5PZty0GyhskpFIVcj2Wyo6Xy3zjSyjPCAWx7MT2Hor3Hk
2kxj4DnFg3Kapdq+Ahah7kiL5aW0CKBJiJFdGMMHlwO+ShR/iE+djK8kYrASbh/HQprtuq/dEJ5F
yX6ZB/p6+w/ah1A9R4/iGWetRHkaLwSFny5ZypeqnqW5SBpkRrrP3vG8shBW00s0I0D+K31V4ntj
kW/jrOt4RTDyIkktpd18YAea6+Axf/1AbLolaP8qq81aNJlwjvaMCLOdu/0/rumAuNvHCubi/nNn
VxSGvH2QwxqW15TVwXJxNraQUZ6VlSKf4J94I56Iq0sOpAAaHAktFEDs50idn8I0vUOb+zskkoTZ
o3/mci+kAjKigIEuKJdxAtT7RCPBOqNGLklrcRG4V+yia4DyA/TCrVX+t+fBeOu0k+aRCh591HoW
3hxur4ilGOjGs+Z9argJRCzYWzgkfXGgNHlKkqbz6qh9MiNftjJa+Pktc9HAhPq7/Qwk7gYvUX/F
NBJLSYAp7Cyl42uaRDyfJjcZNDWWXZ9gCivELAw3z4dZoVDbsNH5b9QOe50l4I3g8PIK5o/ZlpcR
BYTwZU9ZwRVfYjnjD4oGfmE6DFicOg68i1QuA66Uoh+DqXZshEAtH53cG1sF6Yb4WuV9kTQY9ciE
PdPczWmne0dQVJpDjG7n3jHncMQINa6Lavg+pCdQp29flJIo1nnhv3IrCpZoH2kAdhW0NBq1AzGt
9yieOXkGDLQbpR2KPoPXYNHAsHvTU8/T7/PVnaSCwiBZDHMHiem66HioxSIGiDNtEEbeCGmV4xHU
RLAJqhhRO94wIjJrrGe5Ubej1dlg45HW041D/CBVlPQMbBIQhoF4JDt/iyHBGeB9msZNa9qx/S+J
n2JXhwaMDeHHIX3f/LjoPhO5+WS1ya6HslOxaN0larzw61ed5V11fxNnefdh6mCfsojtigVJttkE
AzsxZ96PY9A7v4uWaxEpVYezYvWo0Ht/AbsaRdHJ8TEg4AsGL8IrcLWcLLiWOJezsh2hCk0GjEGt
qx1013HOk/L9orlAk8MuBZOOoDYZxw+PRDttg3OaNtMRvgBLUKTAijL9dBasIeqJ28Bd0S+GzMfZ
8yWJcx75zWbYAuw3QMwNJT0LPjITJMLSxl+Y9aoDjGsgrqrJ+ZOICk0yEKT0dk7wU5heUlrOrdkB
YzHNv3YaMZKnBgcmkKwTCSMS+wo9mkQU3QOEHW2dz54f4wo9tUSy5tUYVjcIQp6reNmnOwDblGTI
+TAXmb4HIyKIKZ9KAWQpGuTDPIwHvu5yWelhn+yVdz6D732w5o5g+8CNhpborTUdLYBxzWou17Kj
+tJEGQ/+N/+aNqxM0E+1sMImF0hocXDgrWr6z417DiwqKpYaPHkpoEsAu9d5Z9dI5R9E2CKIlVDE
+ozBedU8dhM+BiwcvkDfwUMzjD0bZmZnebu/8SeFlKKG0hGqPb4S7iqEkp3Uj5+HNEq4+QF/lTBX
yKNyNAXpCCkBGZVP9vDdgG0pY5m7fqnZZZB1xs03rK8Vzb80A5u1UCG0d6ETRLj3c81YdQq4xrVt
itHii5RcpFmvzZyiGsyLh6Dig35wCA01uyekBOc3hewEgDN6PvXU/EYaAWFgwWZA25f+U6TjcW5o
ctBpjvJibZyhfkZuFGGNXYIvO2dmA+TZn+VF8Ga7SAY0EMfshReSGaZ8zrm68fD0GATiOoJPYyHN
69EjQ/GPwfLuszTbnC86ORWbjXdy5hGD+iiz6bj+rPwTI/kinCVstZozNMuyImQmrt4LihAmH++u
Q78zdad2hfRpk+T/M2RWlHqIFwuaeNnmDGseLdYJOUT3GH0BoYlwj/U+J1PqqbbAddZ6vkvYOfgs
h83G8lWEKS9/wjY9ncU4m/aRuLEgxwlpYNh6sDLWuYiT9ZyD0fLVLV3OPDpbbVXyy5VFh+SBZ2bk
mOIiE60OF9zaB8mjJVaz9M6JjKz0Uoj961IDVy6GU7xJb1ktFYDn3E04FYHkHTcn6KQa44CAcYrr
E8izYRiXq2gHnFkUvp419jY53Zna8Wq2Ab3DqKbKYCrsI3KXTVcTY3CaqTYgiuO+XwIN31v+0EPT
/9QnRyqcbE699TV6iibhRTQbl0M/0rTc3K0+eyaUCRTXeUVYZzwit88QkBXmiT24Xn7/46Fe3QEs
KbmaSm+tpmBEBaI7wBrUoRrKUruEEGwNUbXerA68DHpuFmEqIRK4sPQYh6UtHLpE5zfN9YlpSdTX
NhiG5+XwfNwM94qCoxqQXIW6vMtAhfZMvP7Ybnk8bg9JHPcvYG7ZCnWxEi8OFPFp5Gu3M1X8ZPq3
jFr2spQLRdlXqTVKpCSWwEUyki/k7O4orpxN1Pt0KyOWwYYG8L/j9eBjBl0P0/hCP47ck3vMOCcq
srCX767J4smHb8lzqh3Bo81ahw2pobf/e93Mxqhy1TMB3duOpHWRypQwrBAuYL7XJ2jpghfjSKnj
DvHVhk0cl/hdUPJR3O6wJJ6KOM0BaJIBiD4cNhswbUnVX+LdlOL6kN8IzvqdMd01F9Vb4HzC44m1
OCSss2sZlkrwXCYhKWO8AKSUYXWTsdT2k7h71MorBBm7vBykrOITEjrs9GgyZIG05xKbUmWAqUKP
kqQ2AlxCwnVp/lWp6/2E8yicjxp3+OL+YTFoOF0fvZTGR4JgmbJ9Np1pqjHSqAtLaX7If21NoPqA
dyqoC+UbYh9KK80sOcmHoyAn5+DZF7UcjYgBrj9nGoUnWqJZfwpKv0Nxh11QtwwGuyv8LLBqL7/z
G5iTGW43BIUi26rDD0D5EHjISBsYpXuaSPN64L+4ItA9BLyJP8r1XZPPb/MklgsH1Yw6aGrKuRXl
yVRyk8qMcA3z1ac2EC6m3dFM44bPH5+Awq3tJe0F5FXyVBqSSds5CyAo+YRowS5Xr6M3a0DIdmDT
/FMarPrEQjCZ7TZ/5ZJLKTWvlQiRbB9jjv6X97h3WsAhbL0YjnM/eaPyjr9QqXfCZUmbfezJSgWu
KOWcZ8xpwhTcCEPOnQ6QLmN7yqyJkaVY4haWwArfvSNS+JAFUTJdskoOdoBHCvAFYBHET8b6PNzk
TpAa/qrXOF4+iU1sZ4Kb0njpZ14GkvyHoQQ2bnRtsqdxvtPyDsvXRsaFT1R4ZPb8Aqtb3EBEIZRD
ZvLqas5s5k2sbqCgQ0/zU4WajomOzzTeYbMETrvaSq+pF2bi+PLEwPwJk5Dc/G2Yt8xCwffeYYPw
AOvFcH4PaxcWfYsiCyJVxRH6iuJrRwOjOCMZb1XxxbEECm08jiigXS5+RHaqHyIVturjeFHLbjvN
2C7CuK0zC2adelN3VtA9vhK0VlJ0UJCiww/V5x50LsaHdMMtEHLaduLMdL9aXA83S/TXVhMDgUwn
BnZetYWZU+00vJde2+NeMtAyM35QYa/Bs3cnDgMlHNPq62f2Ntls9OMBhTIIq2v5S2OHwsz3CQiq
y88FtkL6ndx5hdEAvTgb06+olLlQWO7nT0/5nVE8Tr1F1SH5m8mRXpfB5ed+crhB68o7Pi9f4Lpp
WTYiV2oOvplxAYYO2OH+bvoBFuisGX5GjCpQEqnqTu3pFhN/E5CgulnSwLAZsPSummU0bq1L1Ifb
fwTldBb0C3ZIsbcETjCEATk57/8i6Sujhst2A7IEX9CCnHR8MeqfhOCKHWJd8RdammQF6b138FA+
OqBdMlb511tKKHupYKfySOrv6pawNxXgy4L1cgriO+h+HHOi/nT1X9kuDYxzk8T5om1GZQB5WizT
0NJgP0UvJU8L23tF8h6ZDkSRElI0D4lmFbF3YEUbQRuen1MKze64SK7Ba+9HpnmFsXBtn5WCuj0F
Jbz/5YD117Uq3730BV6e2YY81aBhXmLf9G6+Uo0ebMN8HKdgRoJpNC2jouvATV76V2pKJuDcyC3M
PzH2R2hE9r1ek89/7OqrlyXVNf4V+XW99DsetxaLQ5j1fyGN07HGxbY890EQIGPcP6+w//njWR++
fipfOJd/gY/bbQ31mmbxkXI3xn7PfXlUZJxDStLEYzjueTcG/L7ol9Qkr9Iz7OKbW7Y7ymBRCzKx
Q8jftMDG8pMuLcpesLuZV/0gH+e3tSnRavBl22d1JN6XSsAQN9kc7DtVqA+bVwHjYyiMZlUf6fCJ
axNJYvjbDNN+4VW9bipWo7Ghdn7eEFJBpVmlrhmXlfOErdNkEYfw6h4bjTartVQ7HOmQ6WPtjvcp
pVuiYk6+p2FwPSaKtZan+kLPOXXB04Fgz/FtZ1IzcIWppkyYKnB7+D98gNie2NppGgP019n0eogF
C24wmsQer9EAI2OSpjnr3Uc/PA8FlphEqb11jXg+aElZgjBt8zKKizOmK2sPgQsKVhN88qwiR+60
Coqpmnjcrysa0G8BG8Ex9DztKtU6S0buHu01Hvq6YG30WJCUOPBZSiZgfnPUB/OHgxcFueb/fpUb
1lgvBnQQOqK43Im5HZVhJWR9JJDXtTHVy3pv6yxEnoWcN6qVqx0MZ/K6NlJ0OoRO6bT5UkSl+lP6
wA/7m0GR3T+5FPMtwJHqeXFKCLnpXPWKH7cLLNFeFZYGKFYn6vclh4vCYd7hoIHwIr4jmEnFhldD
HpWx5KgFEfovwf2Z/NQB02iGb1Iy4LMq1WelrG0hAH9F3KpK8wsuVNUW6J+qQuye5wc7FjhKs7LD
soIaT7iX68kyMzfcLDWFAY2QnCUMl/h8ETcxzT5Tm5gRjVfBiNj3t8xlprqzNIfyUu39GbiMRM4G
JX5kW+2a1l7NXO/uFiLuaaL7rYqRCA6er0RPE9t3gqln0BL8sifjRpIoZXzYcoRjDs9j3R8Zdhz9
gJtSeemeQ44CjD9UczhsGo31qBYiSjNwmFr7OtwfoqU7sXUpSrhE9103OKoIfvjH+MWUsQFjP2An
9orTQSyE3fGqGMKk/fWdPYxDrL7aMNNusinMHX7P9BFLKXoV3GyuRwgFEelj8OAo2RmS7J0N6V2y
SdBvxUD8WpFzm5beQ/sAdq3tp1lUYngPv4H0Y+BoeMz6BN5iSDPRM9CaqtxTXT6oWyHMhpINqZGu
6tPZP+D5tuzc/GF26gO3zYSmwwLVY7gafwQPe7VRf1Tp0KsiLC+JeYr1HglwRsZyUx4wF5mmQR2h
z2l83KbbgvtXUCANymP8CDE7JL9AHPtsMXdibGnLci9gl95c8m4ej7Z776EYfAM/OocVXqdkoKD4
Why7dMCB9xlFOf0jdBAjUSCrsVteIwbOHZ8CsfMpIMWmPw0XRuOnhIyqIFg0BlTxlYcVZlX3QeuV
k5Cyckju/6+bcMOOMqa5dVCBSFRG0MS1g2MmmWaGMMcRaI5dR4FjxY0IKGzCrxmJ89dUwryhZsBX
B0vevQuQWPLWXm9hdrMET7pcXDyJK/A2U9CjOnGIksNYDRmOfQENwC663LZYQ9Zsl2mWwQXa4peP
BN116X/xUm8FS62QdjTdx7Q9+iRh4KPiNQCbcUJ+OSTwJxEHol6D3347gL5UUkckvxGkBpbZwwe2
6WkIglghz7EoxPd4xvnaEaPKq8XWcpLWCngmouHQy7suF8iaGEgS2z7M7Glig5Iy+hzKfrmW12ij
zuoBXiWDb/NyWXqNV1tPOpeh/QtQEOdzkNH/JdO2lFf9CMj5b3jpGBACYcb4YB0vwoma8OjcUa8G
14xV4WyQaoihwv2ZEMwbLz6PJvxcQZS8hSAeFom2uWVmwoXbudJhZVxRqWYdf1WkNDph+aCvBWq4
3KJY9NUeY6ExpOosNxHVKrBLrLd0M3Ql54felCej9nGeaCoe2Iw5C+nTcxG9GGxrNO4wlOmOKCi4
TfdpCg/IYSfApJifCJEXmQrsCbu0dSj+3reV954JipkpdRdRqnf8zwkyffWdKuQY6RPaNpO59e8l
ccRDds/kFOZePk3R2YCj0jkfrluXLfZVAIjM6q5P65oVUl73pftyU5kJ5xncBo6wEEEbnpfy5yeW
rg3WcSOCvNLqrsdArjewSb1IJnBw2kfS21w0s8SXRnK+/PZmEoiXdE4D/EjVMdEJjdLtlPMqpjlM
SjsFS34hqFJZPB6/1EqPCXg3PfG1goqV6Ohq2jr/IiAfHgID0qLlA3Ikd7kOuGU9vRJTQEz96ifO
YSpy3hvXKedsIDp0loVIgrAVF+dKonpRfAcfdwqS5/KuHYO9nbzm/0W3IKWlfKGJtIPEtDwZuMyo
hC8hXw9C/glRFl268TidR0Zzu6QEvTidDvzR2LvDTxtdfGuLLdxEeMxWwWQWA0Rz7TI+H5CRV28B
64UMCTUCX/VR7nxhzzRPn0Pgqr56tANiTYNZsEwQtbhEucBjbyAwo4RQxK5Ao77sQi9/bzJDTnnZ
oHFaE7pE0OPhSz8H+k648mVnZEzqDJugakgmlCrGm+drB5CtflpAuLY0HuuZolidAxW1+XdJFZdW
lD9libbdhBmP4lXtq6+fFvt7a/K0JGR9+dbTBlSvAGXqF+Kj0q5x6HAIkH+VBNPF2uZ+qv+RMUPf
pn1C0+7kBLAW60QMODB8Wv/fzkPyKrFaWIklzkiZTLjIQlN2D6ugLfKkNjbmVLKWVfl7Vv/HMt9o
c1MtXs+0VJ7xWzUI0DRHA7Dj+O06GNAEks/wK1SVR7mnTp3hS70iz/hwpm8VLWn2vBSxtfSYrXKG
+CnKBjuaUquolAU/ZauHbLQa2mZkLtrbRbkp5oHlxivbBZzvXmzf6VmeLuUHIq2SiUNXEclCpeRt
4Ka3vDWRhKErxjDwNn6HyCpkNWQgLLeOhrRlwp5PCv9r/+um6e2x6+Jq+2xhjYo7jW/WuhEwT2sn
/9Yre4kKUnIUI9M8PYx/Ue9ku4kJnaM75KmE6fykT5HlQJASTxUphDgXuCDbpgO+v58ReVf3Cebq
Yx4HCeg03Fy5RPiuC4gD9YQOHMsQ48g10TzL4y0WW5F/JTYfBySnwNHo96PMXFd2RxhOZtgF28dy
68qfGb7U3V57Ya9Sa2Pokj8tRncety0X83w5G0NKy+0ZGSZ+JMZ8KA9n5raK3JXSraUkgHZsJ2+s
lnqe790BLtqB80YqRdt4kRUb3XRuJ4OGnSk2teoN2Oy21bP6GerYfff8wGpF0ZbfBZSbU3tUP6Ma
TUgZCawZPuJtsremYSEQ8Nn36VfsiRJTT9IChjlRi8X4gcWxHoHcyi/hjw0ityZfQWvnnuRRD4dw
y5FWJG+jQnuty7uENK1D0gt9EPeR+/SbnmhCl5fylULe+LB4kCE88LU2D7TNbfjnAhwBEPPridVt
6fhXqzh+6aZKh+B+Vp5oBUrPbFNZdEfYTQCzFl5dwziWTLbH5Ty2yX+stmWDni9Bbwb0AtlKxnUG
SjfWEAJNuOaI+v110lXLYfukJJoqruuLGjpQPZULGIBWPeBRETrRPTIs1pq5789n3pTMq73Fb7sr
AL3K2wkJP5ZmSsysQJk55sN30GD4nS5ArsYOD3EghqrSFKvB47A1G38Kz1icHKBT1ppBhR5okw0R
3l2LGSPhTNSC6QZyo4d7zA7KZqjB5Fs7w/7SEhSQUc33Mz6n4T2jWwYrb+qYX+xlV+nkwzl14P/8
t+0ExdJ47by6XfHEpn5P9hVK9NUZMOveMM2iClKTbj5Aw/vVh2ssGQL5CE1VOpzHwuWMgzzQqLOL
PJDzj/arPbzrdUg5e+FOGV1Di6k12AfkX3iaF2HAKx0WapJ2UOHk+yacmiKDPTYuv5Bz5dkxrIAb
1gebHkgBfFWGy0AAefB3Mll86oaaWuKIm42hg+gHv3lVcsKpFWoRIZuQFbS2lSCE5Wb8zizFntsi
jZ6k0grOUsxN2B8VrOPCA4ULV6RAYpRJFU7AlUIFI8rFVWilgIYw4kbU4pKdnZ6o3AlvTrLjlwS6
7jAA0/HQsUGqtER2MzeURkWK3RzkNpraLVz/sP9kN6dy1aGM84wZ21AvEh3TOi1wOoudSp3tg1Lx
R+yDh9A0lBz4PxT6UDM+hzRnmvBEKICfXebCbmU+Wxh8q3mxFaXG8UWVEPGzxwC8K6GZpNaIDgJy
z5vt0qV9TpvDfQsnCX79FTowxEItAlzf/Eib3TKpNCdEknL4B73hSOtWIaemuWVy/aLRwts4NoYc
BBYdxebp+WVWQq27OoPhwJSqzyg4WwUN06tGdb42eyW3bJCw/N4h7kwKNlnTaIyCTE+3wpBfAZB6
7hZp49VlPREHBE+odKlNTcaqEECbzcMvWA2Y0IK6cBTCzaTGHPkQ2JCO4S4i4D6sKOUuTc9l95BQ
fcFK2zvhxzaf63no6cjTqhmBPevlb37zBnEjJYHBELw3QWss3Py7Pt5KLcRWLpw4sv8VvP/TKIhW
ovVU86ieoADnl9zoPY8BlUL3Seh4JEOHemvXiuVKKXvUqZXk+yAu0PZicXuH0SDhtd1WlhTeYPIR
c2vQChvkGLEYltdjojK2pUjIvsoZ0rn29hjt8gB4y2f82a4aJhGKybaKPS87jbi3kJTqbPhn9njZ
iGP8PCkllsR+Tt1GD6hkfinB8+qvmyzpGpyk5qK9EadJS0Gf9QUb016eS44cnHQjeO6UrL9mTNXu
vXRm95e+BTzkhrx37N/pQ8Y9FKQjAunAoayVOH8jUBVBgVGnG0aDWwHywo9G2xPPaSscSkzhAO+a
vpYOKz+5rqTSDpvpylTkjVaHzuCBX9zKvHMAnNFJfYpctaLP/N7cKZSnEyBPlZ01uXg2voc5oBTi
/obh/VpTd69u4l9FTA6WWgz9UW6AfQ/2uXsFRsXa1Q6vswap0KNt/j6nwaJ8yPpRZ2LCeVdgQ6he
jC1nfXPLB+eMLCEnvEXFVylDYgi2V0FrQ5/sPzjMKoPV7BB2P8RoiVmVRugCLcDNCugl2Oeo2ybn
34JDX67mgBmaGnqVuWyV9f6kfSuPnmYEM/Dv0Zkrtd0kCqpW5VXOwmznvYMdrGC0DEJvS4a5k7yV
U6UOmbOECerAfPtaQIx/oNz+mzIDP/p7i3KYgNg9eKt/Jc2m6Mn7ZEvdEDWtldV1U2m+iNj5PIxX
cE9yxwpHkgGC1W2KOaX2EWlMrUjfFRjsQgsbxTlKxXlkg97vnC5q4I7P4z6rmMJHIFbnDt4ToQJ9
ClE6SiCzrbobytwISf6J+9FRmq83TadaD8sUjViwXc7JbQR1sutZNMfwjz0/Hqaj01Vh3z5m7ZVH
fHL/UDThocuNo/qYiTuH7mMX8iAUBHyQ9spYEV3z/0H5FKoIEKPCT7U3eWXhHw2hf5lz+RHZ8+kj
s+1w/ixb42RNuZJo4ys8LmE4aqCdp4wf5ipsEpq0s0iPNl0INw4cQsuePKVZ0XglNtHaopzlbsJl
7pDM2mX2daqp2/iI0WYMj7yIc2Q8Mirzlol/v/HCnm74eA11N97PQNJoQhOXEtxLCuTowkJMOcOr
ptmrQePpPTAuKhDJSfRv5Lt5OJGS4q62etC8urQ3xEgWxeaMXeJz28uzvkEhAsTJbWBDvjjWvIVZ
j6G0bhTP6v/syVm+mMiJzNNN5W2DBSRllHDKeveqDK9CRd50fbV+ab+eeHca4RhEMqHA+ytwrASp
w/VbwdNW4rl9DjC8VLTLJogq+KR5opsG2VqTSypvDjR0oUbAi5v76fOUEj/ybuwxrPpeyVLQZ9N2
c86vAey9GDICHVnpeD7LUwevZ339Wv5kj1wmZfcqPVXFmYyEHlyYn86Jdjzg+nkp69PsD8oiTsdG
jtW44ckIgV27D419TIMfcJtg6pn7yug8mH+Ch/wO1X/GXlH5/7mfpb3w1Ch+Xx04gb0qeKfh/sLR
7HgD4i85IzfYnMphtoEQPmVWrMnrEcLaxxZOqibEQ0jKhrmpKC5ez2JTG2z7uJLQvfLf0ROTijVU
kspG8I/QgYuYNI8e4vxPcxBTaK5HCPtI0uk3WkrUGChisiwvflDfun/mGeKBbrARj90eYgvT30aZ
JxJHVrCH0yTVu4Nkwjsliv0XozAxDuKbijyuxl45A+9mezHp4O5Fxz7rmstgJfe2968uOlJprEn7
sBu0V04TnzRGrBPfaNCOJLwbva4uHRZzjetvUPhKcbkjQS/40MruITL6uBt80qz+9Ord7Um/sqAn
UVg7JxvBDhEBTbBnbO9Xtd8sstI/lF6H/4fx83z4STAifF6ga5zDxzEIzwoAon63n9zkFU8nHZ+9
/6LNoxVQTc1aJdeaUJ9Hqg8w8cEasZEMsXm3ZEAus3U7PPjFeRs8nDH3uvDIcYyed+CQi5dVA0vb
DijQsOYmRlq+jd/4KNmcc/XflZVrYEOJ0oqa5ameQMIrEdj1Sh3Intt05RlLHljrjV7MuqpAZzQF
9VsscknC5l5pBocvYTTiHnzuSk9CgAa1ZNHdUDlEckI+rbXpXD/EoHWgZo0VDFJWvB1hqYks+tys
7D2ZaBo5uRsi7bBkjDtZ94sLS6HSTEHHCayCiKY94VqheACIdENEawfoUKsGvI6gv+oU5arG877k
BftOcqeKT0NPu30qp50BAc2iQSD8lmlLIbiKQMW42aJx06Bze5wiSZEigRtbr+iSB4/7iQuCABeP
Yss33dGJZ6KJbY4YizmFfGLFjWRJeOzfKS3+5DQL25sJMuQXGEGs5m3B7+kUhFa21DGLUpiGM4ox
fX1D0q1jfOGm/e6VEIMBzqbcKVn9N2NO2wgCMgFCwn0smhn2YnwgSx2uHirEFG0S0KhVGwqfDnQG
KemeSuaC18IcgtzZ5OAN0FWoj573x5wWPeYFLviNu6EBfMcsHiPztvT7xaisw1acBIfwciIR4Ztv
H3xDKW2Zhoq/vysUe/rhl7PdQebcGitABLVY8S7Lja70FxsEvHCCSwNZlxPVaEPR2vtYLyFNTMZx
e/xy+QM5LORZQR6SoEe1pGpRdHKAP4fYwquq4amKJ3pTZ2Nibf0DeevWXQr867F2U06muSCD5B0l
wOMo3hgN621ykFFU3oRa8/rnsdwFU56uN3RfDQ1iCqyNPOi3L0PJt20M0ruzTPUJ2cqAePwx+Zri
o/O9vTi0yrY7Eq51hmtX54KxKsa8l5iRW1YH+xGUFiHVU2m7ZGgGdCPt79vZSbk/+K39BHoge2kp
FOj2Li3sUVYYMQPM6XJw1jI20LOEYKeQV7Ff8Rds3m+X9hHBtSozCTx2T0KApSNK1Mt9snSmaoh+
lLXcsy8EMoA0c63yU62KR1k9j64eJLLK6rZKX7ZF+oPXeTH+tl07YCJUmpD5hAmkWxanjkdNL7YR
ZXwuL3UO2EVm12RCx7kzmMz8PrkoLwCHe0Ll0CHmmC3oYZ8WK0FoX4HsKiRVyJ2s8+sKpupqApif
/z/mU3eDqdc2FWmI4XuD8s6zInmimV6YPAMA1jtuIfPnaiTP4rxCjLvP7cNESs9y915723UmWA1z
7ig3uEQdtborSknpZwRLZRdrXplEAn59wZRRadcOLcy6m5hpt2gIsi1R5NL01iQuUCkLlopGX0DV
iXLjywWixG8HuJGx7RS5ZQSRPQpz/UhjPflfS+hn8xcxngR5FhXDwp1M1qvTIcbzmKRISj2OpFgg
VBjdsDrlHIfpctfBe0iJR4hu3Keo1uhVtGdasCk2gTONOZolZeePhSf6KRf1RskWCLgiUYeJi6eM
gPGB1PfOAOWBmVCaK9rp3RFrFa7zJjOOC9YMDzT1+D/OyOB4VfIIBicAABuODBuexNsm9Fc0F2GT
w0Qqel0Yy5wwac70CTqUPmuEPfIj0CUkey/zfnX1J3zs7g7ZKE9jdsdsdh2G1+AyvYuAt8X8YHPD
M6r2yrzcchKJIPa/vQKuwNPUDc6gMwARDr1nfpLNW/YK0w1bGW3zbsBOuEbvZr5ezCfMwCO1kUQF
fSlm4z39V+Gp47h/EdnGifDNJl8fv/p/8kKNc3dTBqJpR0sTPRLN4xEQ5zi/Cmg3tXIWiiECjQlt
5d0NwYf3mNp+/Vf2uAmP8M4OlVCA77ecqR66z8x/jQO23naFpuEtTAabJ4Bmz/ubmZGbIvB9b2yS
Vo3ucV8oBvxL1air51BLbzOh8dns9fr0COtc3Bd28eGiOVTtVSlYcBKK786Ey7J36EpVoTAFzr0H
2e/Rg8rk69ZcmxhqHxB+W1gAQtjxvOTDl8zn2vemTR6a1+KpoRIyYZS5z1ahYPBrOrSbFgCQ5vyG
DX4+wVhv/7fHyviJcq/UDpkkr7yBc0163Qoyhn4Q0wXUlMHs3Ua0QFJaBReF7xnfHJyd3xtWrZE9
cGLJ7aOGy7WZsXgb3SNx9bWOXjyidrtdgUJ8f/V0iXMq++LbwAlf7UkNOeExv3sEC03633iTLvod
9sAjXpP68nMz+WBMkbzlWVaXePwb6c+kfAUIgWnyXswNni/idRo0bYj2v65C4xF3dTdT7xHjVs63
WM+54lQMpQoLJlR8XiTGj1nwEwENiTvhY3LFQSb8Qp5q6fCrkLQoEseozOElxTMuiH9KvzbkwTxr
UqlG6rbSwsZW69xQVDvRhM8VCbk+PTtR8WqhVtojxmw9YSMLIKfLSym8GODXCtZkH9TnpL62Ushe
hbuiqOe7klbsY9Z2SA2soeGskJJOuYa9NIWgvq2z+4kFq5slODqGv/ATpIypgga3H2kjOevFzKrS
e6t0m+aQw7EjsxBRNNsIFjshOfFn3LoAH+XjMQDHiIqmxN8ijzKCHfQmML/M1fFNSpeRl1BtTxHT
Bx6oGW8mUy4HV9SnhrrcQw6nZ8FAPCRYYm2nBouCT9oMXWCMGZN5sYk/MLqsmBlNN6oS7MUdV5hw
hCzBqfGRHeBqUmeRJ/5nxQPEsog9Wm9/8zwa4f0/9N/9AiD5Z6E4ZSj/fLv8mxVGQtt9mz4t+jAw
QiiFiLbpz2B/FjxYMuIMxxkZNg3eNri//U6KAp5upnXjfRAl8f3kH9nT/K7KBeRbO8TRq04G1/iw
NBHZOkRyZy1XgZi2jrzttbiwq1VneAEPP7aZ3C/CIXQktk1bil+Smttw1jf8I3VklqHf4XMgY7fz
otqCb12IZizD+bSSFFXtVPlJKmZfbJD01yB461z5j+uSbWiw/3vpHZycrVS7pHUTjr2bk5W//ZwX
r9ay0Ct2d5USFiV7cwzXNUNSsB0K3GMtOWFVEYrAlCU1yoStL+vnej/bJsGmKz6wwBtTgb2fmnGZ
mSIeZcp79ywFNWqRlWzo3gzIt2YNjBG7DxU/aYj4ht14NtRnu+AIhdcyB4uhd0/O0ydIk6ekwp0w
QSmQzKEp2ltHniO/CjbnCyR1wv/qnsruYDi13HE57J/TdPW1IiMY6BJhMUF1r5MXWTFRrCaku5jR
NKyQ8amgR1ex5K0Xtunv7LwhYQeMao/iBnWcJwD/x+KjE+FTwmUCLT4LkgeuhDg/rQnT6MbRohcO
o+J9kzwNYCP2+B+tCTppmN2eajIZKpMRjbH3UD8dYIKVoD2NlVUpwuh/iMZRSqJvBlZYG33QQdr2
g+FfcUk6PBcDTAbc66OoyYWJemnwXQL1YpmPFIvDhYUCzj6VX/8uXPt8UEsH01bGu7ckddnUpsIo
y9sWpxYN/xuF3ETpMRdpXpOlZPEjBsD0XDjjz8+4rdkiVTGlUdRS0TrSrBDyQ84YvN5rhyzh4s4w
emKaUtKQpdGQeJVkftmfK1E+ZzFsaw4IwY2Ram9p0tlKOa3S9CMlBnm6xIyNtSsS2JCws5p0wm1/
VbET4ByuIZwtqatcgrnnuJW0gaYKHGS9KfxKaWvQMW9LaMH1U0GxwDSHkY0/EXrnKv0aG1i13M/a
sOxM8RbQsjf1Co2GL50odd/tw9D1UzXtExNfZBrgg8XRT4MGx3cErAMJf0ugoVTSWbGYnQJ9LM5a
Fn0odQL4QHPh96RQAAhVNs6CXP9Og143b3F4sELFnFproITpOlNUwt8K4xk1TV4GjN1cIEzQEMv6
H/zOYonryxs6e8v2l6g2OyYjDfkLhqmSnKGCdaQXzPyeFFJIJcscr/FigGzKmMw7KyEg2QK7wBiZ
A+I9h+7FQRdTwmjJ3WM56nTA6xJwPUtQrnqdxTNl5RfLL7zwIZrHKPV0W21ftM96XKNnHUMau3VQ
YTcVtbPDf+oz8odsniybwoMDL1bi3kVR7RumSSGv//MHH9+0OhE36lq9mozbkT7bSmXCj6wEnxVC
XTR9gDozTau59NcWj881W6yP9RGM5wmrB9Ge4HI5P69UiADfrI3DcR+BPXHKKQvgH/75XTZUyR7M
oagzPTC2qXYWN/PVehOCef8PZItQCA+UmZCX8IZqg7AunFtOfuYawqqNNANfdZC/HT2FYlzwRv1i
MWtschC/HOTkc+t2v7lPbGjEgvG6Z5+cc4cZaZbu3CpS7E41SN+/utjg0HrTKrVXNEgDL4mvCmYo
nEhQTiACWMhkS63HoU9EhBWykGgGjkkRI0JVzh8pTSJtw2ENwipbw9NhaCkv7h0RK1LXRhkppLaD
LdpI8sCp/IzdNxhkCwJA5FKK4bCLPfNrh6e94B1306oEiR9ytHdSXlLB5RuJiUNcMwt8yKvj3cTs
CfcSWl50q2vZjA7reM50AlqP5dDTY9QtUmojg15eX2dRlT3LMzZeMxKfpfmZ1jo2kJ9OFuXUG/kO
93Rk3oksGZ9uQ1GSZscIKjvaY6VbiLBWEU+sqJvCFcy1z8LY0PvWfAy46T4EDNXHc9ASyGVhkvQG
9TOMQDbLq5YuiblDVzl43VfD3flfcZNg24b5BY8PYjjijhHuxWuD46qteRozBwnNvDf9yy60yBmU
bqX4RkVgmpv/RL2zVyNr8kMjfkLbnmrl6qw+8uMHOab1UQDMzPXcXhMKnz/Ndze2fKj8R4KT+O7Y
HuVa5fIZNUPiKvSaGyT6dn8eJPOim8NhVfAs1hc9+wtCA+C4qmFbOpE1BQeF6pvG+EPEgoSyyq4C
wyhAjfijrXUgZy5fue2qEDVNjSXCiW0ShoNMJx9HI+HqRTTlBC9RGPo0RCY0WAymosjQTC8z9khH
M1ay3Lz1Tn1azMp89tYz4cTljlXyZ7G5JJZvharI4srWxHTZrlOIYMAgYTjxthqDaxWGRZYgJQ/B
jBBmE6NcT0ROngzBUZc0FlEu1A9UbcR8eOGYqRTtbZ1ITcoC/MGH3QvPn+zV9HMQQgqYfXmKxlRM
QQsaD60NDEcAzG4l8AAaUS99X8QJKYUoC6kyzig0oLRG2dGYFyey3np0GOJ8QxsxIn2zorRBy20F
GFLKTCx6jJHhD8G4+MyxMv8x20Tr1vb5O2qbTc17E2XOUuj6WvsS9txc7H9soulmO4Rcpd8IyqPH
AvI2OCQj/MBdMkqRyE4DzyqcaQyAb+tK0F+PYMAfL0VFpQy4t20Dg3JIX+MErrckVF6RFCpBM7Sy
9Q6KJRlGkmdBemydckfTBwQp5CVeNu3DhTBiErehNX7v9QOZM7mxqcJhcUmCIdoTOO3uNmivFUuc
TgTA3AhHpS9iqerb1rCMqrTxCEzpkLNh2ULFEQjUoKBSidYURO2sPlBoOpNcKMocIKhN9+THw/O6
WGLS5eJ6W8OPE416+GYQcbrNBLT/7AQp4AJdnxvm9xVqofVaAf7eGTZydcCRMkLF1voUjxtdzcGV
AodksObfzrG/utOBXh8X3pS8IqylGD/KgtgZRC76WbjbdmS0UfZwHaHatGQQCr4Y+XTfuN0wBiAd
6PIuDon/oe8ESaNjCbBFzjCtFA0q69m5jC/yjuuuUbiXfZ+Zwyx//lKdkzTFkV/qRbHShWw8zc1u
O7kVJUUWr4FhwFwWT5l4qpxz1SByTqnRpLwZfKUYusYXzga6n5ycQOKUiyosmXhGj7Cj15C8lJjL
JVWr3o/R5gKw870lyY58KbodqJTQa1EyX9kmf2Dp6VyyOrvc5DIjwtgk5xPN5lhIsBYfhbSZDcWU
9YXRM3VA/f+LwU+suaktqVC4TcJ9E+fGUo2zEa8/jyXncgiDTiOytxOH3TpA3yvKaXrx4viZ8P1f
2jzeXqDWARZqmk8Q4O8fPoVcAztbtlSHFcohbQ/ADCVZyH4wr2n7DpX22+ORaMT2tBehRtAiIJf9
wmBwReb6DCfyi7D7N+cTW4N++KIvPQ+u4jCcEqroKGCfCzPH7HnVwN4W/edPARbCyOEdKINCHkPm
w2JL9CLx8oMz75+K76JyJw8Ey53RiXubjujxRnDtLCD24mC+GoSz93BNazlvUGqnGGk8Nj6txAeL
mmKKVaujwqmNDzq1zkwXsW+n8CNJ18czIDEVJDMVGaAl9WA9by6HjmQOD/VjGU4Y8kWWXk/Cdzw7
ULmaJ47jHgK4iwm57/ZNxhSCelbHp2JjwEDHfCgjfPnY3JWrQkqH05+vuLb+OO2a8H+fCjt4LPeM
Ptx/0fnbvc1aRDH2wUtWkdiF/8W3jq4VzOkoFbvIw6gXBTf3y0H76JMTnpG2+pVE8OhtthW/7oVL
sm/tiZ7Jnv0B89kwE5WLoWs2OLVxUcCMThBcCpZthxoQd9VDxo5+7tilUB+uVyPg5rmp7xji0nKx
EoEo9nIOcIWh4gWgN4FnDY/LHATk+7Ze/vHClQmjx211RZpoEzdyJjHuRt6tbv7E0fJC7Q5aebwe
KcTWoJy90spORAR96J9cqtnvkCv0DgaI10lS2jUyIO3ZAw2tI974rmGu9FT01FyTo7wXghKRPX1g
ictp8gKMarc+DtkOQAJ6illRo7NMxoEsQspWj8Va8l8aTpwR/phnTxRx/gSS9kawm1UqPa/VpnH9
JV4Q4OMxkJg4WyIgV1i21/WaXaODkJ1WAndyjzjwEt1QR85jCY/T9TXFzHGjdq6FOVy3pWE8sqXR
dCFn9LxaOXVjQPeV42xlYV1qGj+fLywOa584RQmCQBbN9qtl378KchtLrZndvzD3FjTY1sAVT1py
sEqVIt/apFn0HeAo7VeepvZlVAesbwxPZM06YTose3WNh2iZt7Lg1Sn2G8UTvqF74/3+dKlnKsba
iYDEFGIMCdNNIoTJVcqx7VEcFe6/fxljYQMJlkSR5ZpYaowPb6/9cjdTpnxMJk3xQWGx0BmEyZG4
NXl74GvuIrsxF/rr26Qic2He6WMhQ/AUwmjwEmr66kAimcqsgGBF733At4gJz+MV4fQUuBZ+Hwtx
RHgFfEVkKmLPxhjddK1p2ELxc5iYBznQfiItvliMPVLs3UoOM6SVYTWbXnkTaG5fhRw2LRliWQSh
W1HS6aNCe6cF1rGziUzODb3SyLguY87Rf2YDIecRReAYc308rIDobim4SCyiwQFLC2OT37C/O3hj
TzIynq5ugpgHGMZUHIWoOWhvTHhxV1EHb0Z/0/L1oOtbSSMeJBdTpxA6G6kyxxBsac2jibKj6SJR
FOOTPO7BCrraK+Qts9LvIfYRostY+CssS11hXNtS+xxUXkNY+Gzv3o/Dgku2ft3Yk94JGmINogfO
PsfVZi1DIMTUfjs3i4QlOrnA/Mka2yMa0nXmHK9Ko0wVw8r5kp1CxvKbWrv977oiG5QH/BwSKUXr
TiTGb1fjsevGuqtg/qgIUzkI7hhw6Se/lPvd7T+8s+kSWqqWB311muXlsiKva9tzCsSpuBVrfxv+
BKBmYLZc9ymwmX0XlnKiIC7BDf96mZC7WSQcIy/g/0vMTtDQvAwiKGg62phsEOyaHn7tHxxuKwWM
p7nEulEd10o3eXOaLOhSo7Zl/1S5Kk34qHHvBcIaype/ifoD+c1iuKWRrQq/ptRL5dAjqC3lmHex
V54u7CtvMl9lCU4aI8Kryk65AKPMvc4zhaqiNuCpHQ+mCjzzqcHcj0mKivIIU3KjMz+A/k0pN6hg
BWH7JNhJgfw52fx+Awqm/8xC8H7BXwhDok69rssKtRKqK+K+4N3A0iSy+gYKbESybdF0Xsz7WkpF
BWnpUWMTQMlTsMWyVIgPeQo1V9ieXgEKEZL4+LcMKdra8HIcM7ikbCSb7M9rCQGIkvxC1fEjbNWC
VqrpS4zf2dbJPidZ66neZu9aeKkaFwymtFTjFBSRS5JiE0Lyh7MEEtRPCIzqd7pVjTKowh+BTCAS
F8fgFDwB0XhzTqS2l8/IVyNTYzgLo579opeJQkvcfJsG8/x8cFUOMq1maLzD+4nHinVRO8zc6TTK
bN8u079YNJWeI1e/ow/F0XUviBMac0APMFbbw+PB0GQnR8tR7oz/1Z6Zf26S7cJX8RO3wrR5TrI4
3iDnn/kCNuGMtP0KNy23K5WZV2aiaql6dbhDhiL6D3fWyEaR4FUW4H+IrwieWF/rBh5XEyj2t7au
DADlg+r+JiwNi9Oio92EUcD+9n2Fd+YkjBdh23hBDbuTHynA8T4JtnhKWUm6y7OkugbLEXemUDgz
awisn4ZG84wgNCVGGElFWu4VLdy8cHYa0lb4VN8XNeklM9swB8gHpCF2WeUoGmE7T+4hZb49dKiG
RClJHoQv52KAcr6Uuu9k+Aj3kARq+IKzmHH88Bqv2ClDZVYcsUvDDuBkqXjTnsI+fw0NBLEh0RyX
/V3nqUCktviC2TdtSZAsm/6oLEb6k7cCrwhEFhYDwVCAcuTy3I8LJ1xErHY7M97lQbyyc+gr/Bpz
B9J+7dkJBff5rQdc0kpTUSFwNJ3nm1tGLknkX+9Qc+Sbnw4Jh3KFnUfWFWC7Nhn9CW4u5isWXEDB
dA0sEfXHsDgJHaClZu6+oUQ3RpPPObwIJ+Ch+O4xA/isGxFT9eDUlV6DoxL6AVFhdPuKyODq7r6y
K1Jx65h1ZnEz590PJ+SA0yUo6TcslBR5H+9K+fChQjlnEksY4QB8a+hTiIGeQ0Jw/1dE98AHZNB4
CC2tsREq6lQowfBqANIzNH47/TZ38s3RKHlUmNORwD+iyHTBcfqhZ6un7lO41hU94ORluCr5VLWb
dl96OUfGgmeCwP//EdzMMzg5AmKrpXRr7c+xba18NN/jQkJoDW+py1NWAGfznDyxVNPaZhY7WasU
zDC0d1+FhXss+sc9Mm56uruyWfHlg4k6J8SYRKY4qOQjHg7K7PrPzFEpyYcEXn22bX9D1xi3LLLO
gKisms6T9dQ6dy2LeOWIcPEpIukkpLdTzOde9mWvbnrw0w0MR+IzZU0sbiBT9zKMOb0SEQzCV7e1
wqdOwWTDR6QMu5YOyfLhdPdvA1jsL28JsK/xS/WKB53H8C1pL828bUC9Cf6VCrle9QsCM2BWxuqv
xEbSagt32BaHN8Bh/tM+fNhFRfE7jFMIAFhn2pVCt085X52ybY5A+LRIEE5qLIvvMb0Mw76O3nBw
d+LS8mEyQolooiMHzRnkPNTIHzL9eRAWB7KNXkJ+na8BYrkBsI+cfiDKBybrtppUmEHJtu9kgX2g
lcNhZe6uaoVnbc/SA4mj8N6/0ZXbSeJ0dA2Q/ofnGHsX6wsfbZkgtd9PdsaSdm36EpJSK4hl3xGD
MTPGVzfBclL7IhmLxcxumEyxc9XXkUle/MzW8uo7ZpdZHIjOXFHvaNIWSJbqNz8Hn/F0xyAfpn16
y0NrdkwTgkUhjZKHmAhA3B2zvpUT/WTUP171+hD+0y8I0tVM/RC9KVlZq1GzqrJvOy8IgPIDHT11
8/i1EYcgsv+T2Ez+JJTePyjpb1JzFlaW075sZQjivPucwGJMxByroCx+GDppPpTTzs56TXB97/TM
ATehazNd4hN2ZI+eFNKKC2q1zZ+MH3YW9/H5Z6FcyCl9N+xQ0L0itA15trwCntqMuC05lrmMw5qI
TS9S9gYvJcnSXeQyDjffCmonrQqkESa/9QvIj4sPmo7LFRbENUSEHiYUBEuKMtfcgoZZnaxXT42H
rjenQfPH3zhKoOS17NBB2iFpiOLC7ehJ8FgvdBMV58PB770IPYpJlbhJmJddSiwfi6ar6ObCJV33
j9K3QlwD+Bwjda++f0HjWhUUy6zauTObUPKZbQy0Gc4kJGWKMUYpV1dn0xzE0GjgTHML4cOSXg5r
yD18omOD/FbWlFqoH/Alcu60tqJUOGk+2L81GbCQA8JFXlA0ffxxJQaJCtdYE2s0Ui2juBsWlQnc
b6nHaEjKGw5MtOkMDwgoJScv2diaKVKcFJU16nwAEL30JzJqp4fWLL+NuvlMjjNbmFWaVGhpchE8
Yyo+joqfTbzciNbUwSGvblCzUZplwPEaHHmnt23WdpKfNWL/sNl+fnm5PKg5NGF6iEugCEQS2ccc
7jjrRuYc+c1u/lydvxi16zKjTQm3/cfe+32/MEGIG+gJPtO0BndkZ04YNrqUV80OZ/F7uZ3ub90H
yMX6hwUFvnu0/VcdNUQG/j/dG+npnX4TfomDgYyxabsEorsMGmIHd+4S3Tlfyi7oKruskC7he/2h
0zw16YvnieanW+c1I380sWcGxzke5ScQAZlcG3Pfu9KFcdYjIodYqEn5HTjU5ubf15n7KXq2pRXi
y51kjP36/IsaKCnZy7RXhIbfExrILJ78pPULukIz9boNx071X4zFFjoCrKW+NJt/FtpKMzNP7LPT
/DhWFtLO+/utCl2f+vJ6FE13JPP7bd5CyGW2v5x5wL2jzG7f1exG7YJDDmSKb3/4BgmF86aBomW/
dJXPwsMXdAdIGHLU+PE6IDe8vG0gxoAJ5fWehmhc69CbhdHUFq+Cn1k52Uq31ekNFTUAulQ/7vXX
4A+3muz31BvAqStj1NBM/TF+8ljIvb8+VfimN26swhVXjcU/Gu9NCAnXjUHA4j8LwTgyUChvP6nI
sJ1NjsdLZpe3QG6AGd2zMCz+pf6L/VeSKxK1K+TBbDGJNLFfZhvO4LZOiJk3qBZyQfVR/1RkQ9k5
nrisQTWWpqyFnYU3cJIIKws0MzHTakhgnaaDtwPKAXvlsul7WxwCg50pElNIKz0/qG3IJpMSu+IX
B+YBl5Ws12AyadHYbPCttZXreGNgBVjmcahKSONx31v2KfpJrJxgQY/E+V+p7fhd67960WnugvJm
ka5ynTkhdMjLYK+Hq5S5fqE5tzYwp84SV8NFdbO/mzxg+p70WI8BmK1XtJQ5w5erGgz285a8hcoF
Xs4JQWlPtqEdTOxaYh26IFkLDT+TcjSXFQa25/YHc3DvUycEVAjdfbaitXItwhUlVhAbrltLzCCt
UlamPSlI8s0nbJNi+pgOSSpvw4tyJslEU2rkFBm4KFMljxZbsfqU6A/OB+XK7cXRaFMXfImow4eF
b5pVMukj4ShTIcM3EApI4PJJSi/dkpYbMvRh1zHSvTz6MBMe2+PyLolFHvouEgAn7/23pNqmM34l
gqOQcesAl62FsPGFz8OB7WDyv5FZkMKHBIsfA7qMBdH+jQzepTuFwWh4LPe1Xl9ILKehG5ZboNEJ
gNmCQnQh8IthVPcJTG45eCKV0YZ3+/VXJutV1iMcg75t0lyg40Ztv9HAPmDn7AXT08mkXNze3ClW
q9tZ4MXtKy+EIZsXWQH+mpLq/wupEO7e2pvEfXVe29HjFuTrSKOWjxsu3qZexvRd9+/MK3Gy1ziz
5iGsmnzXMZI118z7jzUGL3Pe+SI5/EOUuL7S8tbOPvdx7tSmHQvr5pLAamCk5dWnSeCtPrnfPTiA
mY9ZH9XXDxFkc3azeqiHGcBYqDY4Tkz3KpXIdI8pGiwxEYYsdGZL2eC1QosujvC5oW3g57F+lBN0
xNuWLgq5G4f555txNx4vM+G1QeHfHgBrdkIzfvyFMekWAD1ktpRePPfGl1tRrL/wAz3Jyi0lY9bS
GxOduC5oEROXrvKJT4ZHyCrNGnqlC88ZpBUdW6lPHALikH8CyO0jsLPXvUqgL/MTRVLENlAr2NZy
l+ikJgQtabM5VrK8wu8s/G/67WlmF1EFcNRsfJqOe3+KS/DS/lAGnYRRtjeFtm6Juy/Ju4ur2vCL
O+SGEzr8vcAwoS0CWVvf8ZIDQ6c9l+kayrfoPLEjCpMvUBmrjBQTeLIgXe9YMXYdHqQ2RKd27bpQ
DWpBEsWa3wxbqOSmBvQuz8TUsOSL78O4D+lNP2CdqxtTi5kIN0X8KZsJ4qO6oSt7Ix+h9O5zfxa9
kF665cJramWCkNhwygRmcfM3Qm/7GzYSvGfJGxxKyKqAgjBeI77ETrjHHd2yv9pZrIDJsrio/6kk
3dmnsmkBST7CBgPDtNK9+HTUwagGzq/hopfGelj31bavsGSZK2AH9CEcvJ87RPJrqGSO4qepmFwS
APP2O1/SG7GjWEe4kgKDtslu93gMjoDN8oFea3sQ3x6470IF8TCnr/VkFJBcgji86t7zZI7IlqUg
gV689BI+5X3N4f1edDY4R1IBZJ0I+uHpgdDrk+zFfR1Ah8hXDCg56strT/F+TGwu7O3x2XC3I3z1
Fl9tGm1Ne9V5iULIYqZu6q8vsnU2e+hs6Rm37iSaYD3N7UuN356BVMH5U6IrWQv4qjKKIzpOvMh+
/+V2pyEibKAYrmesl3RSxx1ULC1NL1jdCIaF/l80WRJI0qHY8qRiFf8ctMfgsqOQJXA423ydgI6Y
rx8znqbor3iwtqQ+DfLh8BMXaBBIZTkQJp97dI9gIYe6o6rmZkeYIWLLbB1EZpYZdIDx8Gr/NdE6
+/rVPfzYwt0iSB2ADNhMjbjpc6Db6S5BaSF9fZ7P7M8VgwM/jbe8mwW0wRD2qQ642qfdHmByL5FA
QNbilmv+GNWFkhLLvTVmm4xMSRMA5Wv+JcOYNmXbxQrTJaPBUC5ZMuYWmvH5dsuVW8dnkL9zhUl2
X+8EOavIPFq/MLIeINMySyEC2iJsk4XgL5XHXjVuyYN8x59MsJX2P38hjoidYMpmfOYCBYzgL5dA
Bdn9up3MXDucc3ASTO85I2+2URfMVrUxKvV2oeAHYor7enhktVYy8vp6FmL2+zfBSMCTh4ceMbXh
vvlufmTdVOAC2p+O/eFLmizTUCEdl2YRCTS5sIHrrwoz2nnZTjwY4wxgdYpHfTMwH3WFfKDW5D/X
K9hH/MuIy1oIpr/Ep//WYKNn3VP5B6poGdyX31PJL/1zO5z4Hpcz3sjzl+ki3eT/LpCano+zYOvu
worboNYcrINWn5ZJvodOtWfzzEdPVazC0l4GWbk9nbbti+7UJ/kj1vy0079jYy3KxWtUuf7QeXe0
x74Ab/WwHyFjlARkmaFEkZ3HdI9M6n89C2ZR87lr4CFl4OgSaifHknvD8BS/C5G38WnekYm8/7IV
18BRsa1zwwMKTOrsA+iOjx9/F8Gpj2SuMhACnqpBBdgxCuU/T5xJ9wMZSWgY1x2Gc7dgipoezJC+
y+LS2pFhTT1YpjEMoz4TglTtOK6PDnwiGyHAX8jL/4B219X57QMGwvDf+T0vLIcMkxq/K+P4Oxhy
Vvs8pcEdY3KDVcB9OiND5rgbexWwxQrfdoMwCRzrkzcnLmlrW0Bh110RPDis4aOtuv2ouF9MJ1Co
1dQ/8a0SvvVUD8IlYhjE10lP51iXZEn5zqESqmiTeaMlL+HrDbaNtMhTBNwwblCrcalgFfN2aszf
UdRE4SfFGO/fVt6Rjquu7b+WyPLo4xHkMMOCCi1F8ePABLQWrjfOXYWxRJlpbaaHZxxUPBHkFAso
kNoNo+RdqcD4fntiMDmPbV7FroMgprxOVgSE+yE5AfLMlgIna4DUH/y6Z4BEzLifn2gMYsuafJg9
XgWwWXTdEezbnyZLOvCz/K+N0oBih9UqtPX9ACjCbj5LH1buUKT4jQjGTxQdtS2wtM0mXgxM/PbE
MDNfMBdreIcMauSIGRfPBEo6FlKoFrwL4UHMUP4FCVKjlaGK4wXNcn/v0vP/A6vekR0CU34tJTif
vypfWnRcZ844kEIUxpf7sqPwYAir0UkJiOH+c37afKJ0pA/9/jMu23YgGMXdRXHlDVYx/vy36zjV
JbLWMjjEUZxEM0ukaJXFm+S7zZaZRjNCYYXZVIICiPzTqUr1rtjMt4dgPHxWqPC56oAnnJI6oljB
dBB9sk15LsQwBfLUnidKsCUQ7i4XrRUhqdL/fh1lMMmTY61NqSJIGa7Wqi6rT0xTXr7WsS8NDXQe
KaZkWw3QUlHuVDClCRV/ittXZw8tdpsz99sc5bi/Toq7lD3QmzmVZGXTAmnCRdG4L7qGYOf601Lj
dhR5/S5YKME9Tpf1PInZ5bNEuTbwBraKtjPUflIoc/WNEVlkuQpJn4MXfH2c5piah1yYFj6GVEZK
I9pzXLpj9gGgz5A8uDB+OQ58rWMwvr+zFyI2vL10cjK2GqX3uneQ9yq2Z9hFN8CVjDHHJaY8FmZj
c3D2yM7pcgVgZPn9Cjt5h/DFYVlfLtDZrpQJsJLSVNP9nYa95RcmejXOB+fml6TjpfyvsnSUrPH8
6C2/OQyNVYcTkdUry6U43QE9d3wyTnR0TZqjmO6iHuQ4nmqQavYNHGQj6AqI7wuet9dN5+jLaiJT
FZzoZeX0UKXg56kGODh51r3ywICU/PTE8A68gjfRwg1Bmjy85lmlkv+FfSdJsusVGCpjpA8K0GXk
TgeDRoQqVspUFqGDRUz9ghSfeohaiHepKg0N27vF8fYrjCvoNSOCvImg1lRwlcCNjSkfLfLQz8/j
KaSgJzuVi4XFOP7XcYCqnMeRVTIwwMXuWN/vopfaOLjibeywj2BFEhko/UP0IvYZZHOXlWjd1wNU
JHsa6ZVZ7SnyIP+y5GZEDKEPje04TxLDO/uTj6FrqP8U+KedW0Rbt1dK0GwRRDQstdOHBb6XwNgA
g/46szXi3GWjM117RWWSsFQsEZDU0JJ0efX7DbjHa81+YOa4L9XrszbUMYZ/lid6OaWodu+RfE0R
e1mGOo/3rvCZ+m6TC8seqtLJktarlYiuab5pj/H8x0SAn5FuCikgL4aGWEdGEkv7DZR0J5zayikF
zq7q3ZtNY8qlDpHJ3RgW/aTLCz/h8KqfIMaje4kUznfLPGQibACr30G2cDd8Va1nTnLddy238S7G
D1707Yz+dhqMG7ewnbJLaXykk1phITr+GMg6u8Bq4oBSETviWGHzA6Gco6IRiFKchywsSIg+02GM
o3jlciZShDvkZPUtgP4Kxy+Mpxy/BrPLfF9Prjht/Dgzj5KRkzjh0CBMLNOIQdXYfcqziVLdbXtq
8M/9F9vzkpJ8qX60ZqO6Vjh5a5qYEq7TETe75SfQ1LINhqsgR+91CsPAd0Y8HYkPXbhMtABWoSjX
qqo3JI2W3gAVsCS9i0W6UunyEn1bg+7REh/Nh5ZxBA50xa5uwbcipZZ37M92LcX5FBMNzWE7gTCW
PPzCsUZs+tTXM6OcFX1fKU8CYDYATD2/v+hF/P19Zmsl1oh0M7mDVsOpUacCbOenZAW5CPSLuRrV
/0Ov+culhqh22/SXg6u3LTwcTHDcDTlcER57vWrXAF6+/uJobqQdhL/zgBF6+/JXyBNpHrA4878w
Ac6zzDqNdHBBUeAVfYFrpMikg2GNgTkEEPmOaN8T1Ol9T0uMucCD52frUWgNH62OBq9M6PCtD0Q4
G+2gb/aT5Tw78HMz6vz8Nz2hBlvui0ohIF+U4idg4/v8BKtxrRQr7IQPbwwHv6LPJgSCIEE3vFKF
xykrDSXzR9V7stqxnvLmdN/GIkpfa6hv2Bb/USvwyzvB+I6B3V59Idyoce+mp8XhS1tFQQ713Tzm
Xl4IO7ZBT+tQzvBogahOhVV8fHxJylLU+C3n8xDv0R1mLuTpH3w3EO2Hf4Zq9Mo3Ex2RADz7fHgY
JtTFEmE4ofASY7wIDAK1T7oqDeupK7QFtIZBd81rLvGnoLQs0DJoOzTbglpopKZsMEAt7KuIa6/n
5MbeqTKiZ5TRX3GulD33VBKjymp/n2Dtg+vfvfb/ldvngwcZibb7zwBHOzW8l+5CZVkrMT+tLdBR
nyCBLceJS0Q9olWt4sp7udSIaSpivCsTNq7Yns1g9alecSiNIOknasLzrqE58KWuInYq05er8DjQ
Yjv/FiWA6R1UDhXHA+/bwl3O9iGRSyyFLPxtd8LKjWNZsKAYK9N9KjY/BkPY1qMq/+A+TjFInL1V
rX8q7mHNMx1Xzhz416xSvr8+vLECSHqH2L9VSjdRVxSlix9gUIEdFYG11oYJLqpJaPZWTMtnAPYs
hZ5rJnL52yKBu0yRs79pVSRp/DrNqu+08CrguT/QcxSsJXOBySz9Yqn7rwpRUoayCJO8n3N3Q39J
OxV0xjI6Z7V6nP5ZhaK9Si1fbxboIlmwa6973SrIi9GQ/chocfn7pzErgDwVJDP7VybWNKeMpEKF
FIRzCGa6/HDjaQeEkbuJZREqj2t/4FJIFm62HfnVWvJwzWeVHDrIZlvMzV8j/T/38R4ZbEjcgvSU
CcHc3G4KbbkQBbQPA3yv9UkxEl2yXiI8KXnCelC21Y9wwl4NZk4wHLSMr3c3jKVva/H0DRiTB8sj
OKJLr/JAbY93IftWHhl3bX2uQ5EKAG2NkXz8yoEOQGPhzd1HiNjjg7RO0LRr+ewfr2xbREh6pr4x
bl6yTqzmiWyeqR25P1GtC09sX+u/nXxKzrDx7Hx6AJTwajmQqJia8ais37wwFQAPvBzlrTGO2e6q
ZTu77uQuIliuQzzO+hyJbmUw0DwnDpFvklJQhrtVla7Q74uSJI4VrapxIZzW1zzpJKpeeM3a/OiO
Wx9e7C80FK9SRc3MN9GCzuGQ5xr7zVHtBGYThZTiCjsBNQyWWaaH5LIhynvjGtTKdCVbt9484c7D
+Dn1CFlenJPZpFQa5N5g3Kd84Ekx8nv9ETM6Kz4LRwf46oXGGGpF3fdwAsSjALiq1fdgKbekd1d/
rAPX3WgJ0D3QPOzTC4NRSMPRfaO04INI8MX0qbwIcZApYSJk35MR4Nop+rtxbhgaJpvwhdWBkp4A
wubkl00WFn8NBpCHW/N7JrVbEifp7EZ6Q5+L9qRfLseLuxBUMhJhe+H2fLITqDI+MY6QGjx4t3u4
BCQLuOeMSUvsD7vRtzr6/YwRaEnivrZE9tYLtwHNE6pcvq+e3VilGry2V6lcjqtcLMTZaVqq3dNz
qdb2oMt+NPX6okoO0I7SPKWJwybNauikTuI3du+dYe4Xor0eihGTuuBogIOkuAefWuqtqWMlEimS
OLsQZ1dg7/TJrNqvDEkE6Q7Cb8bUr0TPaDC3k0zloPcMXcOEM02gY7ZnXoKHg7XFGXa1nFLazG8l
LOwqHjuPeCp5mV45DVfBF3rksEpbtW/doctolqm+oUYrFQc9YleUibI+48BL4v45YM0i0prd4NdK
DLJYvehFUbMCXMzgRPydAU3Y5WUZKqM9Ee6thugKhq77WHfqPqJJTnVU3rjOyz0RW2pIFVDqiW/0
MisTgvXqZW5mFd6ni2Js3OYEPO0QzAS7N5nAxCwJD6QjiEd0hqTeUYCiXP52bfneTzTdwScIr2sK
0cwtcLzpM5c/89tih0iL/lDpm+Q+pua25AwB1kNitMGeVI8E6bXXNmTqmuT1pm5GYn9/57zMO+6g
FRVgxgbTEolRMdjAel0nswrcHaXFxBWyIIgz5zO5fj48RkkGXk2W5CUPSX2d28bofYVYDO8Lfqhr
i4FB0t2keUxJs8G5DGN4YF1XVw97V/DiQVzke1yFReafKwBjyJtetR31UAiLZt9Ut0OdYiJZ6MYB
2RqF7Be8B3fxAp4nfOjP9FckWfzTAu/fHLMrdciKSqEXlcR9CnwTkLXiNeR/S+k917USTCtpzlgk
GPhYeWK1Q73zTg6EG62pyIrpB8KkjzYVijf03C+HqYR9x5eDAS+rtprYbiETxuz7YMT/2UpfNcj3
HEcsT4KGLVK3u9acv7nHtZs+w1GNANWIfzzo+fSQq7dKRulYhN8vnbMMCMxwr8LT2vRqCOwsQLpD
OMZHt1Vn9dGJigEViLgg1iAAVTT83GI4WHQtKESx5lrC4z90fGR/nWiE1uRqjllduA/mPw0c3Sae
YREnqrDwztNG44KknT+azbLLKBa/YXYkRsQ8FvGVJClQn5Oi5gkOwQhJQBeAkM7C/g4RvC4d78Qk
BkQh9rgbuuteEQ2COGLahRDg+jKdXMsFVVTOFrRUl0bQ3lfB1LzLzuko8M8RNDuOSUe+/hVCke7z
Cbqcd9sJ9X1JVwuCGhzNvqLZvxngA5hzy994D8KZxb2tmLafaA6bXKJwY78Ph9AfSBGaLol2+6hI
jzqVDhSBeFs6FWfQ8fPbVPSRwX2s5wlkWPtZW6sqZEt5ZKBs7eGWxuki85wgtdArwobFmCHrLzH9
0ZqIadlcs09JtTMG4hXvJ8FrwB4nonYtHUWbi1ALf8avek8jQWCeSIbAXbsHmfxkPG1wFX5reu0O
UjIvUqNU4tkE/Dfxe0EYAfJw0yklen28h4xqOOCF8MVpXBv1xXish/VIMGB3QMVsK51CHBUwCfEI
zOcPD6A1GLKZpPeNWmCEz9nTGdknUgMpZXOqeMLdcCg4T4TnlkTgfks4MEhHQlkeWUqV+sGTq2ER
YJ4yTs3WSnS4SiRffi8sxucoBsgzcbxyYXzhR0O9ZKh4nN2MoGzKWE2mOR/98Zg9Pe0px5fLsGhT
s21dRZgB5ZzEeZ3zbLdYFJaIhuvJW206qUYqsEsYa9puJtPvmYYsjrdgZc98jZcnewvgTtQtzYPJ
sxandV6MLiEsJWVcMyxnkTUB3KMwW2NvLuGqBBdTmDpFlZyF5PTGE8DVNVeV4Qe88mUV1oiKwznk
ozG01ZB4gU+Q5jbKTq0drLKoTSQ/bVWwWul8xLGZdr995ig18t6VVmhK310ZV8WnrMLQ7pPyaGlE
41/i5TgZlVGBcj6z6emlrNC8IrSeOux7RLPK7/lQV0Bf2nanRMWRmXdxsxm7EqOmkMC1hRoUq4/T
p9NGGxRcn6Wt23mvlIUe5U7vY+89Bo0GZKVtbx9KOjKWQ80o/nUxIbc72zs2suhTStJ4a12MuHuD
L/KEQmPNJjzBb6xv+DRbe+oqGxPGQzTK6qN08U/GU7JOKkOu1WZgbGVFgZkI2l2pMmQV25r1bgQp
P6cJhZ35gU5gDoebJmVCLA6EBWcnmpy4VajOSFaHEeEl1yHHGdEj9lGcCveLBEtRDCL9ZkUxk+3x
NVeiMDJg5Snz8LX2XwELQcupuBluDUFzJJ12xksBxqxO2aWmHwh1p5txlUsodHb+p3pmTQmtYyS5
3dsYQvUNRIb15N4tvN503huc1kiZhmGoVTLSX47G9CfEgY2SfdKr4snKy7UQgrSKSoOq1oV+NmuL
LaIdm2xxmfsUIeBAI6NvnUYAXWDOV6aaMXPSIoYPNAYoaYG4w6D2H8lA00q+lKTqVYkJtlYd04z6
VTM6Hy3iqxkTJYcV+eC+D1LSBeU/55Kwso10dg6eS92IKM9xxoU7jqbt6HQ/X60eUwcitDzg5Fz4
4YmR3chrTK3eD2S5tkoOulRdZCbz6Ojf6RznJoNEyjBZfNl0QFR2wAWHIJ9Q0oJ1Qhj7CqDTJ774
PvFUFBRugd+ldUVADX/qJKD81SnYO14i/YJrIEDJiydoYZeD/WfoZZYP/CIyQSnfT4MXhPLtWeWQ
+VSlg4574xEmdKg+SGdoU7RCqEESwFONB+0hoMHg9u6Z8Gt5oZVJ1MwgAgJSjioWyH0sDWXv1Sn6
XWGEm0AhtFuDTDTQu4yDpSp9j2iOWehRr5fYCacjASpXt/UO1rokRQp1wfj0B27uT3gKNU2Ic2/M
8wcqItikK2PGatPpAKo5OLWAHAQwkA9qc/zd+9idlTzfT7Up+c7gLrNet8QWUXiPdcx0CCmUIH18
cmcK8GIzNIwRTySPGfH6Kcp9JKOJc45iEKycp5OFxcaTtrPPPFdjj/I7jJ3RgzCgiY7SFK1RyQbi
kmqF/kBn6aBHuAM1n6YY8dv5rEuBzpLiIa04AGCgjhblXervq8FnlC8WbgzSQZ0j6YRKhs/f5SNU
L77CqTBgThuwsJ1cAwvxTAdltU1WOwcySyDb96ODY72IF413NBALrye0LP4luf5dPRSR4fbHDm6x
AQQQRwwK109tii2z4wA5/+LlRppGk29sWz9/7jCJ6vJ4kX7lEIuoA6Fz0JzSYLbgMn47AhadY/3v
R/PKIjzFs2b2553eqRPKmFpDoWjCyG/7+dRejm1BjVYj05yJmTLdsvQz/pMHO0+H25HFyeSNDxWH
eZfbiwCop+GAX+276fhxhS48Y4WNb+JyfayVV/zbAunI5Gu4upDKhzqlBhERjlFNd3y0k6S/AAke
VDG1Uflay2AA76qEkNcpHgy8DHUZqwU2CuoYiNaNSHuhPH0ewHoV7wFxRhGwOcrItOtdtklpL7Qy
lxD7MC6ocrPkeNRAPq0ChsIgq3K9gHRFUlQedXHxVhPDWrY9QqfbHByE6hKctIz7ixEmeWuGtHIs
mGdA55BrFv/TUlRG3FqIi3NdlyV0LGMwG17ExrctwvOOxvN0Iv6yCHI8o1RZF/+h9G9sSGgUQBk9
azZVZAxcHbTLcZ8sz+rp1o1DukBSauQyxT91YHLPXo/0BIEyJgna+8nqTWhsyNWwlg9zWy5dDIqI
CDQL5HX7RmPDtVF7kTFSW9pOjlQ4ouUXgQL9dvcTCWdRw0X7LUpkDrdG8vNQvARkmXHvJojfanJZ
lDKXpmYQk/WIAdUp1qG1wpApoOZvu0kSjCwszoJN++SWxscE8XxPYKbCOnxFkJwP4r5n7cqr4Kxc
rB7Nr1/ZMZKEnhZT+2/K9gXVfK3jA/BavUCgboBq/YxdGApQH1xnuM2TrFA1ErQtJbjo/XS4dGOs
23OGJiXrP1jVIJJbx2XHlFziVyNMyeQ4Aw6O+6SpV5uzouzSAVPKoAp0+OBi0UZ22jzeiGTDKJZI
MoAses3NZdtJrTdRicLkorpsWreleOG0lsT+h88hXdOW7wsQ4D7ZSwSoCL7anj1bmocRVXe9kT0Z
EJacaM3YX1vTkl4oSJy78UHrGWMz7OdBzRdIIgBo+e0DIukicF0GJuyNxnzPpbrX4sQDde/+4aPa
iYjx7XzZnJ0hFrwfmM3FavwKLWj5ynJdrsFstWwHhFwpYmfYgblo50Yi+rRj5ychn0SLfdU3KoVI
k5wq6UiXj7SWwLXapyWxKeVVrsxUEdQXDcTeXVxU4H7T3eh0bGbbNuNH1FsBODBTqItb9KAJx6uS
ftKoCifDNO0xqfxpfLI9sGqq42QZCsa+8zBkoeBjpqMrff7GiKsdffCogjXZVa7K9++pYLwapyvy
6sCEg+19oQ1o/umZoHvom172vA0WAvFncF6M/JHNjTSsBqahKtLc6x5CCyY2uexJeH9oN2nQe+lO
sENSOLkSb1mjgUYrPhEn6CRKZ+WVddeL2leXOIpUNgCBfI/lZxO7QceymKK5wSQHJGFF8Y4ovup7
bU/0rCj+Hj30GUnMhBbtcX4ZBW6eM18zrGIlAt8Zf1lIZZtvuD794m/k9hhmwyks7QTG/c6rVkpc
wg/z7X730gs/LJ+InWh8fEz8UgOaOOKY+t40FRTuVrqhdCBcCuWTbYW+ToKC5R74mydQNDXh5kNF
vLeiJs18SyI3i59jB6W7ebrkL5cr40T7BzhjiBbpkslgqXn/lgUEQj2QBVqybqVleUrJSvPK0l5M
nwkgMhEXGtSXVrhUjesZ89ud/xT+yT6vO0CNIQjavAic6Y8uFMCNAwnS+A9o24V9cGKrNSSS7vE6
aXwB+hVdn+R/Pp1xp2ukuK3VjSc9P4a71+oS0kdOrtlcng5eRgqMqPxC7czCKKOadmj8iQP0h7th
nrQfPmvQleUdIXvnr1vPAAha/pWdDwaXFOOOBilc7pk813LzykykKk9GU36fg8Ctm+bJQRGcKlzb
8B5J1fzQmTFZZqwHKn/bOiUJaya2mPOVhafqZ45lDcIZsaTctzkmxRTAiBi8w8XA9/7Jl0nFTTBw
l6GAYZUOuqgu3qkW+7fUVRWyNCa26/eh2TSuC6iCQC5VWrCiyRU+ea2GIeofAq4yJuSJI0KjfJjq
Au+2A1tgC/zpbWN8Ahq0YZDlm5ZAoMlKoYj+J/zUJmwatuGevOyfudeofNKX5azlqapTVKKnYoMT
2q18t4i6ItL3w69d1D8B+6rYGzH433B3Fh1wQ+uuK5NmVLVhMvadk7i4QU6wVR9/I7Kt+a5P7iFS
ozXDza0w2ff/MXGkOojBBZ6tU8lEHjswl0CAqQNLUhEDjv/tYuA3dXXMAb/zjCHj/Pr6brRl1Zyn
1cjC7aY+nOkDNkUjDNggg51O1XCM3rZZJURQ9Aj67507CROoPNsh2s89ilyWfm+IGf1kOixvHMvT
QKDxuLX2AiyQjUEb/2CZxS1B6N2qnN6y4iDrIbaDQR2hzozT/cpAlHPkY+HwkoMxULXqWjDWOBpY
BqVcZJukMg25f/7bZvljoCFmV9tdoHePpN7o1V0xb7KZF2LkK2dwRYnmmOr4UviVtWTT1Qt2nD4u
09duKgPZkTwwpJeMgudKj3rJRCP98onAVL5fW5i30VMemejlkoSscGqLhcb430v0MOQWbzGc7lmP
bK+mn0d0d8g+AnIsVmAAyKhgEkNH8JU0kYQObE95Ti21Eg6fJItcg2lv61ATvXa6jZ05pcaABm45
X46KC7R/up7dxI7LK6zSrQvDptyl5xW7ko5bsctzET3u7koi09H2Yizbzo8tvoJTvVN0wRlxqQTy
7tVmaKapsYcPRHQt/sT8BdcWtcWqCSRs7vuUpY+m3HCkUZkjBkgBaF+q+2Ihq/zlq12mMBAba2Nt
7O8GxuWn8kR6hM8X3hZCA+zMAMTnvqEj96TpnR1UVs+Aw21IShwuAYIvUcTyfVCLuO5NMlgBVvhx
tAxET6Hq0e6jawR/3CcDiUMXftRLAexpxlKMA/2gz1/Ciczzu8dvzEq9X/H2S/hemqm69WVpDe5P
Mooq1YnLQKooyIBV3IiAzxUx3LZhpHpWtQB+x0Rqwf0ZZie/nQszR+S4tGEGPLjRm+CNKs3sQ/Kg
4xKeq73LNfV1WxcpLGFXG1/GIaN5syGkPCejdwE0dH3AyNo25IhtmEgQE/dtv/oyeqf9MXi7aHSb
eJEYNLgeYbvq6KGIIMO8REm3923+4gxO64Ju9dypp5InBckTlEY0PDpDwgEpqTGHbM6c4H+f6o1f
6r9s9KScDBqbg38YTgTaWV/emar9NEVGxbSNH4Ok9ErOxnPA2AVC8BLk9qsJpggrodzcXLfifaZT
IcQm3zLoY1bHV5unebT2hV8w+/pNutJx9aIicpUTIYSGcl8aT8zxiC2jhiv4hMmUNWhcB6BApMdT
SoRBuxVP5VUTgU8/3470oRVFQUbWsEiIhJHE/whNeT2De4MyhDrhww9kr5HSaqDKmR2ohCT6q0E3
Y1YBS4AHe7uLSiDbJhjvv1H41JJK9/O44W49Bv2Ks5TYHTfTVaeYakG6Hz6vQrpRjC1xh28wzZ/L
og0bJDASd33RV4GFHmDqOTUyU+uW5GRDDIYS27e5ElCEp6V4SQHIDTUJ0i3A4GNa7TC8yrhVCYSZ
Oq/s0xzh9mSJ33myXwlPhg/HtYpulL92dgRvUz/SQOVspV8oexVnyqUFOb7G0sOcayBdvswQQ7Up
s45eXm3GMey74Dh4xHPnGFxIdd5aWn7uSL/8/1RVMKhdXSqxSsRyOo+ALCyVMuv1IW3YfRe9c1YP
TBpVf32Ux/kYMpw4/aeM3EeR4Q+2YCBfys3LhBNT8y43lUxjTR1y3AXHgegzixPFasJ97+1qmiBk
vspYlRA3AVekh30iqnLmQAH/jKl+dC6HdIPtBuTnnIDiDs9C7r0FVutQbnaqsxwmInUxTKxQ4t/w
VxpCiZVlp+RfrV4ncLOeqeyAyDRBh/XhlvHQ1D+Vk2w8r77DoE4ZWGaUsN+AUMt/hSpI3oQ9Qs9b
4T0fBMqHf3zjupIogg4rx8lmpGoLB8C2LTI9AcoO/MwI7cIgQbtSaoF8ScZHR49tNJScHSjdJxAl
65/gJvmXHosn3rps7DMRlpur/byklWPuaPNms4Bb5UABDcUq7KzV5rW4N32VC7xezXj6RWSO6fEd
O8j6Tl74zlL/mx7HP131fDaJci61qoIzImagQoVm2cvL3UADMsMynKGQ4Yup0B+EmwwGLCedUrJG
K3BS5h+XB4gWWmDHFxT3hoa4+wQJMapewV6M5h4Af1tauamYwQ4Bb2dPHNtu015TU9nXR1K5ToXF
rUNAyIueZfqPyoOGz2juk4AOh6q4EKaGrN24AJQh65X1xsz3GpEBV59cxQj7zx/dZS0R4Qfkk9Xr
3JNBhmEAEogFQXnZQ1e3O/PiyHhi1H6Ljs2ZVKP7EkvATJfC3pPQBF2zY9Mp+5kI8bqiQHwnHc3k
jHgdRQ/koCRZhlcAg7BdtrXaMvXWLpU68mVLbql2jbNWIP6zntxQS49oonUXBzTk1YdWlUCbID9z
ppwHUIy2K+95irfzCyDdYGuc+9YoVdH4xqPXaCnicPK/Kl2uK/1aFxYFhPaqXSO6OaCK0YmsZgJK
VE7N8A15rtTTVVMAdMwimFVUFXMkW6D+/n+lUnZOhAWo2/YmqQ5lhwDwmMtlfywKf91ZtRdOp63E
Mwk2quppIENkBQraN3eLWwXni/FWbiiB5eXPncUVUgHO0DqAfPN6m8oOt14NfKLQ0Rft1FoAn1CM
Z/c6WMOKYHAykmVlgu9NACIJPtKrLYH4jkEFxAY1HHxwvv8U+S6RYGhL0sn8iVkXmJhuErrzX8sw
5e6TEN5tjp5rml+BbzmKs87nLxNWxs9u3os5PE7wc3s3cngcPNF0ta8kAQNnEC3MH/aOw1zwxyO0
7u5TN+gvGJjcd7VeCxoYNKBcRm9n2i6Bv3Yp/4MmLjmp0JuBvphgO9EQ8tDdc4dfKS4lgT0ExFXL
Na4RS3h2jyATZTQ2omYfppInsOWb7MwvjPP2VsUlHzg6aVaRjLgsrqnOVw0qFzr2s30QQgM9oO8m
YZ/WQ6SgDcB2yogbumD0wu9taMe+0+AKDljs4LfAL+h6V4ne1HRi8/+ePFpWdQiYe0BFm7X7fAYB
CPxCUSVe5sJRp06Cf/6Nf/P4uwjGISY/Dn9ZxGJgzvSiW10bwv3DNWdvX5n5l4kJhVvB5E15RMVj
VPpky+4xwTzvW7gEwXXqsGOPqONy8KYTsWDaPbPc75bB0wN4vkSBYgy5tZNgdRNZ6kH3OhB7CRu6
kECLNDxrYlQhFVYPw6S7NDvF3eT2B12jGquOLslSurIqKRlOujVXMej3R2TppLaFhZUWZU8m+/a1
Pk4Od8xrKxsn5AVFOs97dqBgYakxMGtZ+YvQp5PQ66CRGn2y8HcoKD32PoqSFoGu3MlQQBYVUAmo
LwDWt0owazL0wjYFukn9JuvBfP+Dhssz9bWsPMZZji/tpYl1kLQ6F41X3aKeIMwgbcMBwLFSDUEg
iaUQ/fxjEtRutl9s3A/HG+YPKv0q53AUSW1012YSjxj4idPGCJEkuicGCFoT3CWgMkqBIwtzVvvA
zt5/9YKq12vjQO5jCLsSX9Wb9bTwyamEDmaPbsxsDofTOUw7bI9luBPmZHV6OIKlHa1FU6mOcRwb
d2DO7fzC3DCKUbJeUuDI9BTIXPMop5ZlekQM0qNOyNrso43MKFJCG/0JtapahmoFHS7f5kJiPmEb
pFRUncx6SbGbSuvzQ4LW8nheDsQ4ryMHh7UiCQAdOxCw2ge8jzjSMaMJXlBIAQd6UOhurT55hGaF
hNp+j9OCsNMqmmmMQm+yg/erGEDrEkLlWc5P0xqUawykIpaztIlPRHLXdlLu7itokLiUQQswfo9q
mSMOherPoV3bvQcYUCcUNGNJsyS1Ft7B7yx9Fb9vAXH/D3ZJ4tEDkPX7gTVqox6K6EHB/rXoGvs4
VEKg8qYARMGrLiqRCT8/ZWKM7NluzC/P7bRSp7Y9xtrjecoTpRyRzSQKBn5Hd6mb3+LfkeiAYOlx
6unmjks/hPGUNm0KbBDZs46bKRxD01nIDK54ut1sm49ixZUsw2nf5IPZQN3nCOgrNPKQyo7Jv9zb
honCWLEMrabgSOwQO+o0fBYYe5Afhrz5sCacshzNLAUt/3k5HVVBziPBcdgRfCXCe9Bv2aZMJLaj
vhfF9KCqtanjLrPWsTcpVi01gbyGBxRKxrdIWlTN+zSA+mmRF8tC44Ld/C/bKI9qSjib/UGnVmwA
ZQhUH+WVU03MjKrZoEPO2OVjolxmKgHpmN/SmektqXKAYRBM6EPwCVz6j1bKUFZkMthZNIWTlKFw
SZ6VmZ11UMYMgu1b4w+0JKM3ryHoODi4VrVWsZAluxjMGfdoWRZMH4RGI1UMiFTOimg7rnWKAX9V
Xo4vcs/b9yz5OOI6WcDMftr3W8qaTh76vBEsZbDzVf2qc7y0Gna4UjlX70n8O0hn4s5LxYRHWaLP
Sxc1abJp+afQujekIzfuqVr/bjJhNtM1GbuYvbRSdzkVtpbDxe+0qb4AwIos7HsZk5ASW5MTonxN
4KWyMHkQv0UdS7W+vjeO5pg7IhR77F0kPAGmWa8Yp1C/bh9FrqsIoXvovjdKuxSfFJ7dxjD25PUA
HoA4ChN01VbhCEQqIgerlhBCjE0g1rAG3r0VxKX7DTMZTami8uBhffuIPAb+Li1O5fsXXyBdHoCn
r9DObWCiG5TxuG+L2GGOw6+033ttLGFvBcij8QOXCCF970s4qzGIDXDcHJqxuvU1zacxyB10gDnK
Knq85YUhfCDzTFMOrxbHTjFs0scYMCMuGtlnqw1QGUbfMlCboYlJpOpNhEtgQgovuZN7IizPGC25
huTu+7V1MY/tSbPz4HaBzUuXBFEq8KSnmmwVexsrI9cIemqiHVf4a6w2q5k9MXFVEQ3j0/eynyNJ
3x4x3An3y8gAK87xDIRjout5ATkn8u+pCOdndAO7oFvViGxNnsiVFYt7NPwBQBzvpa+S8Twt/C3k
g7ryGbAzHG5jNQ2B4MncAy9Ovsr5tw6v6FWNGatC6GAvlKmBzgRQIty0+E5Cwki5J8QwpxeLvaNZ
sMG6WDowjp83QfNMxBy+IMSjGsxZNwCyavJNXr/3BpZCp6x2qt4KQjYB3ru5nMdOQYAVBfP06afM
cqpekf7XG86BuEyip9y2bVffWe6Lqj0/OxJNc3O7IEUwji6HRq4/wJJ1Se95aTce1W4fgvGr/+ak
McDEIUCXXIsJFCWBC6spPUK/LPt+0JEAu4pL7OvCHxCoAkkP1/WOp+um+r8z6K9IZIjh3YDSBMDG
6KWunGAhgTYPPAGDkqkO6ehIi29g9ozQ9XIpla3GEiGE/b68pd5irCqxZLcCaOwJPsaAcejOszQj
cR11lz3dYZSZjjg5JBGSVzBn+N67yIGhFQvRgqeRFyqJAaIQleQCw9kLe4DDPd44mAZyfhYkitDl
bDFdAbYnnInuC6hK7bROMb1RnOUkQCXgMDxyRmkgYFag0tYFa2HDQ5Z5zVnxKXb74l2m8Cw4vjQe
tvfXxRdOxWKN+RDcRMYfdFsk09/Sz/xE1R9QNE7V2F1a2RBjHyiDNGuvRZRlTNCxK0GZQTbunYhC
zlAEDvQVMG+LTJUmsyqxYz4zi7KW4eDKbUCEGkjr1CE9NRoz+mr0OienZY2P7AamLg6T1x+Sidb5
V7kDBXW76OZzBOTaZi0YWCq+4X09DiUxUqyQN1q23pEvD9ZD1ylcdHGmQda5oh+uRGdVfEp84SCI
SiM51p14EZcsP/zzS/fm+G+/Q6LNz6orytdzG2xyQ08yp1d0499lMY+C1n2OoTlvxwPKuZnp0aUm
cg4TtmtyYXlt48/V98PX/CZ12rcSPk0SHdpqPqdIXAkrghNqi3hWzORORZSQxjtHUj8c+ERPZpnB
mw+wovWfOdmihhhrbxPIkJeJbX3ucuZrB0Wg1J+qYq+uBjQ+3ZO5VepFXzNa1NDFuAOWsG9TyNl+
3Smqg/I+cCuGLYt9b8SYkcEuxCQ4rSJ7aIHobdzMhMGZyOzs/yKbelLQ/9Hu265pyU/xlaUHzPMV
VLiA1GHfQpHB0ZT/vQLJVvJVO6vLMfvCct5YFCJ9qBR6+yod8Wotf7g1ljS2rmcMjuaB4VtDmDOm
Dfd6fe8IVdi8HqUZuK1M6ch8ytb0RnloW+eYidlKTaERoh8L2UwwBK1CeAzCvcq1QzgjUXhRc1Af
/vd801RKNNzdEMx4mcPIcp7O/Rm3z6aEvssFOPWaCChv9iDqqr28UPLvEisPxhpe05HjcETV/QHG
5fcTl2SW2AllPi/2Cr3dTb99A43GBf3Ha6tRUk0qSBHFPUHq5d9zfyCQmEBZJlXprpJvOVAiRRzh
KLFsntyH+Ux/xJzXwt06mMCckPcSec/v+XJ4eXCXwjUkiQ5YK+SpP2oHcg54JYpgUpr/5+dIpuE/
Xpa6iH6swTs9kgxo2oHb5p8ubn3A+XPasjMJIbGKy5FUSqOSW/ENp6ZwVNWQzg8tuKO12iyUcNbm
++ZJYIaSsM89PvY+MdmTo4/Mm5cDisBR2Sufk8G78KlMIvtCl/FycJ9C8SqbcNZPwEyPKEJkhyVx
beowgW3itKX/5WOWDTix+pqrH7LixBdgvCtc6TKuIeP+lK5VpAc+xUlIUIIHQyZ+siN87P+sotA0
AnYljLrqZokGnrpx6HRUn8/u6byacEbdiFYloBWVKtSF3meIbVP3dO/UU5+SJqeeztpj7OLoVk6r
9MwFP2xKGFWwJLu7fc7QyCjkgAQH/TfQqG4OcQVIphS+Eac+D4FMw33EtGv+/TSKykAEIrLa2TVr
Z8usnkEr64lj1+OgsHdXuv9iwtwVCe6WxRBETZE2odkhsyqethy+k2kOAgy8yj+Z8ER6BiGdBupY
Nvvyj1Yjz8Yj3XyRN/tDaj6OSQ1fw6tN03yNWO0sryvtDnfl2pGk+E+gkQR6/iDZI1HDtWJHd7Xs
z91nuQVmlrgkCicblx3QIkRmvYbKtyG7VzCGsTfyx7lkKGlX4D60WBRjfeq8mum7D4CmXpzwdX9o
IniiuOJINaC6Icg9O1cgTLm4kdFSJ25vpRZCG/OJb5oQMFgCC7f61uC0HcOnPnJl9b/kAQFz7Dqf
xuPYQvBm2YogiPXzsJCMX24uVx2OSdnerEBwPt72mQZKOuqwp6JUm5yt34uIyKyvAlPtKmIyNeHB
jN97vu1HFhJiemuOsNtSIHIlTn0bYAHoWfPxk/eFxEN2X3KiTn2NWVB7YWRMGvqMtO0BmuYCSzNN
2tu72dgS1bh0QhM+JVgXNXyeeBQ+2r6HxwcbfMbxt7z0yVqgwyA+0zhXghrMrGld7/e7okYHoVVe
gZvPrHT9jusXkRDtYpP8XWHk0XIopLU4h97SlM2inOCzed8Lp/t1ppAQK1ODj6PDtFBS3Eih3+id
Fs0cltKGeuogeruzNL8AgHGloWmy7tyjoGyJ/pf6tY5eOQCposyxppcf6KJgXBU+eV4R98UKrhJs
mE/achyQsGRG7lrAtsjGu4L7LcfSirWOJDFzJc/rU5qLr7BtvLEeWwweDQ95sQVQ4kutAMmxX/qs
Ry4MpcJjn+0b3CVpaT5cbfQvMugOYhOZOIairxP95pRaCNszU2HMEBeKwJll6hsRpL5dNvVwFq6M
YzVZaON42tNtfGtQofuBcza07AL+UWspZMswCiaiA3N/DiFjPVKqgPOKYqBdQr53J3Ls7tizbf6r
PvAib0KfEz7XusL6d2JcS2ouL6XvNcWfDzTucsUVghxp32JCsK/WqG47n8OgtMo1m/+hOKBY3WXm
NGIaYjsowNXd8gMkfmjxfKsmVRfKMX/GV2ZjrisWjBi94Kj7xRk8pLeg2B/SLVKdwANpypP2xmcS
7/NX8k4ia391zNldM3o1PbmuKJFbGJJhzRAxQCm+MC+nm39sHnLQMGyGf+m49ZX+sTRvqzEAwIQ9
eKSVyk2vuQN6g1FN58N72xf75noJ12jVVCSDLoqyflWIw9ayQ0hy+DkAL19FbPExNor430CW+Qtn
E1Quchyndd7Z5QbOTkDZ9xX2MIseU6fJtIy/i+fUkpf8ksd7Hm13/gacJu2qXuolr2cHZ7D/sINn
6NjpKspuf+jPg5Axhvp4+ybesguJP4h9kBFoh1UyhnQBmdgD1lOIl3zxK0VVbR+qM1U02788ZE2G
/ROKOTrATCCToRFhQmbSfAr4V0CMb/AC08q13sLAtSetYcj350BiKjrBsdGfE+1QZUsYRcWoYZdg
Cu00Jf3RhOb/wmGd1JENOyah7SCMbYx3YmbOAfS4S1GyLUCr6wUR2zI2VGRGZBZRWl6xBnSX5DIz
Z7IRiCV1weNKUMkUPIplDfyRBP3UV0sRG/o0iWZDsKYxj7RDmDL/MgaMJCniX7D6IToLO0AVKuge
hgGsGMQGNsYjVY8TIAIR92n4kTHEm3UIFQmsj1AH/RqQWorxYt8PD6M0ncblZuPwZbNEVPfv5feM
SYyGNBGuf6jcIdCn49GSMmYVNs5QnfdSKNXs9D8PnUEuA70s4s/IKJqzo33uRd6Rgd6CQzciuIpT
PJKiDPn93JkSrQB/kr5vrYXAzRRb0R4EB05XxISsqXMiUxOKU6i0Xo9Nea0xWbF+6llCB1j6o3sL
qTVYtJKaim9ao/AOlp2iaDYeueoQCAFeguculQsf9nA6bbqjc2wJzReB1ovDP00m/7R4Kn30+0sW
GEQurbLDbiuCDN2rk2dTmvDHwcu61BMWLsOoS6EcWcukGi/p6C7HVnoCUXttUNDjeACiqHDQv2iQ
IQmKedmwlEZZ8F0D/rm62BW1Yq4DVD38rn5FzEe4weKn2LJnxyq9joVlh9Pf07HR2LtjpLIEMB4s
se8oXNBN9f0t/3s8qfSyomXqyIJMhGNMg0Z162nmezcBXdlESQR2ll+O3kt5vkKXpkWCHi6LzZiC
kkCW69NS5vu3RHT0SHkT1Nw7SLNh5JEgUXgm4fTplph+8C8kJXy68RKPdauEhbb2AYoy/LlJNQE1
DMXTBfdhbxNLNyPc88/26oMPEqSkQB5mPejiMcLbvvZVyXzRlWipSZtOdBgr8U0cMGIXBOKc2s+P
96yBhbxgc9l6gaN6Ifjk5ZD2jhP7PMwkjzet80Rs3WIAjLxQ4UV7154fR+8pPtCszSKVlMyFSLpi
VuPUDgm9PzkV+bHvP6+Is4b9pMNG+u1tamjqqSNP2O/TzLrCrvqx8NWEak43pO2DPLHwDWJiKsc+
MLbwcbw7WyC34D/1xbYQQ7tPsOyj1dTb2TmRI04l5WNWEWjFSdfJKKI/UjGBS7DTJbmZ11KFHB35
9UgR2ksACvYOTvjcWey+Y2HnuoIeVAOfUq6slTpZruiDBxs8rTNhVGwJsMhRxoszoL4rvFXMltYe
vgoOcKQZ/97w4/QyICrE8+3mRlQ6DbF3FmXd+nwp15W3Vd1JPGD2mjqBj/Tax6YdrsNhaE9yE4Ib
01liXMJ15N2bahsNX0pm19Th658kXd19Xww7kvgmfS9VLc+XhQfrM5g43m9CjYDcjA+UQJtoTuZS
17OPV9lQxZm2NbuUnscM0CqgO4FQSnaKRd8AHxNCSZfSi6hgPDsD+PzbAL1yq+ZE5117NI7n4ct4
xqgK4wUFnFB6myLRQjQtnom6YXCrJMKykhspl06XW0+JC5jfS467jdkyaYCHOBziCH5J3VolH7P8
RPX1IvBiEjttqzrnXGM4VOtlTCKYVwu9XAycIgqvpasW9wHhorZmDNkuLD/R1KOVQltB3f1e6POI
ZICq6JezeMw0l1HSB/theboeZ6XwRLMdJEeW5JqiW4j/uxd4LxhXl5MamQgAa1goEyW/YTlRrRg1
toqEfpcTzsx0+ZmOd+Jta1JArEI67VThfzK7t/8i+pzRzscuytVHzs236+LPeR8ojmcSkab4aZMT
TS//rsDSckNxFZqrm/CRO5vwzQhFW0QyMB9mRS6KiwtnHGRdWzfSdWuiKr+EzzEcx9AyzAHFPWuK
JL2ui8AlXaQlKq2lqUSZPC+XPdYTGMm6zRTNZYQ3I6qLQ4RjGJGyVFP2CkDacJDT/wD+aAfW6Ix8
PcknMtsxZt1cjRJXdPtpiVh/Xr4R1WdA5sjr9HQ1vzIjJv1iMtAkuCcolr/qqH4eUdUoKEX0Lsis
NSkAEPduVy7hGKArMNH1SmGsZEZjsKlmafd0i6Mqlm2E4KivKxandhOGTtjf76CaX1uQPneEchU0
LnGLBDvVNnU8RU+VZjwEXbV/FDrl65WmtpJldJHDUTxrmtijoXW+Jdr3P01t56cPZyD2LCkCgWRd
+MMmRdULY1mFITaikbIVKxrb8YZwuGT+4pQzPft3FcPqkTDzQDe50oJVG1lnE/hV+76A8ba7MOi7
wzoBWFwYyNtDaZ1LC59zW/DOEsABSp4qvTMmaORJvzez7uJ4OZ/dPyhnee6PJqRcXq5vB961aSQb
jN/3y1xA7vcb3uNa7DM7yW9nOo9IyoYdcyxUtqzgG6tPlJsFMa8CEfXBpPXrgvK5WaAvSYNZs/YJ
DcEqVXYaz4p9fNcRJCuqFrk87pHoGo/v7Zt9M7y6VcavNbVJzaU+LPOp3ECrIIYSR6t7RqZixhXH
klP0uvYBabtdSIG3TgK9rZgdbMKZSKl2jPd81Jy3YVrd8zw5AGyBHZeMe9KGk37YdcaP35CInp8P
5lNbWTEoeAghJdcWvqeESYrNNa+EknPIirwLsqEfQiYTAeSyxyINRtsw04K7hEAZjd4IArEaI2zH
Ee9Dj+lsEST8y7Wzi+aqJSZbt6cDdzCC+nALK+shs8Iw7tJ6x4CKFh57PEtguY10Z9fQKZeQhHM9
5kxh1QWVDDQ5zUjEdEx852sxVHfzj/N33Y7BGBKt37/xWa99eLzEWhUbPAuIibHMnGt/yXxGkrGb
QeX6kruunLlsG5+Be4h1xmNNrOG5pw+ADaTZV04LNnOsviozrTLQPwV/elnI1lJd8E8WSg0tHdI+
XHGBvFYg3tnDzzoXG0rx85eEfSbkxtV6w8HdKt0b6UQ1UmPe0SFxT7l8ZDtAkSsoNQsw3+9MyvMI
iKZY1wPRhQvQWQdYlXaHAevQ+vKsovwarY/t6kSf+1cDQWsdREw8mClHvVF7lU0UfW6P/8x3FMtr
LJ7tr4JsuVDAEftpTb9mVm2sldWawsqlTFJ16FCucAOe0Ch7l/8oPO6YSwmFqOUy8YHRvQbgIn5H
14b18enhq//ux5Oml5TnTTbtilQa5xv95rlFiWs4wew/ItitEZBg/Is1FYjy9KIs5TCGdZ5BzggL
dLHCopCm1zJP8yUN7D/sP8/IzfAlClUPTuJYOdRQRFoByCYX1e7/EDWC82iG5EhsOxnrx0V0Sc6Q
DwdUZo02Wtw07LkDHLWl0yKpkLBucICsVIVk4AbhwXEEeUSU8ffDhXFFqu11phfx5IWbhCtY5phj
to9tL7QE8dWIXppsXYy98GrVuCpI+ydzQf/o0KZ8rzxfvag0Z1A5ErqnMZpy3xHMJuK64a8De6ZM
xzNHtRhKLHjMcn5ms1GH+RcVJh/iBioBjdQ6a4L9S/Nqc+nqJ6uC6zC8VlO4cw7I+f/F//PWjukB
aM8PNhHk4GVdDqYp5R3h5dG2HoIRHUvrJwB6M8QRBYPJ/Mv7lriDdBcDsq9qXx3crb9SZmHSmXAc
pugCP7vF7KAhjhUJG23e0D6yN7yEhQP2gWYWfv5Tm8njqCyAWj4ExVBd21reDy03SrY/XK6lIzc7
e9bO89UQZ2Js6KokIO+GBbaOHBZHQX5TNCHsKQ1lf2vRMcQApAjvXlT08TXlrMbs70yLeOmYt2Ey
NoBWtxdxZN2czLC0kem7K6df5017GUw9y7lkxKdWIgXAnVavnllhXOFG70CX2UGWrR4wxMWjQUBp
HS5IttyHoSVwCInPqR52Yt0bTTlUBgh8ZrNhGchbWyCCoBg0Mqcc1e9qgjevkuSsHmO7tR44rfNn
Zbfl6aYFFgC7olkEycDfnFADDR3/qwiaCtcEL7b616KnPa94xTmCRRfFKQXVCgLOm94kk1qo1ze/
hcCHiHJWDGtLeGgzZ3dpVV4rWrUlJ+urF8ykpdOOAW7QfYK1OvRvuGaZy2l3DuwxtPNl3QnK7S9p
N6L+BANu1rv6A1x4XtbONOQ5qI8XERy2LG3jPanpWE2k+11vqes8O7D5aFjtLBJpSGvE0hmS1+nW
626N9JEbSYyopgiiDn4IdC0RQqqqPhEfW0NMP6o84reRXxqu3tY+I/OsN8w++O4rtypJRGmMAL7J
5tM55kUIqtFYHcGQn2vMk8sOo5atbpyQIViY303vJiikAzurDl7SCI6BZh0t8RonLIi66TFgQBAl
JUcDXmgNBNFA90krRf4cN2vecTuhr5mXaX/Hk44c/EBs5m+hm/KslivUoVp0+5JfpfWn9CD4d8Wm
8LNJwtTh/UgN+rtNKpByrntFipYGyd6xPRwhy+gcTWyIKLF+0PtQ6dETO8QCU/nz3ftosGeJCnvU
sb1EVPb5+3325HBtetizmzsVm/Cg+VyPaA0pARw324kJfKpHs8r65HouSL8OifnxarwE2X4t5nO+
yWAPKWu7j1lNp0wk+H+aa1xOtNpdwGr/KHbx1XppKu2K8O8tJZlnhcjTjGuq7ag7fute0Zbm/X3K
IXnt8AucrUuiayMSORxh2ZqvNpJoE/N4HOlXtoHCeGWRq4EFl+verlf3VN29i6OQQ1zhTkoMSmqm
R+Bw2Y0dxYVJMw6acC+GA/H8rwPaVUZEHYeaS7zm0GHph6yZ5AhZwHce/0a53xS79jUmdrsNxBzj
jtMfhMziEpMghqroq5QQ3+OaeCiq2g6/0aG478vFmD3i/KzITR1YoLYJFqxxSqK3uwqKnI6Rrrax
RjxRY/oNAFgb/EMhXK7N5YcmOdFki63fHdm6i7t/s4QPlOM44ei3QVeONnuNE5rHCAFDrKodHRX2
Q0/KOUQxkudALF8Z5b1ab3BqkQPuHOXmcPTgzdaSgeVDWEfcPcrRjmsuIA+PKcw/YSw6CejSN4kX
czLtD3wfArcq9pXs7dpEC/9Y0nGrhDdZIJ5mQ+aOCQ9h2r7Z4Asr1Fdm5uFscnEATI8Nk3v40mM6
55H/Bk5Ru3zoBjCQmJH/ihaZlG+hcIwgAywUoHAHmiD0Qd5TMZIChNuDfeAb+k66Ly5m1lysR3s3
z1KNbizl0XVrmHzH/SG1L5B6vHd9TCq5VvmDYIRh214mrVv3CZ9/EMjNrxaB+ZBYmwJjphMxwNUw
xQWvn5CIOu9lc8vKg3x1aZ6JxiJqEYnhPKmQ1oQJsEQXBwNZh4AyqNWoL+nhcm/y1SAUguhVO1rH
4rqJx/AVfPeRH29ScjWRokoNYiPI4wM45M+sXZ6H1ixQzMpI6KwN9nTDJKiET6ebblXRvIsrkW51
S3CKlCHubfuDUH/m9gE/quPZXOEe4i5EUIFw7vubG0lKslGqqRtj4jX/jBrQ9d5B43mzkbHASiDA
/8MMMvAhavRUM584sVXOwEsIuyfGi5DZh1cpn3CJRF3AtccQ2GdqYD5gdbTIfiD4F8WWRkdOSXHo
QVfTeCO4XrdfYDDVx3OguWb3FMhU2+0T2IMvtSKQlKC9kBmtjAgXy9+380MSwaWSFXllfo+CzGfm
yyOI/vYmcvvZpfceDmpW9FnATUg37Z/IuE8FozkNxZdwHyOra6uyF4tFWngJ5DfZtQlLNVjH074Y
uv2g9TWzNkK2yuqlb8xHE+v3VSA3lQ0jb6bgUZGgteFFGRkxCsuEmJ30H/k5NYQWLZlWGbPFIpf9
KieTLFtB5+IYHVFG9nd/Z9PxTr6E61PvbexKSv1l8MvyiLFnlVf/fZxKAderRgbNN2VFv7UJCnkE
sQU0d1M3DSkvWiMuEeHJjaVJxKNaYGy4/8yfbbIszDUnwaU0EyoGuOp7KnvWV9sZhmkbhVQHCIzw
sVGojEZRFpTG5chfo5ImtxyTNdVNHSoLmnjuYPBfyTFjxcO0nFqBUdOcFkOJzbRuFK8MzV1bcLuW
ljxoJkAUX2ki2VCHemQE3nnv5Gft18ed1QUzXXGJbvBY4nv1XqigWS/X25w7Cp7E0Og+qshnt8U1
C9k2jDJjUTpL+fyQw+Rd7TNq5YwLYEi5EIcSENT7HmjsiQELspHVp19smcZrwJgWc28VMH7fTRY4
8irgydIXkxVyoGkPpxuRrzIIwc/9yi7eykUzGHkDm1BHSCZcqIwaJUnWDYSsQG5Ji1AIc+3wTtIF
gUV4g/bmbGw1Prp7KWA1RV/0F9aIgtWjAnTFIgbB3nb3eK5JbdHPGp7MODu9nAHzesY2bnAqn95b
mV0pT2DSb8w78mU2yVoYHOQZkXZPC4SNjStbz1v8zJ06RpVSicI0DGxKhhiQ3yQADYKb0F6gtWeQ
S1kWL/BfT/z3mAdsnETNO0V4MY/DE/4bCyjCXvtXyFUoQdczQd0wgSA3nNsZkYbRCkzqBmEm84up
BR5I6Z8H+Ij/JuW/Yd2mBch7tmtpwhXaxAFuHBaq4Nhkfx6eMWOIk+dI95LXXc/THVg94q5o7Ijs
jBSCPMtFdtscsSliW2hh35stCuav3h8k1g0KuymgmP/Q+Mm6dMf38QSnTSh/XHCpqyJVcspB559B
aInLcEzmTqq3/WmPIN1lYjmPFhE1ABgfWciVHNkFfx5Wa8aPY0xAZ9lG6ih61A162txD5gnCVn/q
BPQ25a96SwmMHMWngp8H3VBObTjy0qPeDp4o9KoTT7Az1uxea9g0MQXOfP8GJkb/3ULgTTCXUNFG
Vpctr228NHf2/IgLqT7QAcXAeHX8ClMfXM+UHAYSqwWV1/xp8qQ+3s1KkLZMFYfc8Wci8PlW+oes
t6LP/kMVYvN9ZDW/xmLsZNHeRdnqH0CWNxoRPsaFCmkhu4NJAEgsMVJkRu05Lig0Gsw6xzorLrPJ
nYWdNgVOxqGVdPZrShZncus1HMIMZQ6N1k1o+/rjxD2t/WcPaVNKRmlOpdF5dEoKYG/6P7TXtrHG
Mnl/epeIOiaRwoGCPCgYQK3wtO0Ese7ovXTNX5oI0vUCAttF5L89ddHix8Fl3weDcahqfNfiU43U
QITo0htw42rA6VoaRtzzDTy8tyldvrJ3dlrM0QNTWY7D8FW725pP7QA5FmsT0cOz6qMif65VtQzZ
hl792pdGu+MRdhYX0MvVfkULEKDC28aSP+5SB3QgqEGG0yzIEnyAZDEIrjJvR6ZuyVJ80m0iobuY
jC2Y1K4jWEweQ5DCQ4rz8lScMjLLc6txSttF6ntDfQgeYmx71tiTHLOYaJx1Zw4YI47z23MnXPcm
zFk+64lyRDkmVuHcb4lw/uYMXrp/IJVahTZfj4dq2jO+HUUXZYc/vilKYsYt5gv7gfX8keANbY9w
K/5nUIUoFkhAhKIW8mjQHE76EDO+1xXvA6uOOS92cJ3NWRDw2srSMI63YJBeeIaYYd8pMrA1kiI9
kkUHZDZdawkwMPh3BIAkPJ2mMrzex9QpR2ZXee2j+8KDVkhGs1YT/ljYDMiUftlydsmeXgfuR9xi
ukChsoLcjt4ISPhXRFpeA1b1SS4biXF3Do7jo3gitVPeTwl0Wh6sY6aQixY5fq7QNiXnWXpIbLh4
EcSquk72lPFmjWa4qa8gZDbq03cgaukmoro4mIaqOp57U+H/3ONm9H1YOvrSdjVfA9fs13USSJ/i
tE+TTde50nlTJ/uclPBZ9VYxpFmrkZ7V3aKm4op9OjJs7CnJuSLyiOsMNNACnJeAAgAeX7FD7Ynl
UvBjZAYTgupWdkm18zB7TQkUbvFFzlTxMVm35JZTN/Ac2/mVctzXHxKh4nXC2ZglvBai4ICqRK77
LTXG0O/g7hASwLO4OklOyyY/EWuXjbJiB38xUcsmPJp2Fp1pqA+WJPPCZTQO+TAfkmu76gTXSZ40
UI3q2Je+tcYfGHTLAVDXDAMMTmy+k1Co+heLcmf5t4Mt2PNempdO/9cpDozYUjv2TPE4u1kMtcc5
0qO6IKkKQT5fsB42BQxFa+xzZEs3nHCLXnNugXEVdytpKna4vg/WbPts94dI6LSmQYAMeWttDuMI
ULoWnZ4Sq/rT1SaGX/BYcAHiu5xQ470HKhmcivTB102OepBDyvhcopbBlBEExtwUGj1WZOC6/BNN
NGuGo1+xKhYq06InHW8OEXzInlLm+yhF8l/mPwgyaaRjUNggjoxIeoypCFWlzBP+mxuQHrhQS6/i
9y/xXrOaQ373weU9WaYFxU52viMRSJqKx8FjKCtjYj05NsDy9M82OmLQllmd5qnhNgEwvAVgJEh7
Ih5TsqmbI0jesqwmtPdJewQNWVLEWemkryocv+XYocIyTh0J+4tZmTcb0PyPPIzArVE9PLeZG1mU
Q/BCSmd+6U7AHM9YVq5NRY6fSs7U6w4xOEPXvPRsMItZOOG9VjKTc9F1DpglN6LJ4HFDDjFdc6ii
9MC4EG5GR3WvgNzk1qAARfdp4R5l9bl8xg1ZezV0iP1EXnvr+aMMwhkftHT7Op0jJCbCSUMsxB+d
l43tqVtWvEyqhbG1bXuU2XWiYA/ge4nZel6T/cI7w4vMFq6Otm42PFNUcrf38Z7vLpJUoAxXjmjK
d/gyLnDXCv3BNEx9QOqAcvZd9ZxfqcpRjyKGwlIQC7u49/GvWk3pa3ayTo/CUVStHHkO2MdyLbkt
4DaJUIoXdZ/JPNN26xVmXu2+xmsflc5oTK651ZT4yuEbMwohK9/X83vowZBK9sepPEFlzHvZpe22
ZoiPU8unGUWRceFWFOerE024hfKcMRtfOESi0YTL5wIOPQNCl1ohfGlDfWnQkvQAiuNNsw7+U3yi
Da7CjSLmyKq0YG5jnUQ8RWkJTMBEJseqgJPn1yxsN3yBSlf03FwUQz1mMelIlqiPotaNs9Ka0QAI
GFCApn225FmXPuc96kzR6bLZ3A/AkHg2mvdOQXzzayxp1N6CU/if4wFTkPUl8i43fNE0SpAzS6tv
MwmAVi9M5fLXUWCENOFMyPiCysS/KyVNIYBNmIHotn6Xxmi1J0IdgTGIr2/ezAX2og2mF0hecHqf
mn0dLnHuX75icVmkT3/L7byqZruAk6z7MgQnVeCi3mFWO3b/eMM9YREqHsqMbHZR0HfSqFAP5aZ+
YIi0hTh4vcpbUEBpugBPDgYvb4SL5FsPnI0rqtN7tNv4iDwgzbTwCLIPjc9ysj68PLdvMxAM64j1
m0w35RwYCJr2JPKrZiRmRix4076S7Dpp73pU9x5getdN1y3as/Yl42wLnMKBIPpZzaxbJCXP0tXw
GoL7n7MDd5Vb38p+Ia2ye2wL2axrQQwcuhz6sb8bYCejklYVBGrDj4EEbigE5eB615w2pbaZLhlA
UhUuErKrGzPp6y39F+HL5F3FJ8PjQTBChHTBQ8Ovm/8ue4+6ZG5H12tkrmw0DUj9wGBh7Rwfk+s1
veOGeK1SG/r9SoeqlWGvtuKspncsFJ/4k9Y2lJvdLlmcR6WiTmJ87Z1o9jBFQQSsan9PnURQo+ck
ctcZfRDMhkmNPcDEoYi5LkfGwjNsuEKxXfehwpjM2adQvUfA4/qpedkCicH/OFAwhZ98VzDGUb7v
oIMynlkscPY7SXiA9635A4gZbIN/QF7mADiOtCjujLjl1U1pP3/ap1ZmJhAREWUuc3QLS/7F+cuU
iqruJX8xbKY/6Vby0d2aDU2NYVh/WuLF8cdKr3N0+gubQL1JPPzlChCjO0K2Dzf/XAPO+5SH1cAL
EgS1C3CPGinSMgWGjS5fI1SEYNcNjFzbCn/fQORW7vpDW35Bn9Spdc4gFsvAmkRumMY8nynrEKKe
3qR/OmFQQvTIBK79ioBhLWVFLQ/KtfwEcfUTbKgCtm8PI3P9tzXtWnxDk/4Nv7r2ES+zuB1ajw6B
jWlNj19p1zVE3l1gTMBQPDk9Yiyl55YsIq7tzkESOBx9GJ61mOcvl44wEW6/3o4HKiGlqamtAzMw
pAPj40YDwqhFmfsMNn1Kamba+6EEFs39wGi1Rqpeijhaw8KvS3RnvZvpV3jY/6+xQx2Dd5MCLSAV
5r1AKc0gJLn1rrnIRbE/GZ0i0K8eDdUDXgAqYsrxF5XLBdEq72SLR+V03i8fB4sG6g3HDGAf2lrH
cKjqTZbI3Iq4aLTcF+28jT1a0sNp6x4OkB+yBzIjjcgLCK1UVmx/CYudvt7XR3Tx5XHMslreF3sN
kOm3tkvNVuVvLUdua+uSwyUcRz2H0DYtRKM3gMRk0NIAwh+5F/gWB+izzo2n8xQrg5aqWUI7SotR
UlUQWSR3jt3Xr4570PVDjt5t6kNAr/4xuOu9X5jkuNaFs+UZ6BEErOPKHgxrUQBDEs8+ICp9M1eq
VunJjtTk9zGD5XgOLBN/f4Thvl2r7vgtAt+2sOsB6oZy8gijNiXunpfiXlUCP/8UxM+V6MkvjV5b
3fhzQaw2+sbZBZMGT4Kc/IahN0iJGSBidF+BYZpvLR+HR6Dws0DraCghKElWyiIXQR4wmvVILjmo
WTm9/+cWzdjNl5nFPU9LIvmXR1Wy7W0OqWSThRGsfVWPDER4fuAe+3xOSqOxExkt/pCVwJ0wZQNL
e3CEigmj6S5O65VIsBcdNqlaCSy17t4HWRr+iKQnVnGhykqtxInIueBF42Vh/4xSA7xkpFt+DcY4
oxzYx/RBG5FUlLpU2lWn2m9zpIylUCqZqA7bJJ6+gIyavwqxDyKMNShD3h3+83BLlO0wlfpqSwoY
Pkih5v242hPnpnUsogBe2QBv+qlqxtzkoe9DkdEgMZPWIhsioFG1yDksLaksiFpp5XbKyeoN2clu
1Pc0lzz5FKr8vWB1MDg32A2AtDVZTgj+tBOm6Bbg94/9S9YoshUR9LHLdjXj6TmaWLL5RMOTYhxP
7SRNsOvOMG1fbt9OUOlEu61tn4/5N56bLhYKin/ADokdpCWjG8+9iD+fKW2T/qVFwdnNaP6nl5e7
xCP+v8wff7776RHRMvo72TO38khRjmIjnO3SvY5ddS2/wLN0ESFLBXDQmMp14Mrcqx/VW1C+LRBX
KuYW47F6A6d8b26AdA8Dq6PGaMgwHGOU6CeQvM/lkGaSEv4YuIfUT7Pnbpe3ticGg72qplzPZYa6
QT2c74+eWVlbFRsQ8r5mPzTjMOeS/gn5fDCWcg70YqgAsdj+oXgr7KccM/RukiU4eYWA7/2IxuIE
XcO7Mtbtvk8JZjbfpvWuVfihMsaMghcnnP5PkJJ1b52eCbu6D8c8Olt62WFBCrZudHene8aMUqt1
+FhSsn58H6LciWdZxfei/ItAJ2AMduu0UEZqnc9+g2/9QYIEYphAz52VGrNUo2b7tsz2TTqIn3Hg
b+gqbtZsMLuLkQttGdScSXoXFPuyMrpEMjl/+oCbbYTM/xcPIXPlHZiGufd/nTy5Z8x8S6fSzzIY
DPJoVxYUGWUdHPq/hjnHFXE2VbpVjUeMydIHWdMycHn9LTUGHQQRQrHoF56hqeiz3oo3mQLIPLRh
jEqu1C3lwM4RSgK9B715iaINlb/JHIJJzaIo3V5R7vTnXuX5FVVr0KLYPFy3h4m3a2piUWcHqiKa
NnipYnvBjctEozrW7oAcWiS9SFKiCVWG97K8FMtDQeShdl3J8n3N8nJzuBh1EnFfHzUIi17m+43p
2+hmeNL09zkSOKzFp9wHZskP4zBu0hhkAI0GeNLHfEciPl+uwICAq5bj5xxfx/ROKq2JAfVbiK4g
wJcW8TIm+N0yxdVxmhyAm7C6nZ6J0H62WIHGhIpG6lo6/Zv35XHT0iQ2l4Zx7UeHE884QV7LhiYz
Q35ZnBSBc7iI/7RuMWBZ38IhTJ5HaWNlCBwdOgcKtNJT49a+7Yw9BNoQ0D1AiDP3MAYfNj/0x/S4
3wKOWjoOVnuOw5NM+xHKRAr2ztB91eiPszqrf6XLLopr5tyaTLuUu6VS5Yg9K0rlvAAP3+wkXwo1
TpyYvqenahfxs7iMWR/VlpFfP2oCJ4kc4w97o+Bi9lFSZVvnGQoZOus4BBrk5hZPs7sByqp78twE
OD23CQ1ujTFK9DJDIs1zECY4pHemG+3qufoCF/aR5Mb4jZojaN8orDnaT7h2N2tIN2A1ZLjGIcCM
8kJo5C/viXdRQIt5yzNEAthqGWjHL6e6A0PV2h/w4qE992FHbh1ues1k3pXDr6NwvCmxHfLUthIu
Ep/CALMalB9UpaSRhuESdug4CiXxLLVh+ooAA1sqdgu6cY3+ZEx4Z5vRvnywER3a+lWVljaJvZcT
wp5ty/H9W++qD9wFgcQ/r4bsndALiy+8LFgxppRtdaQjH/+srr5LdBy3o4TIyUojE8K3bWi0wFmt
chgIeUPbFUS7FFKMtST2cEVja1Y1cLmiOoPdC6qwRkD9/omvOgzHriZModFU+LkTN7aOszQZ4uxo
UYVBmc2uZrjlWtY4/mqvUKnjxS9BeNPq3f1zW4kY1e/3VVtFCTki+xJeBdu1xcabGEtoXuifItdC
YuFdFXmol79cjE1OdrsHA6JX49PiePuhK6ztN18wmU2s+ZxHdsnajDlgBFjih6vXgYLkhHkb5x95
cTTLrsGfqNoMCKg5xrrFAFe2SXYmsgYv2zXCkgGSZ8cS/KX2+ffceAoQZrhReaPULKhPHupsioZy
k53uuC6JzmJx7HCxb9np0ZxJ77FI4PWXulCY9xD7HXdfmqEfV5NaY1Y1G/Z7BW2XmlQDT3oQbv7g
q1/XZ46wiw6ALfZZ7lmhnvqg6UKxgsUIdK7lRxAC0j0o9QvNZRjxN8RA+64wCwAMi2CIX9HF07Xh
hm3B1p++gBI9kljOOUwh5aItEjd+eOSaJZI5eraFScniZQ8vcgoM9XJ7UjSnU0+pPYQsIijsvFZo
aB+VtYwZuEuLniISXUIbH599gfFhkA/e+fM3w3Zl5u4ljG8cmg+92vWNAhIhl++9FAwwcALFCsoX
m3TbNztwsjLOox3lQO7t8mhGs2v/8O5qAoeCiUuH+IfdiuEZ4UC692VtsHFzFdKABBG3viXsPIeC
ic+rj8LfPYPAa5DMr/mSEWWmjQYitkuskOGyJEmzfsXlnCxvI+YgzXBbQ8xEFM/5BdfT/sQg5tKZ
kwazlesufdvY1pEoL7VSAZ135QqGZzOrqibjr5uNnyHpAbkuyOtaZiLQW5hmj35RcrrVHA6gkoyZ
GTVTpxWOgKnNmH6VSU2FC/8n/vSXWhjlJfY603FMTixEujNwN3QjfHC0lpqhFTX22bDgOZNkpVQt
UF00hw02T5Se3VrSK3p6W6m32ycjZh1KW/g+sTkZtY6L4dPmxb5jGewPeDH7pOoAqJVA4pLnXp7M
oE8QIt4rkZsYrlEcnzYgqP8T6ZynCzMUzKQI0ThLbI+Sm3XPFhsPOc0vLvIybLtXvN+EpWfa5H+O
vmlUUgNnlF7mriu+RkPhQmqn/NIgRaeuyJWMNWaP0IS29wDH+HU9CiXPrqolKDaYpC/0n5Mp6S7F
UBUCN2/tMmgVi/cUWHwtHreAc7q2l96BEuvRAGXwdPUUUwsjm+eeMAhd/fhRCilK4xbQpktOrw6m
KZM1BRaRVjtelM8CY2YUdCvXxgnYKQV2rtSnpvdZdTWqDbrn1M0MeBCZDN33fN7feij44lQv8yCO
QqlEbgs+6enPqrQIBP1uJ32qOKV87XKbD/9jyp5jOysHY+3oTuYeWjNWukJX8chR5Pets2tFR/VR
U3RgETfw4RcC5FvPTimZfD6708X316drYa8SCkL4GI656+PkGSpJ8/phqbEHqDlskxzRtLg+hu2W
uVEVpt/sWd/VimuZL8X8iswAYX45+bauwxToZU7qGsxpJpR8aNMemeiyqoJ+zv1UYYQ2OBrFbPk/
URcJWgNxg8wm15dLSM8RDSOIpBpXxAZmTgZwzksIFqT87mry50kbqwB7zbvAQCY6pMccGqlqAkxn
GnO/QOylXRSHi2jRMT/P7GVxqNHEMmIGsmbdHc4UxzmGdVrcrV5IQK2JVeer6W/2xWO4BX+uX4RA
KExd7Gqov1l5V0NGnl0wFjqz8PEAZ4hEpk0xHfca3Edg+W1i2i98FrMkp03PKDHqb3jig+KqDOYe
XNc3RJmk9e2iex25ckS/nEM2CefjLJhXwdhfh/mnt2fMNrje4RN+Pxi4UhgA2wsF/BwK08+1jbax
Sdawmg95SqKOBiqBjEvHnrhURFQgZuhZgIAQn4VPXVDjfBFrCzW5ZlC4R0L6ZCUgsaNPfv2cFfQN
pP3+A7G42utbGxbL9QnR9q/k+WObHi0EVKMSMM5isnEFkzI7pAW6Wth44XidJY+G2oRZRCvQKHqU
3dSi1K0PLeuF0lHhHdRiM4rOCT0EKq+vjKmKvQHzgxs+eBQWC7F1z7XORvrZ5JOrkDZ33PXpPedF
Ja1iYr6cf7hCFCfsLZVs4FzHxYH2yHaWKefSbpicSxuGoZD08e10suixvfWJmCkbOzCVzJJpDJFA
m2E7S+QBHB4BkngUyP/9VjYJEsk7FUrDNtxr+JEqfWq25vDDspbLrgEvsgHNKcz+gg6trmrb/iTH
w7dfKr0p63zo80tCMQUUK/v0k6SsZ2BHrJQhl6dt/D/Ol641rsxTHQrWXYVn17vkI9bt6EeEU6Bb
6GxLgpMonzI/6Z3x8yjpogwvbMeilmBIBSMttxmaynYq3TQhzEunseBA1glqZru8XhpoC9yr1KSF
F0vT7Z9XSbVgT6scn9dISWBqk09EIGPu9Dad4DWWUqd9yfWZxBVsAii01Wb1biVWwWyqTOPOkGLa
ls3TUNhuMHD1Xd7IPnyAWGV+d/+CFbViE74xWwuDiwSDjsKgbS6jiE4nLRHSeL0P4c1BkppcnJLD
plXRMRvO/F229Hqfa9M+A/YFPCfN00C8RvCcWIegOpB1M1v9qjvloe5XhQkWTl01hYCcv4DA/9H6
MlVcjebvZQlLTYw5u8YEzT3rHWEmcC+pIynm/Jlksl0EGKL2luvCyd/tyxsbsu7clW5hcQeOsvYt
HMrDkME0SpZNAi1X9sm9aZZxCbdY0nbE38TiGaIw4CorFLySNzZcOs4+0LdbKSA3HkEW5KYLMaAS
+37w5balCnPUiEOY8UlbQDRxG/OZ2BZelT7pZA7bh92rboAXyccVz6OUEgqiECX1IAhnvNyiDYax
Z/Ot0AfhW2zZ1W3kC9SJvH+zFBphFSF1ciu+wipAr+SItpP3aBEfzAWnGc2yxq7Pkd39CWkdjMai
duBqLh15Jn43vUywONQG0zc13me651DHwZoO3AyFyZHrj7hDM06HUBCwY49z28bhZopK1qN1KrIF
Ola3Wqan5ARm4Lfg7mGPlKq24IF+hI6TA+tHFBGD7DKCz9ZIHKL8e46xDKbaB/ymA8iF//ljyNIh
XzOjPPWx84lKOm13KNZA1ofmtd7t9xwM11CouomETix/zHMCAHKwxZLhY/AugNux7wEk6Yf0SjeR
LqULBDKu9Hz0OOFg1TzvQsyWEAv8SSHuiSPuZumN4s2GYRYkt8686t/YhiOlGopicYluuSfrV5ly
IL5nPxbTgX2ONfIrsVsmSo00tKBvszFkI6Xzz86NIX8mPa7cn55VbcaAQVhuFjyfmAekMu9srzMr
m9i9jwsE5F0WXq2n570lPTUGkE/RHsVIL9dDI+n0sgNYaXrTuG4HbwXrgvI5IXfhMeZHTyE7m2U3
pGBTYS4Ot8dS0cFaDUWO1WaD9TBVGMsKB6w5TNfxJaszNtA3K3uUK5F9MjUr6lcsbCk7ZXG+GMIL
XIZBqQL1nhGlZYmNhmF4FkA7HObmJJVING2VChgWvyP1Jif+3pWheu/lOj0TMaedSaM4t6/VVPq7
NVrHjaJaVI3GErpPCsvCTbBE3yM4wVrO7PyceoPttBDeLoLzeoQsKend9QhiDxnx7YQ+1MtdL+2z
c0YyTm5RnLJEsb00tImKZlHN7Wq+8vn1fpT0lCYLplFSV6QYAXzU/OnFDc9TSQLcODK5inaVhPaj
0rroxlULcvr4VNMbX9LJl2put2o0qHKFWv121cvmdoP7a7hpd8UYBvBfuTI+PQnIMclvaCh9dJeO
Q8724YSaYBCShGwmCxXg/LGsSEXHEszLMY0Gs8gJ64FFydUS22G+s8YkNNe0pzrL0CULolSwbC7w
u1dtaV9n5F0OYW6RdnCQAgN//q1yd3jjOAe+RcnT8NNjk7Kd8jAZH/8e2sh376Z/9mlcKkwsMEOH
6USk2MWE5bkzM85qv399sQR25QJCltYV7jWNjFUEIwuHH1P+2FS5B9JUjxoKD+1S1p1MCdKG6H/a
FoGDyazejXEpXfz0/36G9m9BwrkhE1Itmz1ck6Mce0hoET+rmRsR0f8zu6JsMeyqF6KSWE8wiPWt
HfYv8QguMoUBiAC2ca21WewR83SE40BDaVlkBKEaAwHZffKD0UJQIVQc1sqmyWZg7Ry33TVzwmVU
7heULQi3Daw2UPEeD+PC3ut+vJd2LxKthku3XQRVWpk0nk7EykHZ1TIbplCHhI/XgNkokFMGlSjj
cm7EFXu0EnE8+nRKrc++I51xMjQGbGDXiNCynukpGM8taLvhNptDEYUZJvv2u4R/mXakno2iT7rW
pBlfmFn7ioZBFLWe3gSV2+9ca7TblufgPyTKsXOwhSX9kaTFZFAM8YP1kN94gSWYGBBa2II1I9jv
UBaun2FKGdiEobLT/ZRf0NDZwyyVTS6ql8YNEOKOebmChREvfbGDt80PsjeS1wJLiluD8BR20DR7
sCjjMSEKOk6TOEz4j3J2rpcXf4fnqBSLc1EtxJkOjzDdT2n9Bi7etlA4EKp9Uz6Qhiu6OgHsZ5Tg
N6ERA7xlJHCaml21zAY9RuPXDui8OAoMqZSG9OZP0vsqZ2WJ4JezdO26kt6l8XCrqN94lvsgnjTW
+CxsiIjp3VoJ6fP/ghdk4bSn6JFevP/vfTjxDIGabPmRGzfzq0bKRao+BkgfkR5caHgRlJji0ft3
i39wu01nohBhggtKbT9JTnT6PI0v6YpTcovhh9a/t0aF26oCi8CZfI8spdgUA+BbqjbNNzuRrCwN
opbUxvevkUnBDISrDaOL4KiXGdyBYABapnXdPpqlK0aIy+r0ZrBoHeQg2UYY3YT6f5yVHtLIuep8
B4sACmY8zo1Xfq7XrU/viMPlov0/ndQAoMjd9qAURGiJtshpdeoZH5vghWeXby//EACJegW8tMHY
xoZKuCrxvyymoaPIxHgP8utoXNfqtMZ9g/nuEWV6BR9RI9Yk5BRHjsw7zfuQy/o3036ORjy5/okE
UKyK+NORLHPwS3tZ4jEyCXMNuQY4OscnB7taxXVBsaXP6WXlKRhbGKPJ8IHqindG46ynw6oQYx41
nunITl0mUov4EqbByDGxvK1NUbohL5KHRZ5EYxp5j2hpAUllZzVdVOL5ZCH+2x3JziBrcnMK6YRX
5RdO2eK+lpI7+Y6LLs18DSNSJcHfGp9a94hmGHBNjLp8yyxbPF8eE/P8J/58cHXQU84udjBD/yA1
zqQ7q9co9DWYmsPttVO2ssacVpKihd7M+Z/hOzPgXAzugnCrKDi1Hq8MkBY5K4bCTNDb206514Uj
jcW58+uJoaY+bCm7hPL57bmDM99Fj1GxEWAlRPmAcUxeq1oj6VR687Z+cVR5oEqV0aqjqmYaOPOi
o07wmkn3N9xRBibfR5Zom4MMGzU4mD32WMmfjkHNz1ypzEbj0KzR1mdMh8Pb8Y9TrM7crNl35lHd
Wa3qcVqHbeXlTW/mDBMRpUA71v8CNRjNxkhSRAR0EHD9Gb+gZ6oJSuEV6FbFLba8NcirWoWuI62J
CAmQQkVYRpiFrDFm/HCeyYmlle5MfPajHv/ZSR+2SgQ4SpBGnaZjXQPsyD1iBZ2bKVD7TmJIbZHO
8Qh/ZQl/g//167tYsCJmtyjiJ5oKPXYh1y5kYTpBTceEzbvn2NdIpdNDoheXyHf4wc7rbkEQa+uA
CJo23woMDtILL4xA78pE4bRZRiLeERwHVMG0wdBx7oEZS0okEOBy8VEEkUK9S1K2hRLibNUTRuZX
CHe+2eNi0+FNdAQonRFb7TvaLB22TitO9gimoCc9R7UOyBjKLAZ00slOHwjs7goEXi5YQtpsHzZw
LBvoRLO5s/PJzeHlJlD+YG5141RYqvTCbesZmSg0mV3Akekx9fMZ18+Z92+GWyXij0nxOYFqn5Qs
mgUToSxAuvp7WJ9GkIpsatXQX5zt0vP8pSgdFEwgJafodngUeO0HGn3ESwOEd9WvODbt0k/TEgNa
2LTd+SCywuUwFM5h+aIPq/ovDQF0m5cFqs94et8xSuhqW7yC0dO9Ba25Ay/sJaHCD0mE2yoNSLAJ
dMPlvRVNp2CBnThARZmHZhLO/dWNx+CQCrJDrUFyoCjhMIdSc5SD0os6yDeOpPuoUuvcHgURaUns
KiJ1WjUZOnt8uv5Ho3V/SqlzKQNLainaZO9ST0pKSlZxDTn+0LhddMBddkwI/idWLepLGNAP/sJJ
zzQoh3oQVpC2+DTHncjILsUIh2FsGMhyin+gYzJwSSJpNdZodkOF9dsLdYIQdzAnYM+GVBZjxu50
oYu0/zqWSWiXKGPmRRDsPC/E4xRNh6tUSQQrjLCDkLsivLvTvl6HlnYlG/TO+bngaoMDsmoMdmpT
60vZYjseYZAOA7BrpiArKpvS+0WlzMXcRNFgwBR/BIR2VGHZTqN4or0Uk+zD746Qt06Yjh2LFVeS
KW/LHn5mBu4dse3Yvd/ow0JOMF282ezt/FNCGrpVnRz2xT+THMWLpkwawKGonj4jneIPHKJklfeu
B1r8Ud4HYSBh3KJPMDn8kJs1683X1ZtCZwnZzZiSU3c4lMKG1qmjQwjKNLRWbic/VNC2pi38hzBg
r3ZLVDq+/FABavXGj8JslFIQ3QjYfivs9SH8om+L4v6F+obZ4BeFzTFk4D13ic70ZwD6cvOC5duz
QARMW7R9C1drAI8DG6BQCgyFZmzy+zomVqxK796SJaqqVzwReKwYSIbVWU9a+GbFeFOauHGqTKuH
sLZh6SKRf7LHdLKMlMQbcNzxQit0AGN4rJdFyQ751cb+bXAXxSfuKSJ96Q+2ZMTyBP1h/JZTw1x2
IphNpXOBWpK9uSabTlVim3JZhzlPBV2CVO1L9wgckWQ78NzB9mrwMcHsODyhH0Tbedf83KegDlEc
xiUhaRltIv+YHTJj4M4Etup+L9IYFavCsdG1EAbyAPb4G+bihwzDFnLFEOYvkjhScMSVaPV0R0Sb
q6qsD9cu6Pdd+2Gjx5AN/x+9bPlRhvk9A9ffoWOWwJ4LF6eLH7WIVY8nzQGHr0Ke17+avzOom5hg
19+5/x26m0zsoCx/EpzxlmuHqi2s9rTSvnkF+Xq/YFzEpK6y4+JP8qgw6Gx8cksmZY+dk6zGuFuu
h3fG1Kr/dg+Wjspj2jmteRt0TFccHeMhIFJ8D2WQEH3vW7nYKlJHZV450sIX3IKRs+0cA/yuReVs
RyihByS5ZKR7Wd1uvms4agkiKM/Lk0qkLOxAPQSsCJrgPqD/SLq9CWi94FFIO2nj3W0QMA7dCnTo
3K6SX3nmvOAMTPccdzf5Yy+ALConT7r+wcqOxg793sO/JVHhnU6G1/K9qBE3ymXxJO42ypat9+/R
wroye1abdI+aSRk7z88oQsEiMa6JOyuXwhsh94crf4SAZx54796VcB6jGT5hy+6yn+adglYVrYH2
kRQFNJSQCAfpS7edU2unBXTl9hXTa+YqEidIZi0J9Jfi6fZnkpVA4zZD/6skpdH4XJGsNo6vS5B5
TNY/cN5E5DrwxVMqEp9TNDDWwbofi5LPd+GlUfXCM9F3UIegxVLf+BFT/cYaH9+6m/RujEKgB3UK
GeQDMx2qCPEVSxwL6AfoUPE1WXxuEb1dftH+UeD+ZAoR34L0BFFXJGix/DsRgbOL2IE27XrBp9hP
FtSMtkf7XmdqGJIvCp1PDcVsW5FsWiiabLXuZ7zo4WK+aEGO4PXAGR/PSKURRA3CHREuCf5AEJON
eQ0vWdsf2u2aZ8P11Wk7CWDTk66Ekx2ZxwUEcVh/NMAkTb1B3TKaR7TpQ6EBfGDSrO8gm7FFcxHG
9YYSPZJAglZQXKUsH8ETN5aFsRBVV/OJic8WA2RYvVX+Gt29VQRSFxDCdwOht/dqWZvLbnQHCX9a
KP24RbMOUX+Gk7dtT4xzROyQ2qakGG8NcmOVzmJpMShXrnDuvJ0nnEG9X3akEnK+WRntVw2f+P77
w5xkdiEeKcL/+L56Xo3m8bfIP0u+xhCAunUN0LVAtyOjX99I9yFK1C6KdrkPsmCPJtDfOPIgmys4
VjrX428GNsjn2vEQag7GhYpzqGfXl5RlMVXtGsvqAdIo412oX1lJV7qaTeF8+dqDvh5cvw8dr20r
Ddn7bY8olp6DiQ72p3czXauEl6d4ozJqBoilqZgXU7JfuUSOKGZetqLhxHTmLs8F3iIbmh0w62fd
OeCPYqvep26XDo/D/5XhBZboF4VIqD9SJvLvRe9OR08gIoN6lkyMcoHezu6y2EBIyvPdHJvDg61h
Z0crl/4QXAHmw8PrIcwUMoyh6rfATRYycI2xC6bmnVirBUjyDGBOZ9HE2emPCWzzfMKiwj5lZEQ4
2XxHoaylxFkHJPuw64tEfHEtXJTXmyPSubWDjOjmQ7eA2J3mSZPrRW3QB7lvvxX/OxbfwaHazuoZ
nv77Gq9B5t1HVrWt4zY/FG3TOUgrYcQfGjLTe/AAB3ZXTf1jKq3q+Qz7/PnsGz+kK11f4wrOvi6J
q/F9W/vBfl0FmiW/SEZ64JzWrA0ClOXvZhqPMG4J5/+pJP8fAlbClqhVifVrioSowzNCdM8uVyVT
4OUywM1MSGOgkNjPkKF3j9r3w/W1rO2ekXVTBuIQuLUUymEa2EJ3pdvkxsKrVOrfL6UnyCbOVaaD
mbNT7Q2SMk+N3Te7NbIZzT3qU06/GLsQ1gwWtHC+EC0lHGwVT/NpMogSHW5CjhpTe0Wru2Samfgu
ZANU1KtBXd12zZ08aLzmz6SNk4UYozB344oDXZnGkqcG0bK1a9ZqQpWpU5nP5GdEW3yj8GZJ+1IR
ngtaNLKg2DUrWuDnOymy+TxZOAE31gTCFfLWU+7YZ8ZtujfOCrXUy0du/VzcbLWeEXPRZQ3DRp4/
AuColyxxBQytBlgHKAYoQZld8t0uVZvNoeDR5fwPPriOk+C726pVTYLqC3oYf8lEa7MKoN+IInt8
w2Ttm14H0q4wEC1j4gQb3DjunzAtZmCol8ogD9VlfpiT7Ql1/rIZ7sZ8ByU67PAqFut4qJGAhTAl
5514NyfNcNUaI3R5SY9kOiyA/CELdRTPTEMBDnLL1PXfDWA9I2kEVbWlGPQLoQhi/9sT2xVcxJ4G
AZk6CJgO9VE7xkAqVV2/6FQMIgRi/Q3JgBqveeTNcnml7Imms4bpVS91xrIaM3KGZkDSpqNcrvnn
tfw2PnEsXPAXcD8NoBfnywNFkEvWuAfDX7tgjI1yNPvrbOgKN5v34Kw5d9rVOxyswNZuI6lUUzsj
uDM2LF4UUruS+ZSUMAeb+s/66HP2t4Ae3nhFMs+bQaYRhp91ICKpELom6QFDLHl2yH2wJBhP9Z6W
R/AhhMsy9f+4SVHyLOztR7eDSLz80fHNaFasweKyXaZsbK6yXvyxm8o3wcW8Ms3EyIeCfoXveRl9
+At0XdHE6IXLL+7aeNQSzyJ4BTS7LjRyxLllyWR4Tdh1NvAAEMZpvulrYGhKItC84ZX/Ehjw2R6z
6OzzwhlJ/MHuIUnKTl28jHba59oU0bb1KAXBG7UJR7RtGAeJg2rCWo0hcrid2ECRfug/f2gvLXaY
hj3JZJzmLcjolM5raMtetAX+6tAP/aMMhvZC4z8/4IxFG5Ib456nm67zm7a1EQeeYIhEV3lgmpgg
vERACy21uPBLPwxVNQoDCDAb1U08QWT1MUZXLjQ9Lw3AbaQjHohiy/0sObLGFtWShIZ6pl2Cvh1J
FByZPl7x/KtqA0Aj1jyktG8FBTin/YOe4eiYoNQT56LQv899NTcy5Cwk0USIQvKAhdnO8wEzudl9
GP4aIM8iur6cGJ4DFk7mjzwOyLjWSY32vu+GAbhz1eKI9vTlBDS0PHwmTVtxyOenFqDDQ9sSNP+f
zCeWsM+q3pRd9zFpdaXorUIAEZ4gI9bb8gedEJdatVTbB3ibN8YXk1qFlReFI6cu4jmN0UU1dBBH
924FVKaPg1xrnBZaN9KeG0Mj41PY4VaQmMUH2I8s+U1mDjYHUAFZQVIhVggJ7OQFfCg1pLwGVp0U
Faq1jX8casVFi9faf4SOaF6FFWuHHylAJTg8sW8UkxPSj9sgDOhVkrK65iQXgYFHrw9NwWUSnwPv
k9bx9GlbgR0BCZmR7NAPRZyvoptTZcHsoz32PU9gJsoY0odcWppulJsT+YEXTxAnBkOBnIPQPbJu
kJNt1y+NsnN3z/yYHprfgcQQTI0Jq5iCcjS31Z8zOukIYLMefYCzu1qVQo3IfjbrjK6WZXvZZ1X4
mjkvYMQWV2P9zGaYZLvqWx+WRkSYR6ZoJb4mkc+OxCneab/9O2H4nZsS+Wopeyes7kbCQKW/XG7L
29rsu1biA9K3Kass0OqOlvrUOyB5+BUwnD/MyGU6zbq2BUWpAAZVb0ESDQRmKb0tA6Ok/uojN/vz
XnKTSMg7nYe/drcEl+JdsLN9IzwFg/7kPbTFqQoDj+NvNvWec2IvXIjrzkQ7HfKj0ddaCOUIl4Ir
koiSWfpVMHFJ8MGu4Z9pgVNxNAY/AwV/Sa3QSRZI1fDUUXRUbq8moXwq/l171wkbhzTLtgTED4LW
uSMKKlLKbUSpRP5Ol0P14SyUpEE2HYT9X4OTtGQ5wR3tHGyBn/R+9LB+8GkhPqgaI1iFgOGVZECQ
cyqffwmSeKzG0xT5/oBcsPIXkGPmIqUPMk26FanbhJrO23Fs5vziDKPdUOfsZuX1etlfzZhpew/8
ReYajLV86Bwkhv8ZCE1y8V6S8XCGrGXEUCRo0cJgW/KY/riMfKbHixVw8zQ2UF932yghH9LuNqyJ
KxUICT3T7ykNSnVIRgNrz/nuf8EcmQfe8NZwteZI65w3V0DjDSd0ClHPI0SCWFWjnKWp61fZ26vb
t+zUloK69mKnrNDNft9zW0aWdhhvYm3L3eg6N6ms2mgeLztVENbCGeXqD23qW5KFNxCMzso9KOla
iegFY3Br206IWSCM737lahyWPb1HbFGZ6OpmWFJQkNMFQ2TP1Xx9iNxeiQNtsSShRPFO6Q0mxx6B
W3XXecG44pL1vLhjmTYfClhtsj1LDmn3nCG3dO0nRyugYpVVk4LKuhrrHSIOlm0Vam0Dv6fKP03s
LaLTA5QNRHMW41KtnbbYYKeoIVBPXhiI6p+BC/BTBM5p06UqDIDQtTGjbFfnidfXxlqZKwpKXceI
gnKNis7VjjKtbH/eWro+aRlBe8RXyuPRhPkHSJeGU7WuEY15l5xt4hDqCA00SlE3LIhtGh9Q6rd9
KGP6oFgoU21q6vrRMt8hcUygA+o4TFQ3aTOmAZI0FmH3VD3TU/Cw4jHvKLL400h2ilz/+y2exFTm
ZJ1gg5p93SgZzJ0whYdYH8VAe6soq+e5wZ11HcgEjIpdjPiZcU7CXbJ2LJUSz0PH5kCdzYP468WD
oABW/XPL87Bx4ATxJQ499n79wzvZCvKkrqiARY3MpxkrspSdWU3vbI0GMIN3V3gISWSNE0h3hMrR
IsgZlio2ELglyhocUjT3Xl/tPhF+NP90wdO4UbK9CIWiJfNv+r68ckjm7SRfsaAmQqlBqp95tkyt
42++AGw7ohAvpLxFHTo01N1evj+7IIMhX+2jTS5Ovp8Ogewml4JwnQW8aorkou8CQNBD/5Coz/cR
MZ7hRj/3MSd/V8R3qGsaHGwS3cn1+RtP4iodSu5NIGjDeVjHKVftUKrQPG6eUQ1J3qu4PmUjIfrH
XrT3R/lj42TqQdGx83vC99YDYsUhxWLI5hG6ykHCkWuBsHGD40BgvHbFjsTkxP5W4M6GBrD3g1t8
3JxmIe5H4CXavcvtoQtdX5vFE/xRlHKp7+Ks3XBlk0w2z1/OAU66I5pK0uPnd9nK3yxSJaSZLUlA
SEGPDusa+3nQuGD+j78lPJwtxNP2WMDaN/70PICyzqjQF1FnoAicm+GbCs1D4qk8vOAMpcgcdhAA
tEwjXbbrH/VLXNgteAnSHX63GT7gZe8mL2i8a71Vn7+tkaEd1j+UOPGyTAW7RfI+9nVZkeYA8M1G
pSGU0yH3REVXK9G7BzzRg+/Sn7mN1k3n3o4IdHlnzCUyFmil1tEV453391Z/rICuaign+7T6/1zy
Qar3kgCwK4cES922YobP1b2RwIdtg412agzq0JxT373EjEXC4Ki3PPxaS51fJUv5HK9RcZWAraDZ
4efaUPOYM/YvbCfel84KDMHQmzje5W6+QKmi+VSriTOsDVs8kUHQkHl5JRxZ+3HHdBGmRDdSSXru
Ghd8e+Mmz01pd/7B7cbkS9T+pqR2J2yBvT12ycNRzp8eZfXQ+Z4x8GwtDZB7/R2kbvZObXZ5qePs
xTrYa0lqAdDE8mfn65mZx8t3fyIZsqZ+I72cIRaNF73NqatkEH6kHpvGioSJ8rplNHe2eS3Fg+HA
F4Imx5twTOWAu2ei/AvD0J4zfqCHho/eB6PybxQUryxDWV+EiLDAbsKJojjgoLy+G5SJSl0kLB3b
CyI0MdNgcBLzOQm/W8Cb1jkngofGXLh+oxJWUGjdWKRZWE6sHk7RfMD4OiqrnzsrwVDGt+QZCWmT
KO014KrborJTuW4tbWk15G8ZjfEtvz3wljq3Kt/qcc3f1nSGerFXiEF32y5bbNwSPKpCesU4wE86
bfgbQZE1myMqhy9O2D7eAH6HP3X4hbO5UBvXZL0aGi6zM3cMkB90wU5Y2BJZ+Lr27wuriWk6rj/A
lGuIDXIfw0NDo3qLQexd0Ybmpp2Bz5QK01KEPmblQXbr+GhANGAOe6EukPu0cip4BTXL7m5djmjY
eX2j1CwYakEripFHJYatxFZ7g2ifZJv/XjmSMCshWMEVMP5T61uxJQ9EY4ldNeiodlxuSu3B3apc
4bMvy85BhRQm2yJA/7Aa+Bk6NGscBaU+FD07W/WnLgwWsBdbym/1+C8mhtoGSJNzZJ9rrkOA9jxd
t0Pz0Dt/JUS040008e/sQcXimAHsScIpQe8m5u5vz26ieMSoQ1L2Lkt5doOFKZglIOJThAyRCV3F
dvpixTqCFsoPDXsHOLdlECPK/F/Tcy2pkucjiyoHY3NIxllCHUD1gbnLxiUl20i9MD6LX8XHqap/
Bvg/fA8vCpB97bRmH1jIqj5g4nlSrHlJQaRLxkfq/ve0hFOyo6Iag3Zj/Js+OtojpK/r31fAmDyg
g33ORFlM8ynuKfQgXjjbVRfUmn4VCUdo4fpAKPlrz3T3XFcpwed5wPSeKfh/ybXqMCKvR+tiV5Gh
A6w7jo2zHEQIw1YHfI1WEK7FgH5ZUbEVAjrul6x0OQdVPB0Hm8GrImwJF+xLY3ENEuClOc86CKPr
j+ys4tm9uSz1IxhBSqhQNVKk5x+XLP5oV6z1DPtBRa9wdL1g6SYA5Dau4KfJHduC/SnPwfbLV2qn
rhTZLjx320BEhjWFc0vNcqCREIv2Yas3o4nwY4+859CANQvoeyoKbWFY9ZenWQP+P8i6y4YhbUhV
2AQP6Ol04smsVbAXXRKD2WhrY0iV0VKlp1xNAE2v/6u7HxW+8MAN7dQEFZOwBevyZS8rmezM69aA
2DDlbKSbX1Jh8Ft8bB2fTz7gqYp5jskOENb00hMnNcDpuKoxm5UC9T/XwKFYKx4lncBkNmTERDkL
//R4LRwoygfGD/iVPptW1DPaPSL2JoHO+txyYwuUR0EVg8i4vy+/yMMEblas3LvwY/unXsiLUc3l
uzD82xQqJCEbhCpTeItD2OGdKej/9ANhld/9Z3tcRlCq3GOTA5EzqqNPq2/8+IdMmp+DRQSd6A3k
FNsAOtAsxPeNfJJTZK/bEyIVffej+a/0oBaku60Mh4MyPMjmj6nmS+RO5mfjCg0UKuWOnzP5bFZj
etbmWxLbbFxCmHVPOe+OVVTuDluANrTgLqUd5dHdfnJzpOSpo0l8aD9wVgb3ICivjEGvuNG7fpnj
fgvsesu3WyN3eN4wDH3Vs7+HNGH2w9/byKH0+Kk4mLMy2F5Ppu4axMavZHXcXVtgb8GaqRiiZlkj
hS1JcjiwcVJBvNa5f9j6F7oKlkXHt1A4egjNki3e4HKaYasVRkb+jBcHQw9aHQ7Ug1GMkr06W3NT
JkgOGY4qFEYyiNOp4XMOstgxb8HI+K1qv9csqgGc8mdbDEv0XqXSBeKopWxWzpn7Vpgh03sfgXyt
xs+rNS1BuvFv6y7loaNGbks/8DyEhAmsiFPfaDkwTwHjbReJzNWvCrCaY4zPwD3+uV3YNnPcgiCl
19Uwrv/4qEB3+12bWC5MLlIy4n80iebIhx4iGOdT2MvxqiID5vmbgsTkXztAn/tDDIbtZZSoUHpg
sEoxFrWMv3+F+rC9hd/euamvCxXqRrrk2myR3upo6252F9C1cVToV5qEJHdkibwGU2mnp4rod33u
20uVL4DrcvanxlrECSIEXV88hQk3faPZFKojphuP536Ze8TB7DdNMFBVJ6hL485swJ1oGpddZGx2
dvCSpOSzFUsPXUYOqopjAR+aT4HR23aUezJIXph2WJGrmH7CAS7xcbclmMEtbNZibdOHB1FPMGnx
KelE8uFHUPXcpf4abD601QA50XfMzM21ieb9x05Tydd365Uc3fuz32sjzVMcUynTddq+vunOf1fx
RoDv3PifG4TMg0T8kMchQduInFRJJH+/b1HeKU38UWUYRpflwfY1wuDeI7Rp9LHKIFi1pp9PAYtY
BgL08I/iTrkLYqwH6/8rBkR3PwIC+LRJ7uBnElP9jgXiLoNGWR9fyyMCL1OYeqNkj9raZN3U3ygy
cyRa3mBDD/4HEDZQcMAYy4zFB8MlHaR6YdRbIM8/rUu3Ujxhjget3Gg00GxFZfVdwXIw8VbfCNbA
mzt5lc8ewP3XPvypXY2BtAH9pXs6h2NhhFK8fzpJ6UdeUyZQjspCIiUGOVoQ5+gM6U7LbwNVyZpg
zGh60v8Li0UFl6aUYAoHaZFleRLt+6WvusqRATfklL7+66e4swg9kpARHjxMXoswoh8hcl0Ka1Ty
ksIq/MIHhP0QUJHH7BsM4k1W2SaiYlR/RT25hVFgJslUbbG24KTUbVZzgYqQpvRa1qdW5nRE4qe+
lQvWY0xITo9YxgBYzfVtyb/76vKbmGfW2DKLCXOU2zHmEuKSekr1/x+LRm0IQ5AUpSbyTF8XiDdB
oaTIAL0oAtfVWr7G/H1Nr4CEpslb7W+SHg7QdYLzMZbS33iEAiXySiKTvMV1ZfLRFgxQeaWI7v6D
TJ2Gw8PgNgir8pm8DB+qRhfUDaot8V30+gHB8cKv8NszhTyql23HBnQYhEPFtjfEExevTxwaq374
G3rBd35ihCy9WL3ipk3XLxRB/nd70/LAnQRzWIHqZU0f0/hj5aoWGu75c4dsdjmKxPfGImoLC8h8
IZ8VdrnmUeyV7pL0NLJ0sO8vXawNRb3ayJ58G3f60WBHw1xM3AS9wJueY8I1Y6DcVHPcg9XlLHwY
synh9akihxeMDWFKILjDX0cmt6w43DP89esm3wVoh3e/tCg+7Kq+ehKbV8DjdRO2m97jZb9ZE57m
8GW0wwNcmJ3R0ifOzXpvhcDUACxf3SFlWB+69+4ZFu6vFDjkn9WeGCDel1NebpejUwmpLrpPFaBa
N+xaEvqVlUBSOVuEH/B8fQGXsVHovtkBXvNPM/CYAORD6gHTDYdXdtyP6Ge8eBgYXQ2HIKfCHVpY
q7IK25HC8zp084Z+M633831AiP3hxihcqbi0HKdMblhaIGhTEHtA1nlAibwU1A22lMO19UBQjcKz
XVdbZuuX+mPkg5J5DxP1OyEobjrM/wIs+TV0+2iNSz5KhjLuzkgY+6Wg4PXZEzheQrfSGmNuj99a
qyTyPDfA/MdEJfZpelTlacU9bxdhemg1eDAJ7pbyWNHIMGQp63JZxLqd1B86EswUzaynPa/g1Owc
tgs1QEHdUH8lZmJv54+TQ837bc7jn/TwoBQAuYkbkXweReOZcv2VPrPX+YM2CC1ZqPQ8/FmnyclT
itheyHJYbdx0HSZMDhBpocTguCMhrVCpVqvW/dWGhFDdhy7fk/bqmKS5JCeqmjNdL0ngICy3CUxY
FpNK79Gj17z9THHycnqOe409uvoUPopyTbqn0JhWJT7jjiq8lg/Ui34nXin24f4KztbxWJ9AnJN2
fG68WyNJiTc/9BBX7enzNmTv60wJBLl4CmcXaXTDwOytb/PedsiBcagsRETPCjXNitxJCn1fBkdE
FnvdMtf7DoZf7IcmSIZEEw9ccQQSg2i6+7aJOrUBjNt8W6VI/UDfkEjj30FT/LauNk+K/LSzAXH0
ejuc30yAeIKv/M32zq3pOApBpSUDIgcdi+qrlLHG6Ru+fL4yl7x9g0z75YU71GyQvIGLVsqNjzsY
ekUJ60y8OakcmFTRrOKDrBkBsqOrCz4JjbQ835reDyQR1yswB7kfmYeMWmmQlkc4QwdKjMwIIvsU
InuAlds/95VUnEd+dQSaic8ZVwaMEPrB90h69qeQKg9aMcMILY1ZowKgW86y+ubDsCwv7pFw8mr+
QVA6PQn753M9pc9mSCjqzYxbOzYfUQk0qg1cdLXchL7XGmke1s7H4k9t7v21iKxm2rYXS2i8YF4c
VS+MoAbkiyLQCr5Q6cAbZksaEYwnwDvicGzdvPqQYAhb2SCdwA/rw+6+H2Gr4YFtwikPThWDiKuI
TLQNT8qPf4azzJ15cIs1KlxbnQAmmhANMtSIede+Q+821bpZCYr9x7W9h2Z+WQv/C3HBeyenFma6
PQf0DpUx2xnnbJ251Fkm24KkhxjHReHKOVpfwzzQ4Lsb7PmR/JKSZ35E3pAtuK4rrwYRyMg/Tz3C
P7GBRSGlCCbaLk/4NgmXSMyxV6k5H85/7p6WGtUcGtP0qF93CYAaH0roqfVzkIPIwJ6QpFwb10Fe
+/F0S/teZF6sHy3eO6WwsYbwNfbcG5sj7SGTgunp9vnUkgBbxqQj/s41EnfVvTjydtPYh/vn2+Ox
S1Oz28I7vKTq/LIjhjUrXwyCA5wBEV4WEDl5UuHm8ZB1gLDkT5gMBIcvbvyN7Z2AUwmcpTDJ7ETM
ykKDCDk600NDwX4XKFEbTY/A8YsD5ltEelDMYzKwz6LWcAtxNci+fk9jtlXC3LX2tTT+GKBce6/O
LBVMPVsJ873WPRXlcsSTVdZXo8ksYbjMYCQ9tRc0YTT1vEe3bUmKArqh4SUbW6omroD1ZVVhaXxP
R1JVKFWGqNvmjw/k41Zz/3tjmgce8OdBcvZFgknbY4SyNdwlenXDcvbZ3pjedgQk/ScW7MM33QMu
jIGkbLeucApqkdVCCyFCsk+gOBRDkvuYBDGvHfQB0Uxhd6Sl9pJLgm6HhAmsrCClD9STsOHEzJrt
zX2kZjJUoDJSK5RKxvYaMfi0Ws16DK9l7f4oS7JCQDyEEoB7dVQ+lhFnbsn0R8Ocyz055GOe7G63
HxbPkBYzoWvF3vOCTHtr7QgEhqhbycGIn/Y2nlwT4spnFftqcWWq0xAhwwfpw+YXkq3amqvKqQRd
gxNDBZYn3x/K/fr00GCToZqtk4MdsgfuMixpPsH41QMzwytMSYDy5Zaz/8wYF1ZyBiYtlR6O+Q7s
V2EHO6MWtGlZqoyItg4K4uYuHD/NPQjjASR8YRvvV0MPiHxetg35ZeTKwgrsGaJJi1c64nD9Y17u
Dy7hLiwsOdJDW7RX+xWRawth7Lx71hC+5E5PkHKmgzCNDSKX1daSmth6aJnJN/lFtEsNwGofz9Sl
vskQraqmJ9BM+T+DgYJcJRe5Gf5CQXXHoO+LnjHoQ2rtIaQOm0Aw5B0qzvWqPpeC6FR6ysaDiADW
YdlQczoOOUfTOxX9AZAhNcexuOa0mdm+Amn8WSxPRvWemcO7L7+HvFIU6KO5mPxQh0IYTaFVIpua
IiGJsT2z2ckIqTOCYjLqKDtmSkdQ6Ue/h7PYUPAuYlJZWcWbkWRX6Oslk9S3dZPPYxwD4GD+CTgs
EtAnFvGxpV9copE+h5taYJ7yfH3zBYwtyg/3h2cT2v/bjJIkwdg/rAvEnYyBw31MC7ASl4Wi8XO/
5HiMbu7zVvtqB3fLcmV2cnZ15sRkBbkh1cLTEjQIHDKMm+KrIGP6qNgeke7X4H602Dahl4FbMF9S
Ciao9mja8FhHxGkb8qJ1DCNM0IgsW/zIxxsdqLGdOQVCAHrTwxZ6XFg9kNqO6Ndwz+YKJJ/fwWrd
kJE2GEkIPA9+mvqJCk7mIyd3K/Otf8Q814X0P3JBQIuXTzA7xD00PZiKCeYV3PCYB6wVLM5Ig4Gh
+0erqhVjldSzzRpBRWcQWuXgVmsMpTctg4tdTqrpoUrXM8xGfcxi8VRmt0oXAe8On5eQxla/87B1
RAtEID/6DjlI3l5KyYG7/hjbSuN688d1mVZGeIrOEYhCJLyj+mA7rd2yUV6Iw0+EyXVfEc2DflOa
BRJMjsknHRnhIxvTDklrI0tKEU6wdmARxaYqz4PKj8vyCOP3vF8oOAOWiDLxLnVI9fO+B4GLxvtH
kOMjUz5EGYaf7vCFRmhiBkIwZuCzD9c/W/WfBp+GzpbU89ZRDvXtn1hkuCpiy21qDSpOaDi6/3uA
Idl3aLTHc9xMNg5HL9dfkEZwRy9wZOXnk9nsDz4rOJjm82BJYas9UTMgGd1jNl0pFmVg6gwXMRpC
usblr6l6jZt+knrXFfLNx0+cmC3kEwcRArV8pMoVgzjLarsaUFm4EzTNid1ke42FqKtuYCOaDaJb
0udJrBZ7qJMT9nrciC3wBjPJqD7mF4c6ZM7fR9ZEw/gN11hFhzSUCha1F/QfkhaVFxFi0sfhod5J
Pu54yzD28miLpnZsGxiriqA917wagL2IA9leXc+RWnG09T1FDN5QqnDlbWC4tLXA6LJjdzsJL/bl
vYlGgL/VFLVTRwgmeAioeeNUikRLGRj3zZ8VAlm7h4sLb1GV4QtM+hOdJo673l6M20a0iM4RLhZr
WrC7YmZg/af5RqvUUX4l/yJbrhGdvxiNoJ7ip+zJuecK+y8PqCBxr/5hKM58ozWk+IH19dnqi9qL
SRa5pv8YNilIXhego+gvp3ngB8xqGPaUHGGDoof75w2EKMVjC0Paq77/EuXQufuolSNywZ21h7i6
KWusOBRKkylAsW21xJvbyFeRvAa0DU7+NXYH9P099bgf6lXTVsNd9vxpdkPivYFqBmqsyKivE7+C
1fXWWLSaZBVDJiDC5PnUDrryo0DbOnuFY+VL+/ExymXZAalVmU91aSFfD/AED5kAhy569LtPUfho
/cummK43MEHimsFX+LVdwQtn9RMWiMoPyvxFyCR1+O+Xd98vz61HablPibdgSKV9Q09865WXphZj
1D1oVs4firSKw5DGbovBjO/446MJOUPi5H8e7sLVmFaVyz55E+qno5jCg2b9r5sqpIEOzPkDFIeo
LUfNDH52C0NEDun8bKvuk32umWWhMybOjdSc4uMxWGFMcyW3rTxpmxtgGW1FsHeHYs19KoZ69msI
CM5JcQZEpYGHOH6u/JTXv4hOeu67Lm6oWwL+w92lKkkcsHQ04r1ohP91oI7d3B8ctCrlO7bu+uMM
f9cIMX4gfgMqrJwzkh5f3W7CUx2wAn8Pq0kVDbAzG5FfwE2BF8yNJWaN8hdk/R3b9ct6dPz/KiW3
+jSZtkoYZVazxzAyECIsFryWch/AX0ZNpbiX2VOaHSLgFXwGEXrkz5LDYCHSWTapeTSYm3o4GYq5
WpsrDPk9W2+fJ7ozXefxjZ+HVs/K/lKu4plExHl55ik+9uZb+iqeQfGoD6XjapSQGC+X+D7ScD6A
3yJKxKIk+QfzTBd4nTgu9PrrKLf7VbcdQwJpN0N1198ZB2dMNaSAe0mPpQArj9ic6b+gUbmzQOqC
wLN/97ysrO5BTHMSR1lxnDWLlMUE6POaIdCbRxhBdHTtN23rwELcio0CmpioMr91ucL+BvkAS5BL
1eex/5FjYj3nfhvN/mScXJuAZu0iKEDWzZtCUKZSTisURkNJrviFzFwJjckYLyas2zxw1uhpc8Q6
lQFoZHnCRd2NrTgzUKViP6Q2UNgqp284ED5lH+g6IYAoTWatfvwA99RiJQ2O3BhfvYKPUvor+5eK
SnehTiiTKyQuVLh6TXIrqYW0KBz9kqxzNaSK2cJlNmugSFQWxW511yIzsaj6fjB6r0dwspNCjAQr
GsqEsSvKM6QU8M2+LYTWKlI8KKK9LyEKBXHhjHNJHPB1Ejl8U8P8B4IiC+5j0lYuWq1QtApHiZN6
AZY0rDi8TmZ3zUteYMdgd6Rtwo/seAhFIuFi6prOnqRFe2o2bzbtt+E5hFjMGkQuRsZGhvDEw9ok
CCzBexfNDqo0owdQutICR4lPgHQ2JbB49724/hPXa6OUWIM7nGvyuFcbJVtXnOJTfYwfI9VQ2kMG
vNHyQKnrqI0zeG0upvOYBilkd0/BZkpoW+0nmJvEVZFuj5OIkF0nJV9TNAOrKVTaX/wLi2C7DfCJ
LKxnM/yeMfkmbokwTI+1mJcPVM+JFHiudTE7QlEYotga//PWXM4H34QpaffPEC2tjADMkcoa3Lkh
wwazb3OKrqhQw+KPZEbh/Uiqw9hEZpdbEs/ir8SNB5yYEeuo3hAl+CpylfV18Gnm2+E08g7Chbk/
4Xj+I8x+vPpxsr/xJtOOYfCHGLFWDoeaq6HEimW8DLCX0PAnnHyVBrQqID+ZromcMhFxBSgETP/b
O4E46QaUipVAFjKDhOCGAvQRJyVv0+fhOX7+Ywh/HcinbRPUgBj5b6ZYA6R8Icq1oPYSxZfJJBcb
kK/5oc/btzyy8rCwBuVV0316Wn9waZM/o4aeXdzQ5LeLTImYjVQgZ6PfoIF3IvnrkBLt97RPvOOZ
spxWb2dPbmLREQVYWTJicb2ZhQD1BRG0Ib+dF2tjUEyaYpXwZcYujsawnGgwXvFeTAyXhwDpRO9w
E2u9H8qTlsQVbuMGANQu3Apd0JaJq+bGf1gD6Uo3vhIoacnWfGH3opm8o3yQqRipOV8hB6uYk2ox
/lVG8djih6ePzT4B4Sn4XG2GVYnZr1DfdefIAtaDkoNHp6dR+noZJxJmaC639+PtWBU2w+JSEWPu
uJo8zN2a9zmzQu7u4++CoPtvkczdjqbkJ1d0MHPkn4nTbu5V+4BuKgmDpAOQTF/HBIUA9BalbkLm
PFcZGRyYHe4pQBbCmQd1wsqBX8DeJGLNbahwEzgsTWAQalQCpUmK8xhZLWqHxZoRh+81SACe/BmN
N7NVd/JVv9aClW8UxxSwMtJUdgV5GuLDshjISrHyItt7aLSIf7CHRboTR6fwNoEwBPjs0SK5m1oK
WNkmjFEhBYwhiA/lCtwjmJwNPCJfiKxIw5nugxURZEGt+S51Wo3/TSYBzpyXzTXJpo/8nyvJoCcv
aO+wpSvMEZ0uhpw+59+D/V1b9Z5+vBrbCSj69AkHdmDgAu5Y/vsLYhwOr0K18ksXYjBb5wZ24NJ8
83SF0ClkGL8PqoGz1aUR/H9Fd8uNPcZRcVvT64Zk+Uk/BU8p3YcV22V1hkroz0tg3ALKi55ggEDD
OQx2YWzGhUWQq4eBUcAXrrDj8aaTw2PGF1AxlZZfHg/C+YAk7tJ0e8Judp4ogkUjWEsrDsnkG4Ol
yhARoj7ANtVBhat9v7x2SLG1sn/Dr2fVnVb0rQjNrWEN4rgtmfsIohwYoActj+1J6vaj6CGMIUMS
NDr7FoGwDxOSfH5ex6fA+rAHDM7llfvraMAb8yViiLcsOtZG4i9qPVIBNT9BdVJ9jGffNhYbn8tQ
f017mJZz6MBTKnhYQ7ydMO7BEci8TFUWbg7/+qWXw4hsR0RBiE77jSm8HMO1lrdvSmL83F8Wl7oj
TBVAiS/plgeMSs7UySMx28ywADoVVmek3ZxHSNQ1r+e7J/6I7SfVgRQczDCZZiFZCUAh4zMzr6q/
E5HdkYkfFOPNwU5gh5NyuSypzpI6e6Geem99YujjmX0wi0NT1MX04G6xwKcYOA4aZur9G+OF7N2o
pB+bJcQRXVmkwvx7quvPJwJoyOaYINBDv3cudp/G9/BW6RLnevzVOg0a8lQos5bsI4ynfWeyvZoc
/9YS4W3+XMF6WHS4JLIyYbUa9pQC8pXAO6GvnJ0Ex0vixVvhf10SsDQmnGkQIJDgZSGgdyn1KOKp
Qj2GoJduRJpd7aIGRg5FRUs9WHQHeBpoN4dO8n/EF8GQgzzwnMtI5gABjON1mn/zDv6lMrZnU+fK
T5LJsZbpFdOMwXNcxxVodwj/k8S92XzJrkERCSvh8AXbSBKk0gbfmO/mjQTM/PJnsQcDwYL2TWxd
lwwnXXtEMlSgtmVvRvWNXhYn3hzuu5qok8G37y7gtUe49RI7jM7S4EY06YJM64epYSNJyu649LCP
oZNlpphqcTaudQ+ypYnkeOqFT2Mw/10D8HnOeoxL5iVpihqcdo6ENpEHuZLYntVjwfVHBpjZoCJ3
0nFlnRt0JvWqqqHLu7utQg6Jdvm9ngtLnYdU9/K7tc4p+l1xEl2Mk1IT9ajWDSINzS4TE3oWqn6e
P5ZNY+qlQSP8bdhpILkrpVVhpICBA9RqWG1pywu3GciKRpodPyaq82BSoAguuzpucrVYkz3Z8zau
Y/vl1Z1YLzIZaup20oC+xP44dBK7tuZyMjmLi0gVGGCXAg3JjAVcpXEjPfC/D95Q+46UCCaqT2DX
k1mTDgzzaP30pbi89d+/OfFywAuVLxWydjS3IpbIJKEGA8RCkk3l+vqtvSHAiEmwOhtU7Z5dLQH5
o0JwTTVJT5won6Toq3x9dkZsTcy80g0YqcnvHr6Wi93gAjm6z0GDhRFv6w259urb+ePzwb2ps1Gn
7g9nXMvtS9OaR34DOcIe54VIk3RxHCOfpXTFaXTyw5qN/2lxGWPYSLevXdpvM8VKKxHjb6L15bJl
Y1y+C1/PihmA3yTYot6rWqbQ9k96nGS7x2ujMXZCqygUQPs/46T8JVgJo3Nqm3BGls94bxPIw7QL
K4sINDwoe8KM/z7oU93tIIrE25CEi+exn0gNhAMmyyNxH5Rkn42CV9cQ54KNdbrsu+A5cYKCXpEe
Iefqb3TjG5svJcgBjMc9ObzexCJEj1oeGC61hJhxv8U1YHi+G33f1tjpnRLMdMpcViBUtqUGpXkO
UIZiFP+ZPMHqoTPjMF4ibS62m3oopRcZ+LyM2eSs2NkHKDaqt08UenYhZIpCQdI8nNgdl49sBQI+
27wOY8lft6LjxeDfKKhSgE/iwMAMIzYbnPlOT3zHpx7ijRCWcRiZGgG3Ntq09WfL3xsYmGY2dNy0
+CC5A5T98z542sPUs5v8tSvVGv+hyZT07wthz3RAPTHNW3dxttpC+MpVQAqkLXpp15HZ93tO+Qrm
LxxluqcgSOx1a7CKG/EKzUYO7Azi99ATuklY7ol2i3QnngSXrJl4889MKOmlsc1RHRNlJoIhybJc
3rJMmJTUkOG3Um3W5/scdvd7sQELdm0dp9kHUcfG0dtTk+7YfT4jPfvq99kN9cwlkBILgrrKOFhV
eSYVAfHhdI53JqtOgS6TYkK7hrDjf/xm/5MbzZ5YLrtQDRS4AxkB5ExtOijFOgjogk6i4karBGFp
jzyWPMGrUPRuR1jclgJdstdtn3loYaXf5wjuYVaB5sFFsE0N83ycbrJLg2rv3Y/ScPt3TbJlV6Fy
pbDGlyT8HAUrGWVSKT3cMXFVTsm+GhXqA9aUiobwYJAZ2TpGzcf+Yx0NPPn+jLgi9VJAsqrGX06g
TsR6p8z/2b3XbUEHA+TIttYNYCvZ2TVffuYnb/5j1wWtNduLbgdm3Ev/dvhqrl3r7iy75p9BkfSl
+bQL4bG3Z+ckhraXsFiLctrSCS7jJ4km9Wl9X30X+DQu7xgTFXFYzTq6EdprpzFHQPl7oLj02LxP
sysgdRvZv4yaixwOn4fuQ7lFnqA6w9l8TyEbpRhnq1SAV3u28Llmn71pasJC1KfpmTgYtihrLCRJ
zANjoux7gDU07PESQzi98JRGfIJeYM67AglITBwq5rtzzQcMnJHJZ18ARLp5Le42ubezUAm8uGUu
UBO7MP+HjDFQUu6IBOasonTe9UCfyep19lCDdlhRb0LQUnPAOj0F99l1/y9UO8eHN/mheoKqY93x
6NEtXXyi8I+XzJJzIJZBVXeEXDbcxDFSRL4HOWJr54v79jPJH5bKHRUXo+jXoZqkNmUVT9Jvs+6q
xCE5eCtG4yqtcvfjPJfiREGDprNWxJhEmgLX32aguhPAYghpOmNsSTv7vS3QMmeFUUvetPpAXd3W
U2f6SEXpDGFf/sueioL26JRdp07yN+zQ8qkF9+riQkW6nDqR7wPajwLGULLaTPV3l+SSqHkb+xBV
X2veNfR0MI0txMgY0Ztz7dwzJZui7NquKhFAzdlj/btHs7SYYNeiVq3ZjAfiyxSAjVAG8wQHyGXK
P4qcF9SqYyvexemfxklB7ECNvZhaKjaMDxx+1Bp9vYvgR0JtRDYFYPzueCUw8Od+u6ku3boC+Kui
oOeiuV+LGp/1IqGXQXTRlaXEXOUob3DgyofWDkmbnz/W01gEnAiZqS8hO7rvZZYw1cTyzHE3urhX
3fS/egjpspWvOUqKtd5uqbHvHrt4I4j8nUdWks3R2yBHqzWYCWA3Hqnooq+jFFQQYfmrTGU7hZJm
GsgdeiExbJ4D5l35Rm22nVCB5EKFhsAIFxZkONRWBbw//cI95z1+zTHGctPz93GkoDsbbeksuhQe
8cTqYO33/vsyz1cQbEaTOSkjI0M5mAWhvn/faG5rf7cw27FwAK8K+gjGtna5fIS4vR0ElyHRDPpv
k7z3yAv426frvKwKPtPug69OqBdodCI2Cn6VBtmdCMQP8e+RinmUwqDR2FxNQSlk+B7ujp5hjP6n
Eu9pfQF16OD4lnlXJgYbZJqSdRHelLjY8g2yjvNFd6Z9ys/cL8kOQ/XnA2058/Imqr0oDFbd/4q4
WkAgesskA066XwkGHEfXRO9OqsOktUkrTGOaPPNnOZLaVnEr/Z7QsjQ3Wj/2HxVPfHCDdOnWQSCe
USRZJvgYfOBttei3WvSJ7DN+D3od+uX1jJPhccVJV5wwpa1X9VEQsZ84MEPokLW9W+YA5qJHIitn
07T03yfeIBkJ3NW65FLy7SCr4ZbGq1rWriPnm3s9FZfclIxJif9mYcR/7zJ77vaQHrwQKtrhyMV5
oWom93m6iwzyWajrqlWA/iFKpRpXa+v9MXt8ZGS7ta0YPgpVo4cmw5aWROqir8QaXnen9InJzlNx
zW3GLNqXGrDG1gOHsXNiaIwFaVArgSkk1tBls+zM2YUxq82TqoQwDP6ML2QAi0H6P6UyU+lr/89d
/hIJWnS4l94dC3/iFxo8FsIP2eCcihrl8jLUjpi19wzatuVpltNiuruf8oUc7eZ2cuNYn4f1IZc8
Un+eFBvU6egpjLaKd1ZTqTtlg3t5N6brMQEwDiy5fGClJSBJtYpXoc82fclx0k5PcmmwL8J5p8N9
OIGqQfmK5DQVYLcr5tR8WLzCNFLmrcCuH4keVQLxCXGXMAu6pEa+Z18L+2ESCdriOH8ng3cFco8h
aBk1kIsN1Ldih8yOpMj4ZE4IZyAmR5ghmpyZN/jL+pa/mspCrtIyzFGRGKS629Te9uHhAkZQ1+bx
D3r3o3FoZTEdfOQb36jmPYOrQWK8chX9YeX1q2cJ06Ldg98LaMcT208HmA80gQtBdZ37ofwtx5rq
SEKWcGGFPi7Uf4EkmIhQmYzpC0otQZE5qyGkOfzEkz1/2X+sNNVGvdJ4lY9vrUvuk3LtsPAt6w70
9feTlOwGJ7mX1NVPx6JO9lacamXYdpThRP2arjRa5eYH8CfveNvWIfq1iTh5h37Ngq7CLl8SR9py
UPjbtu+Dp/4NLwXvNw+7arbU5u9pjd9Mfpa0s9QsZjok3TM6GQfx1bTYmTbXYKiIEYFpmXUEiLY0
78ihYoorPGpLnoHMzkmplxbDRpNT6hv3Nr7zHjO/12klNsHTUicA66mh6MDBWHV7w6Ay7GVrGLxE
TqAhzX4foMnoEeolF5rJ0ODJI2V/rXQDDjVGXn9ZBZRup697z4KCIrSvT88SKE5PThFJEc8LiILA
WHPJGMNNVbgvqkjVdMZuKu1Sw2AbOxR9WaNxbgpk6fur7Q901pSCVNnZpTN71X5T5sBVd2GvemFt
QrDgQMhGrqIDPq3vbJAZKR7lAetJMP03ksozC+yfZDW7YG4e0XYv/CKvY3Rr3runL7S1GVoMRhqr
A2Z2T6qssNkAmM4NlqeXLzVblPNBOyCKG8fNctyMfneVc0XJ+d6DVxByu++ZWjw3/9HcRlRy1RRA
GG9Euv4oAWOg5jzHuMvDVbKckHhAlmbiT+xxWRmIg+QYcSXpk/YEAT2LepT5kPa8wbrivUIv0Pty
EVZLtd/s1BB6Rsxg2t/TFwEiA4vpO1Qlz829JNCEur0GaIkhAjv1iPB0kn/Jag8LZs4R1Pnfv43Y
Q8Ek4ueQVV8beJMJHhVfV11RCP4P4oaWuSzh6/c+pXgRSVC3/UNArobGTE4NcHBjPoy+koy7Nazn
70akvPQaEFHqd2cc9Ob0WpkYqgzyzb3PI+zYUUNW9e/mInmnvR9YPsQqY1v98TvPZ9SI6V+cUonv
CLvvZaxM29SL/UcCv2IAaixTaOPYRZPErCr9B7UiGYFTutyxvfeCbxF8IjlBPOTXdy/4c+TJbKoy
7tlfaCEuo8RWeUhwgYY4cby9XYx16Z08Hpl1RMq5mCeKymPjNjG+qJzPnjdHUW4mhWC9fr8I2lV7
e3XQPDbjsvUzDMkA+3OREOHZFlE5CZa7ou1mdBbrFQJYoZAX7L/9qmaH0hAPOXOqml6+/j29ZHuO
ydyn7yOYTU3S53UovjvrepPVYmcUh9OqdXx/QI69Pae0caJPg33PX++L1ZZtxjRTH6l+UO2VLPFK
A8FHoq/MwS5jiiEe8lCJwvJ5DIxEF2LrlxuabEhQvDcloURayJpQQ0CeTc/KCTtUAYJ4grt28eRP
p3oNrL1+7g0pdOkJCgHXsMWaZI3HiXbCoMG6kNiuW5KnRg9JU18Io+S8ZR/sCWTa3hzpiOIn4Pa0
vCLwb2lNrSvEPI57ijBuYqPIu5Bxbbo2pnr8Rx5jzkAq5/1/+VQqtJYT7ut8n6KDsYCtPY0ok4ME
zS27LWzi+ELPRMS838FdrGZanjP6N+3JBHpLGE29P28JvIkVhtoqSYr1SPUmofNnrEAlDUvdeB7x
oUtTULEb7DcrS4BEiER7QBa8TVLN+zl5YmGmLZaRI4AbFAxpjMF9o/6impcxWsmyhgp+vYSU2EmH
HKaf475aL+3S23fU123QWKUqTj8q9n0AQ6dgIcAuzI6XSPFEfJh5EOztFAX8s+Gho6HozWHTegD0
V5bwrPfp3pjv4Crx7zHzjlQHAQhGnmm726Qmm+UYDXU/wglsctLSaZCZ0PffmaCXhbdbRCSdUewg
woGo/lAr3xgLZDrYZ5JbHRZ+EVSXkpJ2Pc9uthXjpUgvXMSVQv1aO0xgCLYy98NCqxjakQTV5BWY
czx661MwJXj0XsC27prXMRibwHE07yTiLvTDVFkmQo8F6S+YDfe9VT+OapYIEi89ee94spS26gPk
tvHeod/TDukm4rqk7qe6E1Cck89rh3VXACuY1PENz5wRLNnA7oS532vZmyTVxnLSwXY1GbXRpc/U
kYglRxRmJdO8xq32H/n4ishCIqLE3kptUA5f24oeDizjM3MjHqSZtvvSxqlKtKlkT9BGHs7JV7LQ
z4tYvhXYN2khZPUpZVqSXobYyyf4VPQ37efDAO7Yb+033OKJmA81ne8VVtQGdrUQ2FccZQuiu1cH
eWoZhxG0gVvpPyI7d0X6We6ioYUv1H7GNfU87noFJ2eSg7wrJR/XqeCZvncO3LRuOlaa/5arOv+m
TBwzATeTD9CntujGlLFzYb5EvOLOHOdhbU9K4KL0qghjS+UhXcVG+4CaZDnP3FenXItVyF9Hn4bt
cEJrnjBeBCD/AIenei8OR9oD9JmZnbwoIanZ2iJJUdsD7951bO3ifEExMnhKYjyfQ2LPo9qpuIea
OqP9f6p1HEOP1jyKZvRwXLzV1xNcmq1CWwX7xmZUdE1tn/E83V6+sZAc0685OxkHMgceJd1fvlMv
LQrfcNLqoTkvVIEx26bQR7OCBSgc6VMnnMFSz+uRK0WE6Eiq8k7TWkhz/99KctDdYYPC8I07Ivhm
WC8NPdOrt5M5ThsBMRQc8QtgTO/nKp2MsdG1d34M2Uo4t5e6ddQ5qSeSPrtvTNiwkSo9Qzq+4122
pnSr6S6RKPxPuFEFDpRWm/rAzREDBFQivVl2zDi9A/f54CjGKdhBMTgcBLv3kKdDx2mZu4+siqGg
VzwSk9rmt+evkl0snYeTOhBRJls3nScuogodFUMenhfGWaEvXvbEDLK0z47CqXmLZ1wGHejUkBm0
HpsZU5vSZy+xujJwbCuuZZkEqZj2ZrozlND+6T5BoLXkHdfw3kFNNX4C+bcY5IPOvBZmt1OBdk5g
mnuvzr+vBU9pH8tOfaSUSZK6qQiMTQDdHoq/dJHI2VtXdMP9XBO8HpRUOrRjBnQfZqOsX1geYTPm
PdiaCMwkRfC6C0oAakwqRPW4zKd+WfirsLqU2DovGDVSsejK5sPzeenS4D9t+py9GrIcVMySAtYe
bwPVQKXFn7Q8VU/lzv9l5zNo4hZ8vr/OYKPTxEPbNNK4MPZLZHotq9fICxNGzYJrH/QZ1JrgRm8E
7IG722E7AfAIXVMiLPlyQZjcOB0HVRZ21el+PEZHPkQxqN1za5eLVEcfryOArcKMWaKq1G1uYXG3
R0ajMVJLs5rqmgsLbzVFspBylqx+SKPE2Lv5owuV1t/3jACaVwsmvyPKKJalrEVkmKwXEo2er92w
MckDVpECpQqHQnmKOLAPTYm1ESZoaqOZ4McKZuSNZ7uLrcbZfodKT1mf4jJQLbIeYaBvwKvNq683
gNacWVgQiRU6ruyDjjhPrPQyOe0ZNkY2kfbUcivvOj5ymA4psYP8yttGBUDILtu40e+accnHCOEf
ewDfZASS/mgz1CXIQGNa1VsD8+cc5J20cPFqj3opFBEf3oqjJGy4hqs7VuL22kfnWj0BXt/KbbuH
uUq3n7OEeR2aADcNwl65ieCUKyu6AHC+M6b2+zHd7vzZV9Cmdms10MFy+29lwL2rnDdfX4H0dIUD
n2lTevg0D3Yha/g8wFDqKle1c2Y124JWFK9TvyU1Gf+Y68PV/eUM+hsPXIX+sz1GA9Q+/MfMqiWM
Whm1e9SP2tY/YaML+7VhpO+oS1eS2eLO6i/mkGcZiW5zKS38ZwpUMpoAtHeV5rk8Wcw1zzsFeJUH
e7QrCREBPVoANqtOGcUKZRJ9sWrywvMogVnH8//hwmSvEn5zYuGRsU+T8diWOeQCsOqx1hJ4PEex
gs+0PWYvNnVhjrqJwtOYKm++sVtUOpgic0pGxpCdhXgp8LDaXHJkz0PstCE8mVGCXcLQtPuSYTwp
zXIR9x9i7K83/AynkEJtHzKNw/9AlS6h+CgmTcKR9AGpwn++b1WVBUbeqaRWqRD3tnyaz8ujUPVb
9VJXtNcyUDwMfFqSjDx6YGaEcR7hS24ByVvr1+1ekClh1fqMs6W/aid3H3BMLPIMVgS3gHqREaVF
UJAV6f8RYQQYHnb528weHENmZMo+tnZZK4DgVaCYJZEQ+/V5WZtwctvmxl+/Q9kgYbgrXYer74eO
rciam4p6HdKKLz5PVE8kXClGS24Z1sqWbGnBq2vYGM6jyViasr3KmYBmhmVYpjlhPpqQHHdlqhHV
PxF9voHvJZWXFEhFEMA2v1l9avj6wEWxrLALoLuO9OPNYQnZFDse1xw+TuXH4m6F29tw4tWCD3Od
Vq31dO3eL77nvOYhfExD/1NFRAA+hPnfagoGNnEyM1V3fB/d+Hy60tJIzsS19Vu4+1KoXSy+zFif
Ib7IH8SKYExr1f43KYE3ezYqK+tLm/zwGMob2nayiSGXQ9SGMlsM6iAvGcG/Yu38iVi5VA8lKYLV
XQZ2fv354bUfWqel1UEuLE9ZpnZqcp8NBWk66tmBgnMWSWox8ZPzSTyOumA3jMPqxdL3W0YMJJuk
dvfboZFCTl9gIthbHR6H2WLTmROcLtrcci0jx1RaIkFSit83qiuf9Mr560JFOE9n8VCRXs3ApjUr
H7NNPJIRpfzjq2ptDiYM5N7Xpw4X26c/AD6lxsliEtBgw2g3RHH/shtbnAm59jos0E8ZNptBorJ7
Vg0t8nE59rLabxYu1/Cj1FS2S9auzx3mU9GUsoQIXz2Xyuho/7gW1jiMpkM2ESGMPAxYQCxglD9V
Iaw0UtxW5NbLyhw49BaL/76SwrUbg+62kDWvGHkhA3wNzeoXYO/DIcdObgwGkxN5TVWXl08sXN80
JSD+XMABDA69kNGm2DAyUA+0nWj9O37iTZSGAceau53LcktLZ/yTFIq4mdBhaTQQosGcAsE/cvS7
upK8EIBa59p/IQjlbZSoEOGUbtJrNnKhMTQaQFsJ03f+hGYYIoZlXrycUEk+LPdVY74r/1qq47ou
9ImlPbaLAGq2qnQhQocINGWbHnBlKN1b/fEpSb/zhod3r+R2fGo7nt9sGLKUnvDnqcOgZsevbbez
gevbPRVGMbNuRB8g1dek8mm1vWDOuSKH6Jw+MgkC4nMBTFF7CrOsYJEdYJN/g6u6g9MdwfqEaDUb
5z4OFn4nWTgBppQ1t3uiJI4dOCeKSESx3F2YssdjHvt9WJA3KgZ/oK+wEa4hscf9EIBzVMq1rsvN
SK/+D6eDorxg7A2wFMIlCROlwPuSxysfOS2DLIQsAuvjj47logHY8sLMOT8fzPeSwipQE5ZLctwa
dbzXhZu7wvI0LqZGq2iE9zS+7NfO7usk3PzVcfh2BkhuUGAaT+hqK5fJubPxN6GchXyCmQRP8ivH
N1q44uqlnsg9JOQ6rZVqHwhv9gvaFA+2k646WyELJaX5ERm4OR2WajRf1r5UGwrsP4YuXbANndw0
QP/gnJnMPKNrslY0SjaC8tbaR6m68oApxgyt1VMPjVYu/yYIf+n0BaVPa0Km6sRlLoNFZtgahNHP
TLkMtS4xJokE+rbWpu1ulfpDbs6zuNfx9cdDhyG6r/8qhCL9Isa1KLst41Bga8pQadXtdwkicYE5
wp0ryI7jpj5wdQGO4tLKF/Y3KW532VaPLDg+N7haIFzKxYow7KlenlzU7fZNOO9VDHGXnpA4BnUe
7FWDpPk1hhuXt/yK+5GievbZc9cnxjQItGQIrS0M13xzHzE9NILz0bY+6gZIntL0ozw1eywvpfkp
hM/i2A0hHJU5PQyMzU1yA2Ssz+1MhNs9LHryZS+HnZfZTaIJLi3zbmDXOqCUiM9AkvP1qgqlYa1a
2iDz7XqapJqPiquy75Ki77EoaPGRaGZQf7NQ2XCQlVoFsCCfbaT3JFf01/fPfwLSEz89IGA4NbF+
yAPI7anKG2V7cWNKbXwqLHQlTLBRRca7u2GK0f3PFJLVNVr+RgY8whehDnouCeAK6DqIc1/9hiBx
WwcMe/7H5e/wU2ak39wMRSMMGQJdba0jRbozhITlSZCAsDuJf1X4SH+AphDxSa8U8CzkagMkGrAl
rVqz6tRtbBrsICe3I9UqQo+7QeRCCgY+R4Zd0lTF2zpCHgGkSt41gHyRAQu1fju7EosWdWAcRNXB
S9R597ZWarS0HXRDK2MlSsbJ85cGJ2DUXs3Oli1pSQQt6tJ5Sns1VDdShwXs/SmbUcPlWOE3WtfX
gWeYhSdBwWor08JVDfImPyhLTI52m2qJ1/1TUBKNby+N9ybjjS2d/AG16BiinVcf2rzrK2+JyiWK
JB2YRX8K0CLyfrl5IYnJPm6A1kI8QDbQouFoZ0CU/6utcDptafc1LLLOWEDsSjFxRv7yiZjGKBFH
VtoChiVar2+ojcxbhl2yDvZkBQxMLRaQr+3dyQLIu5WpqpYI04c8KOtfYb5dU5qpbANgXYA8br4T
sr01ESCmidOQxrRynCihnCL1buzCvRSwnYpReiOKbKGEdgL/mq6sfuG2phRHBm817qsORxvMovB8
3lpgE9WklvgEhsGVuBk2I+VzHinVu3aqpxQzuM3tz/dx7zICvhXGHbRdNM0I5YwOyuWK8Glq6hJo
it1aUkJsF6rVIU+xoc5NdOwGBoIrp3HQpVmg16bauz94SGkIZhsz8LRI7MUPt1tGuD/mgUYO4iaj
jtJ3E8yELBNCYO3KdJZmJLe/fdcUc9nNctngMFq3etes/0LLUce8Ac+3VfgPB1sl/t0xY5fHi8Hu
RjuUOwX0TJ4S2ds8ST9BmNL4gfbnk1wjZpNLqu5xA/W8hlcbSoPsF31nvagquyMLSkq1+FT54X6W
AtXP7wjLbmhqp9ua5ScAse2bBy/y56P9YGqa2Bvxq65y5KcdwnvunI4qz91vB0ynBy2qwrSliAPw
W+9s+rGUXBnA9zx1xF2jnM5eS5IPZdYoeUn2XfePAmGCwSRkVUlh7RTyMQL863uF0uqPiO7Oo4cj
v/tBQIkgADa5agkhngX6kMrlZUXkwtit2dNCuwpmQJj4NidgN21fmz17yHN6EEIBmZW9uy3x4n9e
qhP1jAZt+fg0cvTYqJiujE8kDAmbd1RMItUjXdR4MtJywyuTaAP2xR5dkwHGORnjcBlmOEBf467R
96pcwDkrTDd/Ht9ELaSjArDNAxSiUkidZ/ZxUTkEb9KNBiglkFqMHLg6RbDwk94LpmOoscRm702e
cDWKw1HsqBo3TtWmbH3spKV5oGwdpfXp5JAInzARHpyd0Li5rreu3ZYzbi0lUkpe4WyenNgFunoc
OpFG6qTQ4Oe7HQteqExntVdaLcCA91kFggdUi5t+0aC29I/I21P0P25ocW+LkP4mc6fI2ky0DWHN
9/7GKiXIEmatUj0htDlO1pVioPbsdHh/51ii2SIEcjl+mFJta4dA7vTUZOfRzIqMc0CpZ+1g7Tcp
BUF6ecapwkcm+/W1hWOAWihME5ler9k9bDofxBJ0YuYWKtBRZO2emsHm1X8Dwm/MqPF/FTO7Ds42
C8USr/q1kZD9Uo9UcmEGVJZylTh9qH8JxT9F6URy8h6GlPZk/IQy1rhA2xssD85I2COe+bpEerlz
QgJ5CXeIY8Qnlf3wz6zMKJebSeRDkZpu+ev0oDVBUShFzJu8VU1eyB7Z9j7C///zbkZG+IAA58uE
GyQRfnORpBqF5jfAFEYp/aIlRA43mI9sC06YFPP6gSkNUr7bmPS8pwZNRgZpJUyaUE6vb2duF0SB
tfKQWzP9yEDR/xdpw5+SrJgBzK8lNyb89ATjqkSw8+RREjrr+qVP685SzFUYYMSIjK7uoAAVKfuK
xv6ghZ69YBXjZ8eswTQMy+AcAsxffj8235Zd0CYMkdwc5RaHOXD7ha7I2gMqICC6CBQP1jyPvfXH
9Mhwx2lXywJji7Q9AkMR0lG0lVuZy6W8MGauUtxw8DEPHa03cddLZndg7eaSJ1VpSIE5Ql+uDnQs
tWk6k9CzsCSyQROI28pygdX5P/ktn8QAnm4gcQ7mZqxkwNdwhLGt5/5lTGwrc3SPXHjszB40mW5l
welyKYLss/Ymr251sxtzyRmB9bFyjsExKqXiMhpqKmoRT1iPPeza9+uJsdP25HESUwz602RWfhnh
JaG/uqXegtFb7ttcSqIkeRhf6WRdlcNG37j5tFlApPIKEq+LaTABOGrH97EoAm6X7MM+ZNbO4m/O
tK5JyIjX20TONySVTXqercT//EaGvVrr6oZhdh//cMdx/hdVNkuXpCdMeHkdvn46x4IWlOsZTfPX
+IWboGyZyEhQBKM0cN2J2umcLBL+cQCsGQMotfgHTl6666Y595iVYs24G2nC/hoHKDJGCPnHPjZu
SUA2083j6C8evS+8YajwXtH+dRqK5jtjPqNsmMdk3Bfe/HitnHAKxmsuE7RQeLjSSS+NvsHaIDp2
rN3NTheKnPZcMKX+V/lIQiuG5ehPOoaxbThcD83QRAbZ5itKIsJiwJjwgdZNjyXPho/mKb2S0hpA
OCbTU5Ok/CXGGVWxbQoeap7BlZDfNAfyZCpUicQuPEiLOz/p+x8NqN6Jan2WSrYn4rViZ82VrKSd
Vr1tHoBZHO6j10QTKKLg49zx9H3tzAa5cjQDe/+MUXn4AmCex21QwZerRRYOvgWuHTtT/spsDF7y
ej+RJY+Qx7hT05e6VMShYeP4YSYdprSDvFklCJyinGSZHW63TzXFd1yIxPy/Ugb6G3S5OKQYpfue
RKeDPAJTagQP2tesanfLi0M9JxUQ8VmqbV3Apkhnp5TK4R7HwPiVcsnXP+igMMq/s+PTDd7G9mF4
AkD8TIdDBFH6/5T65nvZEKTI0f9/nuzcyj6OXTr4mLWufxfLdK9IgX5O8OBptQbOdwkJfgxmCKrv
Tkv5txdTZp0lrjBl7dtf4iMhteRbM4/GNCiEE1hB9VszIVM8mVLwtx/ZinTxMxOOusUT5Elq9FtW
Zge086QAruXUmYAq9Dcx/Y1SYgejWoxKRClKvoZ4rYa3yXBY4vYp0PPhu9KukLZkjchMHJo74igN
jflz1y7ffX0XqFPyuOHY8uBePX/Pmbeu3axXmfpoQ0bs8YHmvh4badSZzNOIwONIGcRRk9DtAg5E
rbbQdEyPrv6aEX1kZB8teaLIN28b660dLd13cd2XBdY2db3v9PcTKh/cK+auW9iMbSAXBuiUCgzm
J/ay6bGJlRZdrlPtZKFldRr/tmC6lQFBxILyhQ8lzNXVvsI2JTMxYYJrp+8fv8KKOS6ry+0RW6ao
2SR72xlkGpCyKD5bFnSMkvTKLEcoXEzF/bovPYTW/PEHheZTi/l4YZU6Eeij4zhkMVnd1T5iECtQ
7D4/r1P6hXM5hhx5hd/v5ETVTr0qq0CClCzvPIfbwVyIujxTzfY3k13sbkwgAg4LdpnaoCqAXpVz
4XBV0hEFPzTAH/cdBhAFjhwneB7YGuUT76Fyi0W0bWJJHBrdrTw+1FxrjUbnJixa7Yq8Il9ef2qb
33KmfD1vDYG7jan3jWGjlI82fEDnOCjIdIIPEtaEYq6y2mthOhwkNn3QrdVDQuKZGGofx0bjL2bi
5GBM/rK4eEmRXMi3G2FV1fJ8whWnAxnZyrzzVMlsV6rsVy1gTWQLzA13QWmj9l5zxyVE1eUqlXcJ
E2eJxFgDkir4snnfRSKFR+f24ALWkkmeqbG5FLd4nxaNvzay6XTSPN8R5rDs8Whf96Ri2ZFxQ+xs
7x28dKBtY6Q7QhLtzj4n5N0IOBL5OJeU8F3RZfwWQM1mNLZV+VFq9TPMwydcHw/j2LMBjgZ7MlEX
G6OLQ4b5cQUmbxXyhJx2liL0ukXnjtm+W3v6+KMk8y3m/Uis9HI7bzurWrzS+d4bALfmGsHeMfjJ
Z++MhbcgywCOA1dHBFW9P67xGQrTjmZUV/T2Q4ZsmTx3wontna4TtyvITNvVgGB6gUT7lR2t+t17
F/ytOq0uD0Z374k2xKSW6m43HWXADDighzFwYOmFkCpHgoRn/LagZxRvn4bU8xiXimG8L1eBY1R1
z+ZsoDIfMVmWbAV3bug0lZyrjvQWWdNfbnOuR5UNdhgcpIHjh9ELjjiL3H0GhFkJ99xwePKalcu6
DlPZLlmI5GBpV7hYTzvWaSvjC4tXnlMpE8fYxcn0Uz1W5+z+c3ESkgtkuxnAZqpVvieH7GFrgXx1
UGOWYnFwBmcolMewOlZ7V/2v/I6ELrGlvYnJzcOdwaFK4B+DYSSAaEL9mMTFVn7NbGrFBHHfYND8
UMIDDWOBr8K6R5I+jqeVUPNQZcpq+76n8PnMaR+L2cwJ/KNYzApnAsu9Iia1IuYs/YRpFcOdSt2+
P2D1qt3TgzxJaeH9ZSTbDw/dt0d46CWqsV42V8azB2/at4ptZ+e4Snu/oK9elv+lYATRCrq31jnj
9KH3TUDG9+ZTIn+OYH9eu5SS+E2Np4VxD31iljRn0R1Kxbh4ghylck3F9wPA4Hm/t8RfPf7qAR6Y
lmLHlulyqzD7pG0zAaw8Gmw85kSoXg5EokNC/2NaIs0oxmTqJH7Svr7uhYEfKVMgb0Jk2I4wZvfy
OdCfoLE1BDhNFofC7cE6NvXfPBMD4bbC6Or2DnlDrBTFcddZ5F2En1zANkCC/0VNvFkcFQVqeKAN
kGHGtbm71XUtUzq1lBuPB8z7AjzB82K0c5g0rqm/J4iBVIVgQEFzqBLbMkWH7Erogv03HRzyhJ0l
2KBm5Bn0LPeZbyvwpnjXAMSHkjLkEZCN7MznXUiZh+9OgVG4J9IZs14xzadoJLysnmW48KzTGB7t
uMb0hbxPNgmi+AOBuq5c52+NRCEa3PBkG8kkf8dv002PQNQmlbuWPwyxzrIe44gHEIvpwQEpi4pT
m9zVSd53lGyenyy6Z/e+fWeZOdPTYXg4/oV1nCdDhZF8OF546hDtIAs9eSFsXHGcNleOqXqimMuk
33ABVfC9r91+H1a36lbmfywkKBM9TJCl6RdjjKU3ubYR3omZ+lhna9uqvY2gzwHGTdJEhY1PZrQx
3Bbn5/ER/uPNKpwv5Z2Y9N6B/0gZVAivSQKIUPiFiaUyYzk2USQDeQ/2E3XNILNfy8Hw5pchFaBy
BNgO7V+wDoxRT3ETxzjZEQSCR2DMX+e0suEnLdACXyoDXh2PiNjXN+ZjkpDd8EbHClpx11+8a6kD
xLFh7wtl6fFZc1tK7sPZ42K87WeIr3MUDqDMqkIDq8CFQs+k9jHNaowG0kkxWQ0I60Wgh5Q9uZVY
VOD9CIUSUdzLJv17J8HOrp/ZM6ozGVIBj9wNlOvnLnnQFS3VpBGGOxX9AIMpiJ1n4qfin7ANEdRn
npW4lUx78FLjF+gFtv9USxIz/WreNMVOD8UQwjfF8VFWqF+KAhkIWWETuNIrys1MavCWs3fp6hcA
ZPUNCdJMRii7OqCKz5XJ7icBDrQ1bnnSp1BPuOpWwW8mBNmkZfeCg5ajeBpGXUbkey9m8M3JgX3n
ppsyO6rzfWwyH8cLuPyrU9nFpMmBMS1A12+dBo37Hz82g8z49n+UxgmYJvV/rrRuLkAjCSEdKo/s
Cnl+s/g6rJeSWX/JWzPmUOrebcKVD/a3/MaKiSAKnvYu9AEk3LHjbk4CpeqzBQB2bP9hns9DSWfn
FCtEQbA05ig5zPsJdz2CocOCk9Uzp5xS8REljf4gSuvGhyzbfRK0MzNQwYDMKqvTgbnEHK34MjXo
2NmAiVEY/3JTWDCSSrOf8QxGVcSzdzysXxvrSLjJyZj48mUYoYY7fErxnvjtp7t27Q4y3XhR/sUH
z4M05xj1isqXc99CG1VirgbfG5Mj+dOWUhkwxx8lNpd4z0LGt24SkISVW9v0EsI6c6OxrjbakK/q
FrtteJUWEdWQ+/5eExL3Ev4wGYYFlRu9pixNhSji5OZuWpqUQQA814GIKLJgJ1+0nsCpRrZKZdHT
ySF4T3/J2AugBVOt0Vw5y2NXXwF+mZy9n1Wf4wbuU6vng313patBfep66DoD6yoRLCZCVX/9MuaH
vVshdQfto/E1SWw9R3Gv2P4x2V9cgXTy6+SHW0PLw+wRAnpDl6mS/Vfe2/4aDPdadSFEp9F/VljY
fb41balGN6vTU2w/z0Cxt8Dv4Nrvk2pLVp1hLI0B65oNKd+bXGCizANpXTAJjT6WFfhszLhMjlZP
wfRUdhdaxmv+RIK42CLQkFsD7JCvHr6eKVjfVx+/j6Etu8YRNtcbeRY7lH1Su7cYVemFBL5iahyt
B1k8uufghP88dEtGAF3tGDF/om9/ErEjs9E/Qcyq9U60ReHbclNbHv1j5xSaUUrKoaSPSXScSi0h
eX8K67hXLsFlCP7vHBFkSDkHlc+1KnFWzkmC3xx2fNUMbXGmV1xYofRloZfgZ3dhZcsm+fKEGHJU
aOUctp0f3+REgE4ycCSS9EbL3znp+Q+jsCSLR8NG/sEjljeVVeETtF359zjPumm20qk4UR/JIR2n
/hohKWGBktsTh6xn8UJoeH+vo/8UZoSLF2ssRdTotv98A8inLRwhhVGwbycZtG9YVcqEbeAWDgj8
ZAKDx1VU9nK9A46GKUOHL2W2PcF5yGEsV77uN7GgeuxiqFVxwf8EomWU2d1Id33dWkS9zRx6aXfW
4KV8PGn3IV7B9n3N6lUR75eZuSPqUJ7llrz8wqibeGtWccyxQ86zs4gvYEMZcIhz78ybTNaAH7F4
igaH71F0utqggvBh4+HDWe/q1mDdrDg/8TRz/JjpX1Nv5EWeWt3IsXSSnPuzqTQyZ+yc4OwuKOFS
+NNgK8o/uhTIvR1gr4UhjcVYmZUexcpdKAGuKI+BaKWq7fPzhDbatvR0lh0YqXx01WiV934vYid4
91BEFsHZd2DwSqfYTA6b307xS7/kxwnSkDN7aFGloqaGkySPCFkYOe2zt9nNOXb5PJQQ+W9XRIaT
WoawTSFS7Cg01cqsQuJYozHXBmkK9bXb4WzWNpBtZ+mR7Nx4rXqcaNgHsfNA4XH5xKGZH2x8W1mb
jfVOMkbJOm8yEh4vMbDHSLCVLf+1JzAC74OVUGdUq/XoHM3YPKxA4jExlf7TbEyuCluLvKZXgjKu
WOxhsxi0l0x28W8ACfSUurWcbycT7fYny8MOsq/ZKQP6CXAjjQhKo/fIszTT1fktJlbgYfFFbuv7
j4arHw2LTx0AUSFxNMlFMyu0L6s4bJQCWWfGE09CfljAvPEkGT2iHeML1x0sNW5aaXPKrCjsAIXm
t3gH2/D8B13VlzDB/JMNUbPi3fglmhkrSbbED4+D4pWQ8D1F/01BLSQBkHj69cU+KN+LFDdb9k4A
7MF+bd2QkYl+g6cNqvGQ7H23gbtbF07gyT3L4yddufG4BVtzTyZI1MgcNng3Pu7T3gwNXdIxjYDV
TDxzbDUuaqfvpp5rYWzbqkxhXHl1fEAqs/GwDbFH4NvSqPqSld/SVPVBN0JpSotV/PbNTllzRBLo
3A0K6uCcra5DZEqy2L8+K4L7cdV7n/7BSN+6daHnvvAdDYu+nKcBhDMooJWalT7KADK+UaAqemo1
z1Zmc4C+p4W4Pb2OgkVKqg+cyGMlo+CWijCdYGmw6j3qb4m5ybShuaPLiK2wOtLBGoWv0K8RLrqX
vjXTgpeOuJEpDQ3tTB15NIYm7AhIJEOnqwcWs/dwApbscXPo90E0wPWgVAimkxLdMbPAjWlUUG3u
/G0TBDMhKrQ8lbMLRNYkZhYAEOBDHeAY6b5Ejeo72ggIbaPnPdIbY38Tvno3bQPpkBihRDRg5X29
GSk3f3h/TkbpBSK1qfLiK3WsztZaJs5AZrOn1g3b8jz76aTCdHXA8ZanNx8w9mVABRfaVDwk/Bh7
oaCxzIxy28WoCguP4h98v8XrfLJi28cD7IXpNznFzo74TJfJwv5siIR3I0bamwzaUpItN/D6rhkw
k87IVG15DvpGZnvCT7SkSytp/1M+WjLb5PMcOH+LUDlijiVef2FOTMEh59bj8cPzb9+rcW0hJMwr
Lkuzc5YZuiLnJGq5zkNspLAxOR8NN4LC4mYGnpkoqHhCPatXTwUEVv8EVgw7C2hAkAabKGwBjETu
Zj2Hw9OxaOZJyfvEjawtp8uw9+di1DhAEpJrz9ZFBHQ8gOxDJkwDRyY7Jjrqq41A0dld3YRNaPCy
Eh7r1N3wQAqMhWZXVopBqI4u0j8j80rGSX1P3obdaN1+195Zv7UXVXBhRl3T+E27lcWprM42CpM3
b/7jeClNHGeu/chXUt35dxLvUlaqKkSxA7oF+2ZAhuZvMAk1JGCb+Ih9AYU7uMLwQFutYNzaO8og
BqV8hkiqbhkEbxwplsjswr2YRE7gm5mU4mCPcWmET2GA3yaFq/3UhxdWStHnJcuMbcgONgGNffs7
3L4SLxPYlrwyTxzYEqMBoSJCJxgPdX0+OeEi95LC2BHgEhmM5lKAIySfCET6EkPm8wkT7EDQVi5Q
9rW9nG0oWRnKUpum2RWLHhA9RL9764MlqlwUBOvzWCnrG1d8gMzwbObfi4ZGKNUwt7Bo3pBIixf1
bZNEXNVrdnOhik0ci2tp1RUf+8bcxDuschIFCUiM9DtJmOMciWoIiFcDCkP6s7fdH4sJKI9UKYzE
dUWeBi3QrWfzRapm2197nCiPfUa5GS/DDEf7jleaVmp8M8S9yukPWS9ezKrdyuc3qaAM/6krB9hF
huDRlrg+oLj4JRwPd/bMwTxgcZsDe62oNHdkBnnhw2l+8/eO9MglZ1VZgRFhQHtkoUKrCifh4Kvd
Qxpjgi3BKbMasbsqaf00jdBDcb+MIJA2rJTcjPipeNK8DqMI7Dqi8B5igstWRa0WIgaeraAOC68m
aMISJX6GFxl6ytxTpqVhZtJPerakvS0HvyiSuqrWuXpiSy5ukJ9Er/TrKWBKIz7n+I2NDn+fO+km
sNWehBAJEul59vaZ5iJHRDtTuLXXCWNL4Qqf5rDHAW86C7XH0BOScgV6SqP+0zF703oEhHKIfr7c
uckw4U0GYwunw6Q5KFeNuU4YvNbrSlnnd8yUuw2XcqtbXB+Vpuw7YQ5rhECcT6NLZj327r0gWqJ2
YtrnuqAwYfBXqaVnvMWfKKlD6rtlj4WTk/E8mOH8gQX/J9t6Uz557wY6PS85tErSt6qE0dLdvG5r
Ns6dAxrIC4MtDvIvwFsMyrBSMoo9ETcMtTZgwI1rvB0LN8On3q5XFagw6owJxEuD9326wuI+ZzHt
HLvNkq8aCLQBKlZX3clRHD4xEOvlov3LdefAWHtcwMBXytNm5y6IxtKPlSv/9VfqvszPxYupdwS6
TTe1w2+nwhDmj8zakAEE2ikSyhMCtXRmg0aOtWN1pZOmkxdjEbW08kiubgoLXRg9rMTNrG+Caaac
CcxJPi1pCYlr9ME/l4lgdrQchNr50EZl0wzhhEiagxJkioHgAc1pNLcLwhbhhw9XDwd/D/t3kfXp
9pYzBiXZtVR9hsPenUcjOEqNvDnayPIBJJhq5TDLeNTlqhlHal+7UUwKGVP4PRtmHLEkZ2ZZcLqg
3C4Ivcz8GirMwFTCDMzulkaaB1JSycZ5ar4YTY6Lm4cskKtG26EQxEm93/kWusBpDb8aJQuLLaEY
ja0B0eZg3FANpOI8Dd9Xj7mS5YCVc1Fg/tKujVBEMBOmx1UG3M2h9NuML7Kxq/nJ9alxfdSLDPqd
xX3n3LNZCWtuOHGbo1h3OGW3dRmTGVPtQYZTnrO76C/LVUXSziSO07dNMv9a5i7zhW4aKFswJbYa
GjC7kQs2hHu313pdBRDuik/DE0YE5F6rpGH+Q30XvfLOExqBpbC6AN7Yq1LXhgpDpkZ2bRuISRhw
uY5ibC6R2y/uT0T/3QgYu4bYqQF52BVX33pB/5KDcMODg2VnfSisCnszPaLBObwFcDEnamF6k4lZ
GdMGawEkOBwk8cTHvxgEgdonH6js4Tf99RuQS13BbmnzvoMNA2GGNlIKALLAhc4V3zDbamYbBZo6
8CVmJ3NaLtpnzcp6akYgQD/Hapv++n2x90plg+n66lXjYcXog9elIXHwoZirASahLiL5nZjGns4b
/pemB2+pKWW/ZxK6TeYBvJpMoS2kP08m2/OZ4nQrrU3Gh8aqO8UDOlgUEYWKyJBRouBR8shkLWmM
yN7EwoTP3bIll7f94hWTNksAicIDZ2P6laNIClGOMmf56rNGOfo+ozXbxglNfWFywhdGXxL5Lgx1
NI1J2WN6iZije5kjNpqVdqYQKQ1zC96e3NZuu99RLHdxj0D0TobLU9Llq9HHtDkL5QOZ4JYghsni
qvNgYDCO4ns6PQFyHxsL7CIkx09/jCASLoFWGtvaHu+Hqw+DBYchYvGph0WwDFr+dVKcZWIoj803
84KEk3GKFE4iOX0Awjs7LGJgB4bfvZInIelwFTWNBecEGl1nZcxJe0ynqTrO/uu8MlzxFj852fhb
ge08DXUtnVhYfILPTcZ2ahD5I7sRkvp/OnfV9HJhbQqR4qC28tHRPbfAQIH1tKv8hFydvHJFLMjS
i8wrX4V4RBakUMb/0mrCJYpRbEg/biFw70QVjGZESLPxnrG8z5YLF3fhTC2IpaxNp6zbVhR2QVRz
HoF9j6M5w9CjoHsuupQjU7MpVjCgEobh4JRKTwyI3AlCp+nNKc+7Sc2uaBhE+oz5j2VnLxwNrs7U
aSYZ4N/yptghi7ZfrLZNtwFtknoPO/I03C5EBDI5BsbZdz8v/Hzg6XWf1x5mMXI1l9+0KZN23KPl
aIx7RvmOXe32kLXZAfhjdA4uAwOPh2LIFrHGj4Czf7EiM6gZaZQ/IkHCL0iu14LnG9IHMDuzI9Lx
YrqlxPU1I306KEN7xq0q26N8LTfh4Y2ztYhvf2ikCMxdObLLs71S+uWtqc0B6awv0NlSFOLf0jBr
Hw+ruEm4lEtcjncEKh5k1hKp0v7exfTjrE+Ah63FdSfOKw+5L26PNNGHWyynTxHasNLc1qPKsQSo
ou8UyI0AFg9DuFaosNZd2Bocp5NsALQaoR6T97xwEUobADFRPCXFD7QvODRFCGk0zirYTzrNebsp
DtqcemydRMTa7peOkDPz+2A3WAkh8kKiutfKK4bD9d1EgAxLjjhfMkor1Vk2cF4qSeDmoQxfmXyo
7GcaZF9u1KFQF4wGHkNpYc701VmhGl9Skgf1euiQxPCR/NZ8pWKi6tCbmMV6x7gDEPmBF3SoUjgs
DBOGcxP9z0WWY+oDn1J31CqbXBLEvoA5mwNh+CMP9O4ssw/CL9UGo2lnQ3cCi0fy81pP8d0ZCxGJ
G8IRjff5hJ80NcuO693bvAPI1u+nIWia4R6hq+Cf19Uj7TWO2oAHzgfQ1ol+VxomJc8aNe5yQph2
znUKGPmhwX55WAfD6eYskC3l5tyJ6M5JpGQAyCKHYmhli6crgpUdNBJ2bMbuNZ6WAMcJtSlTRNXj
DHlUrPCAUlUN9J9X0Rayk5AelNWjXFMEYh3bNYuO3KjMvpR8rIp7OMe/HGPJq236B1BEU6pMbjOy
tffKHsqEQVRQ3ZvrJUtDHe7v0mO+0xdFyuMZBxCIbs3iYkVPvCo84M8pF8na6EBoyhj80MdJ14PK
I/lKrc9H3OAjp8prVfOo2PxOXKtC42jD9k/+7CBOm76uHnk/QtXW8p0GtR37eHeAB5tFqJWifTQq
qjHv7uPj8HenyjpQ3kiwiLUaHLOPeCPBbi0UQSuQURKd6hzwwEmVcjOgK9lU0GSlUylMJ0Lzo+qu
EOQFv+b1xU7mGjVDx8zXxau9VvsPgOEVL0NTGrpd5HCCR5fkb6aN5/WKK1LDh/uUAhS2nGub/y55
FyVWIwy/PFpxe40tOhAqNT0FSB81lG/KsDGX4BjxIIdAg0iXLAWFxjymOWpQjo8pcuyPtaIdT7QI
FTK08sm0rZoth8gccDNKD5rPBRIZZ9yjU47rTdSSMf05oeLV1EUYWMo87Jw6U+eij2Rk8kZHVVhP
zuNUxoWnTLMLm408+diph8nYofp3fB6xTbUZrXl7GReWjA2vuo5pG0Abd/8v+/A6UBr2eWSe9Mas
jVZoxXLcGn8x6AQSr1oz0LGlhr2kTQo15QETHAvI/lbHn9u95BKGuKWjjMjNn3hhilffMHFe7Pkh
voMGveGQX8CbZfKJksac1N0pw0kZKErowRFUL5O3/fDMrlJkhR9UfaCofgW7N+o0qYbpWAQ4JH8V
YalhFznAU1to/UtITtxFEB/mXFqW6wT68TE0+4/ZFm7SVU4nOzVj+kJBLIEaRHeu3iXE/x1CZBF4
Cjqcukhu1Tm3WvgUMNhd8sj5NWxEXnTr1i4BTwORVf/dKPyzamthbDKCLiocSb8hcdn8dX7F73CT
fjoEGgOqi/Ip9JGkGYJQpzLaOaRmZOJa0K8Nib0Df81lftqS3anncU+qnM4G5hCdbiou+Lg35f70
UJbuJoPY1jA0YTYsNgk8J/2nhahWFe5jBwvYyEDNM3o1spfQ7FtSL9mERB3dZI33rCtCnpu42e1C
CqsEigCufeTGEjxzsBTnRXMPsMyWZ3n7O6xB8cLNvRanLpPCE3AVuSWu8aeWf0A5NpUGpQC3X8mD
IHmXEcLsB5+FODcZlsipNjMqdoynXO6sPI+D6Gs9LDouJ/6Q4knoa1YwqZ9ufwK4sWsJGAecUv9F
HUr7CZdETTM7OFmAwE9bdLH6BDROI5V/cOCMKEJsz2CjIzXVSZP2bYTAh8kBWaLhAOZDQkNNz39o
Lyxb+kqIDvTxAlvjDOXMJKmUfpCHDTn3d6tG6g/ay3qMR1wEsOVQxRG8JXn1q+cALhgDTPX6olUz
cEeejlUfCfCBbaDSj7aRBRtkVO+NA46psdiNK+Dg1A+hOGfebyTo0vkQF76Z9eW+7RsSXVSBjcNY
NYtM1NSQJrUV8Lz2oDamH2crRneWugpV/bGmp/z0k7j5F+zZIMxc+7TnRD09DdtFn56chToM9ay3
TBoZh1tGilwcCaCNzaP4sv7xZTLZSu5ACNjNaMVmYMgzK0G242rZJTieWVFfwMKRQS+ITQlBamm4
Pazu5u4nTAPPsDMQm3qmFg05J0v6EOW2eQi4QX0E/URJ8BPt7K9nU7lGbfNstNQqBYXtP9FRhyID
0//8s4GfLTefvsN/OKMn0msnuCUCnCUCmAkZEhOfqdpEjuTHV8KXDlAFm28zAYr/mmpEcQI0PUD2
t6Q/XNu8K0NjA4EWdFJMam08UGwCSapoBqkVATX6FWjcnWCTdH1HgO4IgFPDGzQA63ClDnDB2UuF
7RdYF2CbMcudM+c4GRMNuVI7TCt7SneN3Ep+1Sg9r08qc9gCihqUIr1Ypy/9puNoQFQDQ1qfIH0o
qT6GR7vTR1Omcb87EYscVs9IA0wCrN5U6Vysn0bp0OsKg2bSVQYb4Y9kllWvFpXbPxCa67jyAv+r
i+SeuiPFjzF/Qp7v96wI22ErYmEYGX1n0ZS5qcrnC1x/KvSA4uIES1q/DbtdrhVJUoRvrR1ekBEK
bTM69IdIWTeUYiAt3CVOb2Tjxpckh5meDMyRCq5bec+Jf+TB4O3D0a8zjVEmtKWFgzrXDHWdqwgk
xRPJptudovESNIaY6UbZMiZm+4hvKT/RjdPtLDPMwfLcgP7kpR4zlWNd839auIa3gmZHf5FSCJ56
o5lSyg0ZEIugkMLzUwJdRzCJzUG1OkOjIsM+FExwRCbBpO6fdZRI/4Ei8M/fAgODfsrLH2mWaAYH
6FXC7Kj0JXcciDVgLZFBcHWyGSkfM8iPVq1qODObDaibQCY8NSOascaPN6QwKjTqbv95K7BYP2HK
88Y/G7ZazqYJBVJtw1burG0ygX+Q9fVRjPSH5HOhWo6Tw6gNly7W7z/WgPsfxuCESmucgPPQfTpZ
UFnlBsxyR0LVrgO07galvnFA2YpvPphx59g/cG0TeAaYSUQHfIhWCDnE5jzxjt46BEtlNu/0cMWi
t3dYGLbVin768iZciOLIpMZZO0hmyFdunAkTm+rqGwJ//w1cgrhkqJ+7x1OoS00VzaU0cCxRi4g9
eQ94mSSE9hHdGK5nNSwPFImW19AiDpC3US6pGa49ZNZb68AqKe02zIQg9ktZF97L7rVFyUtvEbyt
BMyC+Hr75IJYqk6MveRey7r8iDr/VvAF9IdFM0YmTRSI+TojRTm+gnctRJwDI/eglrcMTSA9gjtW
c9cbZAtXJl8E0x3mSJAAT28M1xQ49V/MmC/5B/CY0asjPTdQzQP+yAwis/5FiDtpFTZBWlLnbu8H
MBkBKi73y8Xq8LK7P83Kwdd1BzS4wTg4+ozcxxWYyH0lN/tuBMz0ioFgxyphQLv35AkgGSRtrtIj
iN62ifR7kNb3bq8RtJ1A78DvtTAuMPRoMYsY+ynoDU4tdb7MyBvCaZPmmTEPbOv1iGx4MEV/WwoP
M0xUetW7Czfmh1oJHpHWiPkFgP0kOX5WnBaoeSAyBAUoIy3iJ/Ja/6GSOnFeyapQ+xYg1ZMMDoqG
ZrXQOady3oXUD9c2XEiZkgJ16pHmziVo+ZvmhZzftmIUK9gW1iCC2zYSxbJCupM9Org4mQMRINM3
tE31BAiYXQvBaWl5oTxoX0ovnbrHtIGrcyQW6tl7s1gJoiMsMzYq9iUnOhEQAf6dIfj81uE/ztDu
6NbH6RBqQ16fhpGilsUo2ARWE4nt+WQw6Eb4w26zQTdYj2Yt5PWWf+TjB3A3R6LOnDCdL9b7DYOb
JpE4z/xHxn3KLli1Ei365bS4Lpl5Xbg1XxPPmQJKmJFrMDhjLSYxYjKGjucCthpid2eLJlNDFJHa
D2455qNwhr+qSn1vqKXvCG+LNwRlWEMbE9EQF56olBZJbnA/aLjX+9WNcQFCirpxd0CKRrIWhRjg
cXqiZjakuw/4krbS7eb69jdEGUAy0IuWjBiGfqHax1pTTOQjZZpXU9/TQ9pinXWDcDpvk5SSPAXG
ljkTiZSOA+bJxA/Hg+KDhqvO7UCSoiob+bOLWqBOE1K410+6rDq39yVao5AxtC5JT3cO4jyaXVJy
oW8cg51zqkqLCXLO3XDn94helU9HS3FLYJ7kNdx9BwFxwM9LibaF6pP69DPb0YbIGl2DJv/5vywW
7OU/WWe0CGITCrhh8j5zZuwngSywHUcI/17VsxgDV7zMTeNE/dkyQPdzFEF1ZNU/WLYeFICDpx4a
fUvrblnqszN1DSEW1NBRMCpvxE5CgIrMLP+yekVctfrzI53sq/T7fJVLurEAaorgwtFEHhE2RtGM
xXwgK6HECV/KYqY24DvqwbZov+3c+HpCf+Wq+5YjWuUxOFAvswyUePUKqd+2JdG/vbCNLwfPGRon
HaT8Vg/dKhET7hGfevheZeUOJUsUMcOHCRyaAvIrxQZtGhiu4IAwKxsbjXMvRARkloKZCfuWZPR0
McPB+dGvSpwjgX8bXb96px/0SAjN6WWRA/YBjS3zkdQYRJgkFAZTlazDahLBkGncOogv1H0EW6sX
ZfsHn0Vy0yIO2b/pxNV7FSUnSMH5uw5rw2xyhftI/bfR2soMjKmbiNpDdlj4FL5Gt8WBWcfOWQrW
houBdd3MNc89IcgahFtohb9Vu4fd10b2YuTP6e6wV3A+ivASReH42yMSkUMitoW8nr4i4RpHLenh
e1NaUqx7XecMbvriHGELH2dz3yH3ttpchyNzzJsATDPxPWnKEdcVXwtn+TydbcQKjNDokbzLeYqr
uXO6SZeVyMC0cY2vbfeXYWhnKEz18UyTZZxKFp/ch0MI1Dmf3ahLcCFN2gl9c5Zz2h3oFMpNykRY
vCfl1oQ5sjOMc1x6lGIVf7LzV0QOpGyoviigyE+tyQDQa8/ny/P240O23OFjDw2/qq+bhoBwYW5w
NiuiW9rlL+b0GDvYCtVhqt0ZQXuh5caK3+SM/Nj5/1Oiv/OJ9sI84K/BGT3gByQDlS328I7Tc6Ew
f9UGikJcAxCJvNojtgm14VicY+fyDIUW49AgIUZ0/4zkz36vWVkZmQYposf700UJtn9x61vfNjf+
oOlRV62wXdtJK4hxLdiccCr6fKuyODiNdjYPiM6djNErfOCufTEykoDwnPCX31LuvweeyZgBLYLX
3GAtA/934iqkoLz8IsIFxy+O/6T5AaPibB06ESBihN5QpoNcSGnjdAQa3KfMTBK924G9YZpTKwrj
xD/sJxscl7r3u665EjkCPi+rf/jk5pSXZpUiIY5ke49RwLb/IabKJ1XGgXkGlWniukgIReapJmN8
oIhRqIus2X8IUuVRYKR9WnXYZcEGwA9j3cPKEhUXzOlUIJsSKkIloa93oFzE/KbtsXlSfGGL3a+A
h8/1Yq6bxw/gb85IWc7vKXYhFxVPWC8k4k5djkLZAnct/5C3mApwhDq36RsaIENw6HiU8vLaK0eH
1ekwpMprnKijHnryUuHCwzB00Cc7ACW5yupMXtl/d+CUKl/+0fkEaj4ErCHtiI3ud4D4KnCCYcQe
+4phEGcm3YoIjkNcVKTwg3kGS1F1a9RXrZDrQqlozSk+JoMs0mMvduhe0wnWRbYmx9a3/F0kWnmq
jhizGD8IY1U4cpzpPc470Zak/ZTpybQzo+67OQH11zqrwt8JNdolCIQ98xbGsE1UCNae9tBcjfDq
ONGRde77nmZvOFDlcIXSU4LV/DAhSw8h+bUYQaNpyVZUakTrC1AlND3+L+OVEhKoFieyWpsgRZYO
ge52ujgFx8fgJ+WMnVk9ufEBCsacVRFzJ1u6DQaLZITPZ/Co9ARHJVvruBCIWrSogKp8m+LE97tW
Knru4ba1k1OdHnR0Amyt9wDj+HWvOLW8E9bqzIUvHpY2G6QDDUWmfQS1bRoW7KFFXjCFHd/tTELa
+HttMRM5zvwScsErJ2e9lfB/V+RQOS0oSQncU7asttM+wpZuVxrJt9xUgE6BajHGzKwgMqQkPZX4
lR//3TU4RiHVunkAb5iZ0Vt6MYibH15pyaAW6kZMn+xfEvTNjNhrV4UFe4xuT+hyywYd/tN5R0Vo
kTgk6Ohg7gF7jxwTrK2mxRfgLZH+pALOcry9y2SQoCrTukMDe6uOEigdJyFYxAIS4rw+HwZQu9nw
maoP+hwBhTES8dKL3Ed4FaHZ7RWXv5C8QIzTyVMguKGKjWhTnOqGcWRdfsY/gx+i4p56BPqQVDc+
KdZDmB9biB9W4vvY9xJtf+xj+1kXw3MIlH63Ksae6KF8KkQRP2w+5n+nL9MVuve2ZDBeG4Cbijpy
gUiFdWrh0B8VhM1AGwis7nXS73F9ovCsWVi/g3IrwuFd8ohz/jxAxE+NomVL04vRo4hhgTr4qxuZ
NgpKcXd19x1+WSPadOd8jev5Y4huc5hFOrG88+1/Gkug0Pr49c0LMI+bQh9X2SIEUx0LR+VNY1fC
p0ksg0TZCVcKrr3TTBlN/EMVjk1rRRKsAWIiD9c6jmebCqWkjoplgGsujfCT7l5jiCsSTgDh2Vgk
HY3+1DcKaTbq1lMixYEGrxOKENAdf+mgJjwdzZ+J4cvOCgqAKXAg9neZ7K0veIA8uYc8N3svAZ4m
CO4haBmx4ZRtSd5kaS1VOWogLt847s3Km1+aC730a43K0ln/eysVijKoBd+b6KCicg+3iOrD/Bxi
sd9CTG4lapYHAn/P0seK/8CKHRgDFMZ6APZ8mxZbZYmqyZDPBTCHhuEqO1nSIwU0rHqlPy1J/SU7
PjSO2HL7ldHS3n07hEevatVM+fcbj5IhTwZD9PtMIehkaqbljS3//++NpIezIT0jtb6sYb1AmJ8W
76czF/mQKKqv/TlPaF9Cd9O+Dt9CeuAkYJ8kH6+ysyNNagBOwk3tOsCsyudD4nTKc/DTh3kICtR8
e2jU4IE2EmAG8bOiPbNb0wydNGoi6hHIShNZOQM9JtofW/inJMCe+1BSAgzSh8d+JcP5i/7h6TLZ
7ArfGr6uKNLV/6fubVxNeR3c9wZY8N02x0cyaN5NZqIWBnEBcizbq2ocruSiFo75BFxH++OcQ2fj
+lBDMDKkcKRP+/5KOq3cW9Rh+OrIGo5abrXR4b69f0ZVDa7gDxcJzmEFV8cc1iwHC1mKa1+hb91U
Ci2N7UXXBGGrc4wZk7hhalPo15GYxjLyXzJQO/+8MHEU+XjaMgvopiVveLdOvnObgUjZUQ0HZZIG
Kf0Z4ZeWyE9vyDRnhyjnD7/5Ohrou1sGd66wvTXT7MTJ6wpluGrL5rRrQWZUXZgsUW9wlyrQ5Hn0
SYOvlkmB7LaRmu4YLLhfJTP7VonakuQTcYQLGHqh3YoWw+qm7PEVpQOeBTpQdZD+N1Cgma5DeWtx
IY0wwdDVNZukeWEal+5ieVEgKfhlHaQ086hEd7a5FBYW/10uHa7Qqq9KhqgeTgtf1g3K5zp4bVz5
pHE8XPj2dnb44WlkDlXlSwY4aSHqojb799uBT88cdEK2cQOo67E2cys1AYXGMS5Pe/eqYrLTJF2B
9mMtaQWtP0PuIYOMAr+TKVqh4x/l/XHapAKbdvkKYsIMoEK8cjnL0bmto2GffoIFrOekY87jp6ms
RaBKukBW3Fo3MhGFwgK8le5CDeoysuOpfiGCCO9u8NxCoc8Z6O8ZOVkNVMGkTPu8XBUHXfJtd/R4
2cln1QuCgMfDFGqRfSmkR5WTiC2uKCaPdkriILoxmPIfONfpCn24RO93tBNMBR6IF45p90W6PAyG
QNDmjvTI3Mo1jnZhsOCeWSOO9e6MDgGoxafuHD7unZTyOfrIcyoA2YVI/VIaMMjYpf6FTE2kVScN
XGlc0G63brX0mWJmoVD0f0lxmYkaujuLFznS9gFzJdNNtxfVQbtIbdUfRF0kKvOXL1+UkU8F2fc9
GziaC593iakQmBNhRUyygUECv06Mt+GxpgqTjF4JFtUyL5dwFGThPDBT5L6JHrnbGrZqdIXDqpxu
i3fNLXuDhVrt+jzQ4tqKWaK+VQFJN28oKcgDplwZtrr746x562A3AuaJl4E1IzuQYu2/UXEvCiXe
OQIyw6gp/d6B7VPoAFnbeMOiBjH5nenmXXqaVlU3XwPSCEtaOwO8OeB7zT4sPjM4MQaKwL5w/65p
DwhOJusUqpOLCIkY2x+iruHKelDu9jdJMM3geFRxiTo3MeBsW8gzd4xKo5uRQ3X9w7wF6L7TAtwx
N5xG2qWMwWYhlopId2/JMmtKF9p1cDZTHpbmxo4Vrbwbm7H7OOwLOEexuSxBw7R/RM0jdA2bI9C8
mTkOHcf2cGtPbbzREKGFpEz56gdbdi7RjnIq2PNpBB0TMsh0YCPhtW1TQobJm7Gy81aQ3OMxtIHT
+rEU6+CwC9jtzQkVyqdtqgIP5BiawZJ7A7ulcP75K9HvZN6LIxW0gSsuQNE64HGGkpG1o6pRKRmX
5RgFGhORGl4H5r9sBsUBz5ZnmXA7zqW/oGn+3011VfPOlPhgeYaWkVm4+j3NtvOWriusKD/LXz0R
8itTxw7120YePQ5svSP4L5YIlaL4aAp3i/I5Kg1iRpEh6J6XERvfVqE5SFAVDzFwyb7UF8j9Eq6U
cBMMtxjKkTbxrP/gBbqOAMTdzgp7i2LdTf0IAyeeDpyyZgcrxzog/yjHJ1rPgV71CNwV3YKs8smT
lDQ1wPJGTom3iZM8ZoutdSolwCwokL5eQmiWd4kR7sNHzrsFp6/VQGx/PS2ITXQ0X3d+luRS1S1t
3/nn6NRpROPqrD7lCEzowqbeBrMM4vqbThXemmqrkFiBhXaeQF8qCY9wUiAvL66GVl/yws373HDo
I4wqmRgqh4Dr+1HzPRqfDRw173B2DcrHiH+XDT1zVu/pIi1b7m0g8q6ANX86yCdOdChMbKr42iyW
H2ll+aFmXSEgX2Ut30Tt/KloL/sxgAROhdHB7uNbB5CicJRP0floLLu0UshkXMpU1WRe+tKEij7o
g/ItRzW422mauLfeySRpCUuoyIonJiMzfjbV1kslludpR1obloY1I86HSMcq4KXHFCWpWVNNw1N+
XREwcOBe8rUbh52LFqw2w20Q1arT1He4tQW4SLi8gBTDXzhonSQIEeUkYBlhju0oomFMT+PkAogf
pGs/nlRDQZb3u9ZcFy+9qey25sweGz3WPAxd3cFYsEnQmvqANiAoWX5aAwUwCgTh8oQ0udNjFSMT
N9ex/3GbiXK0v7lMnguwbC06keIYJMJRZLjVaVGyD0Ufmannx1pih1zmBGzlJbdsIz9vBw2bEziN
pXaWoZCg1lRZyExS1FCrK+pUqdAUY8z5cY3PscxdKZjXg0EFQ3eZ5wjMEokOJlDu2GJPV2gWG7ac
PbNcRR2lGgjc1sNgajJF/Rf/gt5BhZvHpnlRo8ALXbQwSHx3sOkRm8URGIgcmyEPGRG6c6p3bbTE
2QA3lZvEsxTNDUaDSfnbNcoXafF86LA9aP34ZI5YQOSrg0VrCSEXFXpaWpH7277/H3i9ebZwOZcq
jSDBco2tBFtLXOsnItRzFxiwqEHoupidvBlcSDiajhIWqKDKKDiRccMfnDo8472/efxoVMA52qKa
4HcozSgqzhhbZZwzX2aYDBTelO2rcOry2fIKpDkMlgnmZkGQO8DdotM9YtHPNp5DVK/1GUquhxgQ
pQh8zpRklyN7HROHOf+rohKIprtOue5i/ObASF/hj2v+PM7OBYW7z/hqZaSfqa7KMXpc/K1E2mg1
0NxUQUZZrlMvFdAshqTLAmMZ8sh7ie5pNjbOvGpivHXYboro/wxm2LY4ZwBFQElcmGrqUqn7SnhZ
pi2gYWpmTlQXbRU1liQ4jPC0B19kygy8E7Rh5UIf6E/TD1RFkraf1WV9++EJeJTR8INhojeVCuQ+
IUoXiNU4Q1FGrGAk8iPZYy2CUsV8WKSWryV52UK/q/E49v0VX1sgTRWrU9EExxsB9S50AhST38yc
4hOeWeZhLdBL0YmTzljsUG0YmIRkux9NmTuPhwnUHIy+x3pNxXJs3sYIFo9Yq0sB1CHPjAYCodad
1caNUSw7MewAPJeToDq/n6zkTZsPo5TSe+bUjk8Hxlb9IbVQHidZl8XW540LliUQ1BFKCH5HDi5L
rRVNyQUE06eb4LRtonFcAs06818c5DoA3Tw+m/8o/Zc5vxMXk0Rfo+aSL6FH6wmhgB3tIhcPMNJS
+a7tKVvzDz/m/j/+W17eCBed1u57MCn0vbBEX974B5Xut3Q0r+WjD1m4svm+yXRDMmaWzzIvr/un
mg9ZSFCat6N7m1hru1Mx+7OVi6QkI7X0xfvEh/UmGvT1qN/JBy8uCci3Nc8R4+a7qnA+ZMefDh+F
D3gg2pcxS71JlX375uUy2OuqNDwv/HvV9eg2ft/Uosb0M8x+0XjVrRSbrOt0rWV/a0Q8nKZPFSrT
LclK5WGOd747ezDtiqXb9VQa9AfMhDI2rv1cGFBPBYv6XySWJFzQnVopFHKULx/Xj/zPzRvK0ecY
ruWYZjxA+mPX+hsOgkBLi/P+BydYKyDJfWnZpOGCZb96coEkOt+Er7h/wTRc6piAh54N//eLBxl7
EEv70Mi0qdGVq1mhP1IPeWi519fIajA510kMEGJ31VQ+SE47V0j2i43lTJZmSoKHrMxEWOwIa5gn
39dUMm7vrW6U9t7XC+olVFkhacyKbY7rFC9OPuLMdpk73Sextlc5NoKX4uPHFint3dz3tnlrj6l4
Z791x13hxuBxHqqUhS1+LEn562zirEOcSs0ejkP/nldecd4FKhakeGcWw3m+TGiTkuzs0OmFHTen
8QEwW7T4pOymlGXRgg6WRaIn5Nf2aqqpw7IMEq722G9uuHsW/t5JthfFesxutlAPV8Y24YQyXV9b
DS4J3g3RJUIdWhNIat4SDiJH3sIzY394+E3z8KdVPZtt7Z3o3eECJsF2CUZBSIHsA0uNYkF9NaQf
CJ/xNLpDsUCW1iVP92VZe/mqmW2xyFi9wYOLmBJ5gSKaYhcZ1i3WZBREpHmvJUkvndv2kvuRHqMu
hc/VFyZHdiZVoYyvAjvdQsIQX1/a1dlZcE3laybFW7kt9pQmHvtZrriJvQzFmrUj0+sYfoipAFyi
Xvcsp8LYFKZYxdwdBmPyXGnHxZ7RbkzEjdQ5+hAPonX500WOXRfxV/nggFdRFUJ+itagT5AzobpN
vxCZrmhZTlehOu3XusGtiL2xR0sLiQdo94HaJkXoCf2ONl6LPMAyuJ6Ox2PraDjN6+QxpKnS9C3K
t5xzlZZHFt6WdqvXHo5lmzILW5efgAaQrmHkWtL8KDgkWR3Sjs8zJ6ZN+zWKHQTcAoHE+XVa6eTB
g9e8hNmNPRX8Q//MHFH+AOf2o/5v+/GHjkNZ281sDXT4Va2YCSnArDravgU7ZwFM3QPi/tp1LHOa
Wy9HQ8F3DoY515pRtXujrsdv8MNMtmzOUY3N/yu9u+VjUfr+Ahe2TWSE/TMAEp90SvVAl/3aj6ak
I/qqoaRUYTw9sAT/UD3JoA4yjyRyHbgzGjyHPm800NTITRpydwWCCrQGy3IoV+hVGixe3G1V7k8s
ZDKnut8cS7UrIHbWGkmY/F+1dxh7nVPFuJObnKOijFXrE1NpZVsR6MSlMwTc6K2L5/CLHYvLNb+Y
989OPpajrVNcga0aPcIwCXm8e9tMRp21mwgXUuSR5nuY7cpNP9JSxCvVKlSqGMAWosuMDCbQtDiY
1S9Kul+7HbP6GzPuW2sXo+MeQFJ1+F9qB9NKPcUPXDvhDdli2k3Ln5/wq4fwXDxswpAGZrC70eFk
ea+RMyfGSld6yFk7XqjG2G1vU+kPqYUbodhFGJEcOQfWjyE8pHu2T+YG1NY2iMXEZWLn/+/D0GVX
o20EAUjeoM7y54+4swP39GngL059kJKocx01fOdNb+frhIo5H5Nz/b2m2vU1NxEjVEJmOkj/PHcP
Tz+zJXOP2ajGd3dtbHvROCeQD1vyOhv3j4FsMDaKq/oqPJCXbgaBD0DXAQn0alTP/GO7MRRPEL+M
OOaVsQWiIWSGxMRhm66dvT6oJyJHzorDLeRek98UVAF/+QacuDB4qIy6nfefGjtIHJWli1HDkCsf
CHi0IC7N0nnXPDNXuWi/mhHz+JJJQWgmH1enxV/AlxUE+EUJ7XZU7RXX84hqw81URuax397oenWw
PDj1XGzPtji2BtjOgSoS96xjThpcO3vwOenVtGYzyRMM6EmlgZ3AHGfwI/RY8C+h3XMR0jJm3sKZ
f8M0chpT6HfFr6duYb3ZKliDLsFJl6O2lLjvqyPhjEI7SEsqmAPWcue0QHyUtFt8TK8TSh73HY9G
YmIT8Gp/B9tZEEdO9aa2kK/Lt1mN00g3F7bbiCV2Lox87rnXeqwG1VVcx3z6sTUsSXHGX0QMn7zC
hz0Hj8HMUjbkQiHuYT62B0u0Kt+oIpJ8CceSODQXgCQ790Sue+zhHSwjH/cYAuaJkJPBWCPMrhB+
kG/C5gfd47mlVgzNaSWuUgqwdowKuClcfsY2bLC/NcmhWFNTrk/GVNOzYDi6mZSwKlK9Vqa6+Wa/
Lu4SAnDxnIasPcWfLJO0s0sDeW8JmERIgi4doPLsY6pXKhe0n3mwBw71f6G6aTLF8RtMixQIenAk
GCZiI/cgxlYdikV5yZnhWfFeZlEoSJ92QppaMeM1Ae76r5/NbyoScLLetxqJp6AixbJT8ISkyHfu
PdnuEXgjP51iluNQTrIf1M5ivmVHa7HsompGezmzqxd7ttRX8hQibNja9DX8in8o07ecMrlJZsVx
aOB1+hFAipnAHbT/xcIwdYa9goWzcX7ct3XROtETVG3lBDKHJa50b4aQZS8hNZUAGVcnzvu6ks4O
x3CNAdGDMKY1OWFczPLl2CvmS43a6x712powC8LP0gAkjo2pDM1dwWUhJTLB8VrsDnG/B/c3T/VF
mShZOkXS85xWStohCMSgu+/gZehQK/ZiZKxwoAL6PH6PBALCwFGdgJN59MowrS3E8ROS7osoMDqc
pSvhLcZTfJmnqgmp55tjh64ewengqC37uwNS/VRKlP6h5ZPnsrvOGeo/RTmNNblUxMiG5A/6tmTw
95D3GZR1q1B166ZeDTW+wY5kbi6aHVpBeG+fBRO1Usgq1t0XayxAyK40X9nLmrkbSWWOwDKBvoQT
26n56f4Y6857criKgj2AM2s88QlVDZUV1l0prJPs2Y+D/kb51aljVMWho5fJ6iUbOnlpfomzbpLk
R1iiY/5lyuvquVx5fknyDWteJMuHgZoCSjwJ5J4U2ITeiORRdx9VKLzS+1C475vfetamQw0MiCjn
ivat2pBjEBXmqZlZ5XnIxHgiz5Dka2OGRQvwFWLZh9Tcd5WgQMRvtJtDcq6ZY+CKMsZGu49Wd5Ny
2Htw8O7TLyw8XI1fdvK23CtVdM6lRysTu0W7LHAo/6GP5j6KFIBug0n/JJD8JMuQLZvi7fE5aHg8
8ru3V7phChvtDpqEFVA26386SShsC22PNWBkUeHqvt2LqSilHTgSRGxQ4AOhXWls3fc7taikVzjV
jH4tpO9kNOm2GvhnlTrl52M9cSj8xMzbU5hgtohRSHTWXKJOl8Br+z+th3NeSQZ70LenuiWDW/jU
2Yuezep53E7XH5anIu60xpXmbSsKjW4SPa1BA+/m2A/+4o3zF9L9DSzpF+II6OuGVx7bl0tkVjvW
aERSDEIIS1h7v1zz6ENGIVbxlUsrmYhqVU55QWfPTojS8Gd/Fp4ImBbQG+hG7vEhGy8iH5TkwSiG
KjqWzRNl3B9TYrtPdm6b2qJs8APWnS5UPTeDOVAorSVT+FQkF/Eddn2NwThdynjnHsS8d23mFm2j
6T5ie2dj6ct3tnniaBiLXuwKuTCw5/pQ0Vm7plU312BS5cEAu3YWXt8UA7ZEi1OCOqp1ploxCjVf
U3x7Y8ktLYg5IPhCtiVerxtDokT3BpNfd1MW9fnUX0H91V8Z/8urlZCyVCYw5xbzmzcLLZLOdSd3
cbDOW8ztiFM2P1k4z7oKSuQF3pj0RclkBfiJPExaFjwSntcH0syWbuJHfU0YnqreVMI9ndG9i1R1
2pnh+5kTmbuztozoQpavDj2cW9+iLTlH21O8gqx9pWFxIwqOCeYPT/nOV0o9ApyPhP0x8Z5cdyQt
mHA6NU6TQLrTtQx+UeDXLO8p5GJLce27o1SGO1MAaf9L6umr+KIEVQ/FJ8hSYDDVG4Z/93cP9QwV
DvX+mHtU69JmlkqOga8poBVz15ApSTdM2fQk3ZW/v9YE6V0fEQgF9JWeiBod6E06YeNrBjIW2Bi6
5jlY42OrHkn6UH5uu0mdEYnE8Cbsa/1Tt9LzE15zQ63ieHXLla7yKwBaqC5XPEgvZqSad/mypkxt
P6m3yr8jIY7KtTYXqPFVtZFPaIORDPDYrNQSPe/XVS44Nyky4vPUk6uv+k3ExTRfufDk861qLXbf
Hic4INZkc4MoWRUmVe/+QzEEToKOD8dQaea7cdEWjsNhd21UciWDPZWqTul1qVqOS9KE0jaoBWVC
y0cCvoj1nLEWZZi7fL3UYkKqZmC/BazGg/AqLUUHqTox4obepk0WoqFQ9CFIUlO/I80WOAuUQs2b
+MmUlgQlUPuvbT/3Wm5HmUJqoKw/BHALiDQSQsiZGGGpr+Xsc3MwySqy20E0Vii1NEukhXBkXRY3
lHiVL7Mhz2V1S1vmi/nA8jtglnjnSG92jRAaaizlpZ5pu/sHjtPkUlG+VwisCmjo2yniNeM0gwP1
ZrnknkMs40lECVqJQ/RrezFbluP40XSoRE2Hb4x/CZZr2I/f+l+3KXTSFekYkFlsTYtRQaInLGOA
S7RwH8OtTKE9o79RtgaEddPfOn/mRrNJHs1YMzvYFwoK2Bv+VqSbxFVOzbgLYTECysQwWaQEh5E8
VEiPwO5bLvLi2QYOtf5qcoYUJTdkRtSxtYpvO7hVohOhK4+V+1M9glboekrfZ0QHyT81mIiC+dM9
IRcfghmjgCeU7EuCmV44quE60HgRN/9MWr0q5b/XpMcyitiSpulcYZowlHP+7q4QF4R83f4Y48R/
zW8ApsbGtvSmOxXiXiRod/3mKHZDgmj9ksflGX3gZJQkw/N0Ew21LCl3cc/EBdA9ekCWfs5hiTc7
LWH8xkbgrxTIxj6POvxCZxTRZwjcdhnUy7qT3zBfzA/HutlFBICcVMvVyO58ztuJGfJcIXE4GZfa
Z2ZGqoV9CflZ1MbrVzbSOmTC2zelkJXSRZvqJ2C8uNVSybI98p7m+9xzFp1hl6A4ksrgsqENUmbn
r67XPBzqctJxSa1Bwk102kIw9uqMMEJpsi3xQQ1FV6F9kBI0xkLaNV1TpIeJvAxXv5bP5HWzD9df
LTCUsMKKfeyrbniGyf07Fs7/zAyB5dqUTUXExrG+MIuirmJptRGAX2SY4wC+flSVzXAVNFELegmW
7zRlMxTrqhHVEc9jv3fde3rKoZc22d1Z7XZoO23ZwdpGv6x87wTkObe9+eDzuywyomaf6Jakb+ix
lwFYAh1nohO81+xm8HRvQy+ufVoDl5hOYkiUs8vKebKgnu6mlHCCmUJgE1AZgK6/6+dB5vp9u0fW
YIYqy6Q+B/ohsyECVYn14jrtFg1FOfiH8txwk+WgDG6biJTN7trCpn3uysjW17ioiQOaY/1nDFbe
VWihKRdzRIReXci2bHoXivDuMqBLus00fTZiMZP/EHBopcdcpCKeAnd2hhy7aYZGG8EgffmES56w
cvGK7B5Oms8B8SyJHMqv0JglT+rsgiXMGSfTB/R0LrLZZbGVyYpCnmVL/CJKXdEu2TvZIVNF5UwE
Roh4dE7alAtuQNpycZ1BudlqOCWkAUr+az+P9WOytMyP7yQlRvIhymeggNzRVH5bI3j2/Jt/iTum
vdiX1RLqxCdUXa086Y2RXQpXIfQmysFd/Nw6oH79ZpFALEUwXTc/tK7FFwxfynm5n6TeL5AEFB8Q
fe+Fp3/jhTQSMNxmPlulQh9+EYWRskLR3uOUYjRQFr8mdUdyAEHXhClDHC3ZRri6i6+GhzD+f+FQ
TDSAnZyfUieX8k9WL/Xu2uUpm/jLXaXlO9q3Qe5giWSdIjNiZchTeqz3JL81zo8X+xCa3THNDgin
sQwG/J7e5zD4q4AIs9z6QIWg9K9NhO8VjICmmNPZw4eW4Vka0VIHjgi1o9ZmlFhYlESyor/4d8F9
/gOZweGW0ASPHNcm+BYczEY+VAQeRND3otKwS0CWP3sdExbcV3euqX2UIK/1KQ3OGwLssry7Spv7
VcrLLa5bmhwhypwJTpPu/rwDo2+jwEkl96ixDFBXZL9Bek4mgoz5Y42bZnsYxi1oK4Xtbm73+GF5
bQfy30EjXWyKD3nDKQiWoqw5lNvgl/c0p78lxrOaK1Nlo3yGDAJvQeLj9YLGey1z0GieYqGL83Sl
CIVnl0Y/TLLNdhOv019rRjyns7zFyoCKE5vmM4Hj9CT4iqAeLw6vgnF9MsQrfDcz1+xDbdIIwpAP
PTNEJ7cMlsQW5JANH/hheUcq6XVGpmc+n6vEh/yh1dM0ZGYilUJ69HPIWMQ+uHDtHANn72lgGjRd
blG9puAWB0C+h3kF9uXASjM7L/bheZL3Zn7MJ14uR6vRegBm9X4i6w1LTvVENNTJNx1sl81xIYIt
HWM/aMBb5qtOSLJQ+hqa5Ta4S2OsOFqmYdKhpWQrPuvKs+IGqM1jCm8j+fjIVEr/+vEBAcosagMN
fm6Ogt+S3aLlI7yFNJHfLPU1SJtSCZV8RhCYaVjyidk5AqzyZqOO3tMqDQ3shu9adZyvH5QeiBtU
St7CwmBeOH9SejcSjBMIvmNuUXrTlLG8iIZ8GyKxVofQabEQ3K5rhONvcD/gqwAIzTg4b5TGxZce
3VbWMyRg/BnYqc94hBpdvaReLiBe516Ox2kK/GrD6cmsKPH+eOzM3J+FTbArAHdLsLvE56+0cls8
LD9itX88369oyCJtFVnoQ7jOY16reV9iZiQGiQfH3rv3+2kacY27CcX9e2fBRiIyAQjwaY+mJVPp
xtx9ZzoFOi3BxvEVKz3vpOzk7h9lfEKTfdxDks1KAB+1V5r2TVw1XaA/6HPr57GYix5x2cKmfbkE
03EBR/xM7zd5lr7NcvtUnhyNOZcxsxLgd1McVaex4NGTrP3FNM1Gcm50xAV9DDD6ECW3NXFCTy4a
4qdFC8mAK/PZP+sOuooVPyXTEPp4jOm8WqkPK2tWKjkixglplWdgwZ6eMAB/O+VzuvJqeq/KxjzE
2dyjn9ylLsC9y6blQJ64XFUMwZkDiubt3OjkYyal20Q4Jkp6LOKIvmtu2OT8dPCu51cuuiKU5ZJk
Yv+HtC5vvbMq5De5v5zNyBabvhR7SgDd2VkAnti7mr7nRBnRlDlqgXMZeaSCuzZIJdjeqdvQCXjh
pvjx7Lru1Mdov7N9wxKXc0fRozUcptPvRlFKbCm6ZACXfcLxCEZaNT8ZFjKEgicMMqPGMwsiJpNS
M7Rq/ABsDVdOHGBcsRmEPLLpRTOMcz/a6Pn6UEiTFaBUN3VDmSM1IyBpc8PnH3t+R7rabbfhVNyg
Wr6R83JR28WsUm9CPLjdkm1+7qncaqvrfufqt+YDjQyMJWmyKYsRvUmUWFGewKeDGkVGMJTfDOZx
AYot+l47w3BpdxaHyaU7gOCNe1t3SaEhuGPyf5litEl+tX8DQH7YAuVPBfb7jj6Z8YfZXb0N8/0s
c1Q0IO3R7N9+gb6ZAtQwKx5b6s2kW0fe5bi46rTehb1kh151I7gKJeh62cggjtYKK/ijfEqvatDD
Ev1tU5hxsl3mKCDid6Q1UdNbl6T92kSH3/dUYRIYqKz2qA49dCDDlESxqDnKnG0nj3dJOrnmGR65
5V/Xs5gb58T7V0Kp7d5t77LVEUMCdMK9CvJ3AbvzxIx6SmhXqj+sZ/S2YTjuTL9CYKMDfgfCjVfX
9K40VbaMxN+t5IMzpn04DkvZ0ThPhLnWccpzLr2GTn169ODG6iqH9ECv9Zc0D49R7hExkZ0dqOAt
0j4MnAydbYBdP/VrV92je3OdkBr7taWaZgsEQrgMtfo3vbCCJTLKAC9xxanjWpqHmR2ZdjvwmmMF
dagA5OF1qLjqLjrT4tqyVdFcyhLCUKaT8Pst9e1WhGcW2NTEIGtRfJlG1bwI+Rk+lGHQ6yVy6sw5
tVD85U5PG6L4kUsasdQ23PqrpGPlb4qY/p/iCiAHO4L3SQ1XSoAhu2m6akndZCK/UdgiajtGCyOX
KUeHargYaP4uDMeSKj23mjG6SRdKyLqAxfag03SoWzcrY3wW68qvEfLNg9jn6l0DO4gWCmQ5n254
R3Ov1chdTmeJ0CXcOw8tLnVJMoAZINP2ATVPZlvAlitZOK4eQsohHUAb4dnY0+nTsrY45/fYbfRY
duaIiT2GOXyOZXYLoYTqVWjRBgAwFi/epBqPdbAajLHZyPhZ6Ei2yuE2vElWFxin0geTdI9PBHfn
XfcV8Ktdi0dvVcMxySuAgVe/T7rWQqCV3nyj+YoGmKwOIonM8Piqaf/VZ0rHJ7TwMblo35MGHUH0
0j9UwhC3FXSQE4JkBAJ71rAcCrkmeqPhtDYpQjFNdK/vpkukplDKgqoM12P9JgAl9CIo5OD3R1Ho
7ki5O47+Kf44dhp6bxdXbt3jBvpHjGxDmrRXYbgfXoByKY1fx0FPSZPHqcQ4euhX2vWmJW2kV6tP
Q5tL7ZwfeNmzEVhkUhGYx1Ue4kSLFgOTT/J82Fz2XfvOGE06D0FkicVZdZEGwi0vmxSPGBgTZw5P
t/vCVAOwtkpsTrM/Z/fUw59o2Y8gnrWazWDrYtshk8aKMkY4P+83MigCAvbmVmwzZPgj3MhIbGbC
CuAnKnABkGmzcXi2S1XWo3yYdI9/IRwwUYj5t8okIRoGogzj8ugy5ygu3g9yiMbxyW1/GTtKseXM
VZq+Bo7XgyWnqE0147uNg0jluB4flfb6ibkyv1l7tuchOrHjb2aPN+n84AVRUtf0QVoU6aI1rlFU
OIA+KPkJe4C2F8+ITSBBn0O71e9bbiafAyNwyMShoXEqTsIZVh27jVOaquwmwQ5+zK7hveF1AEJi
Q/G7EZwPPuOTTvJM1vjtFvQJaPcklGBWXUBonQAF1y1PjhBTVleAY4D/nX4HVYW4XfKPZf9t2YKd
6PxrMctX4AByx/kizn10AzfMz+B6h8PDnkKNamBeDrTNnzbGUH6+40vZpQUe3/Yn6+iHvFzULZpb
+MHOxNZobctfi234d2+kShE8nbbqPLVZy6lwkL2nCH5PvMP0fXJFxF/SllMTPCs7bOwYZGJm2QjB
QhWiUsIx2BvS9KrIJstYUFMLx/DFh3Q91r8KqBoGyYH1y5Qlw1OaGkMpsmCij0w6QzcPU1q2Q7j2
wG+gwZZUIBeikSf64nqopiGH45ihaj7ozcsHDqERWmtEwesCIO0qoJI3uLUuZkCwpNJNrDQtiJDb
WIsHZjcuAjvDfMTbKyneR+MXFUI8XB7tjpR7uxETNg0zewwUR0sA6UG1+h8CGzjckrZhFQxlozRJ
7RMFlEFTogKA49MVHVzUj87NGPKMRM1sYjtlWdedW3Ic9pqUuIgB1iGnk4zVQlXnNw0NUIfrqW0E
S1DdR27IS9htbbwfV+5JORAgS9y3eRiC+IRnAEamd2biIjgKYD67CDbsH61RQp6msnawq7oQ4Z28
MNrH2LscKUj/m/tkDvT3QBE8VqZyi0dMza87s+D6PqbBzdkRAqJ0UgIl90gKq+yb84E7rA+zp/DN
daY9EwLTnMN4xrJSkj/4U3+Znr48W3gWkOBpvCqOAFs0vTIWO4xaFdThn7OV5XKYNMwu8KAIWmaH
Zq6jNpR7aAHGxu5Al+p31IF3xi1DaRk2PapX6RWl2O3UUQ15a/sIRM3QjBph0liliT5AnNhkwPeV
S0eFlkBbEIOpDW4UhbkIKI2PR84JayV4WzhHWB0FlIfot4CEHaWMa2Tu8Ei6pioScjFFjBCkaSYS
dcUVGN5XptyqyKahxZ0pp571LXhm+mpPGm3M+Uwj/+qG3c9sbd8pumiMKjzro1grMiY+E0vLhiuh
OmbYsh6RT044jfa1/RW4IvwpJk0fXF5cbKKQdmV9mHRMIG3nDrtNpv7ma9b3nMKYHfMdyZycQ/1x
XK6GMpRVZseF7eYvWJGTgFZaQGFx/kOj1NM/ZkoSpJ3oDSzO6ZY1TgGSYrVMdbL/a7PTy/gV1mng
xn/CqM58Qd2+dTObWVBqEXWQZCnE/Y1ndmX35nwRMS3ALxGivtDfJbhtcl5r45Eb49NuQGmLC5W0
hlbLFb8AwJOQq5VhhCLKUwuIJSpIk6DEW15eJJA+zpwDV4X36dMEhwx4Ek1wAcIPk8T9Z9Q5RcPd
SHku7guPKDJLQ2qaKxSTkVrDXBjd11eLNX7l3xWHJUnsVQgv0lRMA3QWmavzuHkRoPZBYJ1LP3B3
jK9NnlK9ekiH09ft0eb88+DJJkGmoICb1LLwamHEK/A4ju1i76yEQtppVmRjdtQ5vQ88LkdoBgck
3AyAyBgais6+c/eGgmvtTMluGQBYBYnd7ohQenrQYK+aPdsLxRBNaDOCcRKDtPBRNwDH6tth0SNr
cN1s8nYdNuJZyAnKiHjeZIo+71pl81larfjCR8GiTu7uKwRwH/xLNOiHOiRbJdZgvHQTMef5Wl7j
M11VRncAeetitfa6zPRjwxEF0HU6//ZnNCOwObKHFQiOL0EE5YllTnHQ5g/Ps4jCWTOLo1UeAdYw
VnFa2qE8keTGSUzQv1UvxTGQQYRXmXRk8mrsL0akWuiMzWnQlcxMdnhrRJ/X6ThQr5+kt7IcykEl
akqcU80KeBGcPsvI2kGj/uWYypqo8wci+B4hbggcceHyAvj8e2fydJOvGbGMaUg9gQXP2p8PbcNz
EGb1IiKcjMECJIObJupTc0hvQwiJMrWoCNORWGYgu5vbwdkd2dqSgzjsqoYhPO1TNJ5S9ciQktlG
dP8+ixOdQp0PIRmkzqbHpuIhhRR6XCJlxtw02o20ETvgF2XhMG8nhE+RenATW6fObAdfYfNCv8hR
hAG4GxPwcsLQSNALTLWU7iOhkAeodhHHsnoREKB4HAQXqcWXcBmlrmnd/optetBuPCz8YY2nbCbi
wbP40cNT+BhSL0wY5uArv+HxT7DpgYyk14I2fMG3CvMGPbAreXW1ekYonmdLVoWV5/aDyspCMOfi
1bY2WUlFT/NhwOvrZKn8CggZ76V6paENPnNVFD/q+sVl4kjLhOvGk8AKo4gbPrjVxSg97HhfNfBx
7JL4PeIYYUAouNLazsLx3Cyzk8ZisLSuwu6IBWDL/ZcLgRr1anuJqyxPRvwhutgMvgF1rptzy+da
sPEPBUTh3WU2ozx+sCFAhyD+q6poUtHYGFDGJyBtv2kO00ro9WHFYbjPY+KoHz+iFDOLTVEj0o4t
w8tMtO0mRUL0rAsrokOsVa53B1b32+20OBurQZt4vXk9e5cuRZnwSk/nYbam/a3NutxhyiblyRFY
B4P6e7Ac94zXA+n//uvS/z+3GH1dMC0yBGyOJJ6xDj9/gvuV7eyg1wogQ8u7J+dATwz8NOh9N08p
NwrjNzXhuZj73L5MMQ/7OD1bgMe0EPhQSLkNno3ycfE47ncxkHl50oLXJ/oyZ807fbYH+v2iqk8N
wXUBF9mLf4Qmg4L4JvHl+Y/TI24BqWCflcnTaxBrOEpISMfQPjmOBJFFEUd5l+keXDQsGl1J8hXx
Vv8aUyDeCtEilBvXrqUhpnSjwM9prRZBDMNbgucGDyp4nkXsf0FinFJASOzmn8RaVPwMA/6ql6RU
9e1s+/ADXJFsnUib+KSJwoS90Apxgtnav8NpI38oKHbGBgvzvOsHBXqwxSEfbiVbLVA9zywsNdef
zvIq5bEn3oUyRuAvqOrClxaKQiqjqwiD/jUkwKNtCvZnciVH0W/RYS/4otz/h7y7BTHYyktqty5M
GsPJyIYnUhUPyOVzLyhy0J8p9YApkrf72vG3qk9FZaM3eAe5AUSUlt44o1SQyjv0F6DaBh4+iT4S
Q7NqlQYu+IIPjatlWJ9+cvwv4S26D9GnfMs5GFp83jOyugo4uQszL68BAgsmI4Ag7fssjl/9o1aK
PB3S6KPdluga8ZRE6042hnuzWbREVbwa+dGbqnDBqCevf+cokRMXHSF+F6a4UxsyQvHkyi8FhIb6
elXToZGaqvPxtA9xlBUus9tiO0mAdiWi/pUHlsopNuNj/WYujrFo6Mv5GhJdXFn5ZpRjp7VzZ9zK
DLiAPLaadZU/g6PJY6TDq6sofyx/9VBSh333m1AYzL/KWIY+D4F50GiuBy1QvhiazrJthT/e+jL7
2244xcEuBXh9/N886RmMC01UD0Ymfmu0xl3jk8FpuOlfDldHVFjrKt4PPFPCs0tfXPDe7aOBRK+d
1hGAqRwGRH5E9O0+0K3ZAaafRkrPKXatDyt9deRqiGfbiq1VqbVAwHiYxCNRY+mLhhyxlOVf0R5f
LCYxY4LQ0ovAjckR9kGQFP0RLXSWxySJ68p0YgUhO05UK6ESx6bE5clNO/JqInJQlyfm5/gXxlKG
I5/dBi+pKQm4xLKH17t0G51aNOoKtrt4AAVvVrDSk0Hnu2dGRKEnwtf7+KTwoRywdhBCZfhKgkb/
Xxfx8IqZZ4K7WikCfG1q7ATUvvIQfLY2fCDhLqmAtgmsZGRFvNNPxscX7WLEXMwxI9kpIaaamMml
F0yqAn0n1aEwobVDhNpKzOFFtTRoHBDkb+m+rdLuG7gxq6gRVWpySm+5UUEFTveLYZy8djTY/WLB
QnpgfZfaE3gWaXrS6n32EpJQWsoJyPJB4ny/o416bDo9HJfqzlR2yjY+xY73ASO4Z0lyh+AZQxLd
ZMiT7vJlJYxgOj5ZRwXsMgrsqTcmWrJjaTXCkSLaAwsNswXcq6tnw2dpOrSYY5cwBNOuZy79Yom9
O0Zc2we4lGImAcEjBbxy0Z3775fv0s7BRHYdoOfLdbcqvjvXilvOG8gqkw/jE6KEa1ZcxFhQwJza
xc29RgLDbyAiwKvciT6tti4PRDpbx1IE1k9wQMyXw64ff8MfvHDhiVAhpuRpodyhi6bUpnuiI4ft
rb8qgSevKf237r5dHpRJUELSY1DllwSifRCCX+4U/26rUmwkEkohjkNgQAPJo5+B9/RGONxnlRFx
9Y3oN/uWtobv64OeDxpt3Om4niWyiVku5JyvZw7bevpRPDzxKLLYlhXtssQuTFQTjFX/pQtPOikr
lB2vkK5LBllTB3j0nGPa8c+oncuoniEa6+b0jXO3+Kn7M26rDDbzVPJZKS2HSh7CUB+yo5tSqVwM
nV96juCBg4dbH9pGsXZ+sSXmyEI/wT6BrfXPTbNs2PobivxA57rPJJ1qsdp0izpWuy7Vz3nCbFtk
oRFM8WaYCJl2dKSU3R7seBEIP6jaMMOMv8ib3x3zvHhJLyyHCqXxTz3qS/6YVvQUXMb2wF4Ov4j5
w9wRV+CN8os4IuKh+LRMT8FGxB6OM0QMP9gridaWDlNGyw/mtWcpSGtSv8tAcbiPL0VWxz+hJUqH
YaoU4oTlXVyjmrL+sCsBDdS2Z30sflLc7k8VFKanSQVH8vX/C9To/wml5Y4w9PLLzEMDmMmqshaU
y+JRoFBdlIWjJW87yILLdrpVPQLI9r3f9E9Ob9ff683D/oy1u+/6xdMwnIDzchKlq8YHXPikYhIN
6Sf2HUZusYsHWm+Wh80peylNzJg6wTWTJ2nYqGoVxrfsnxt95JXAu5ZkiaSh0Fb3i+s4g2OUmqVR
vpNY0BsFtXTsR923CjvATZb6/hOOBrDKn7DCQXaZ8EhjVX8Jne/x4DyuyXsgwULsxwUZq9BbdG5O
utyr16OqTdgaOLuIyOJIfzMBVkk07o9kwJIdzQVdriqasMmvn4by/3SIrLdnw4OvVDenO823WIEA
+geGtaqdSerIfB9nPWbCaBvDB0KUbWdrzkUIKuLxL7dNJ4G4rHq9K/Eyw/y+R13LsGzLEwgLqMhr
Dp4ZoaUvaIo/fDTHjCgy6dF0tK98f0hpST6wepZnRsBVsL7TAPno6cikRY8NQOZm8o9KxyePDvtL
P27aZI9H7XahLbwPWCqW/aeFPlhLhOn6aCQ1Y3aob0RtI7iJ4Y+ulDnjdpEInVDwQUxSCfhu8/Y9
zQ0hw1ibLgWlc70FZe06SxuSL3aHwQh/bclNqLOhkKYmF+o6hoElbSsgLgwfSquOtQQTto2imqsJ
vRA5pl2u4uR4OG+Fr416Uuh9tE0CxHxqri1ySuQC17comFvBIbQwAUbsFd3zCpvus/6aqu4sLNLf
gwkiOnpH4crLraYNQbmDhRR/rlwzC6b9kxIwZ2OoGs8p8HafVNrdlSpDfiaECo6X4Tm1pYKTGeHk
F21vrM17Jo+Ps+hpTl4M78sdG36idPaa+zpyHsq5hWP9/kb3sY44Ea08zw83mQTP0v3+ZBFcf+iB
icIRw1XwUuvH5LISjEgecN8jmd4cw0DrXguXe4Uz8z/CJ9mhZhivwFTQfgzjJZf3HA4+9xP9CIIk
nsM3Nmig5dC5Lu9M+d1zoY3iT8PTeCOesEvTlefoDbpYcARHIzTN7Z2mCwXYHdJu3afuZmb7yr9D
Fq8sGmnAl1XobR0dsdXnxSWi80SMUdQFwQ3rHM1lPqJnEkkpv8asp5067uGXmlN+fMypCUXHlheM
E7M8YJ1bI1C2YwXYpAG7H5w0e3cD/hNR7lLvUICYGbFaoUOUD1P5WbrGN9TXf/FBhS9+I83gFY0t
Gn25R00/RFH64o77xjLjyW3rWNTrcqtkhgGNCyxvE1+Qi3BbV3SndSdXfXW7Mk/YnQBKOON0u49x
M068XBJaVbWCREtQXkt4FoqUydeT1hXZeTA0lUPA0rpO2yymxulP/K5W5+4hJ0GY26ugrPSqQHoG
2W/LizHM+odHCpe/ZMANsjYM4B9w3dnG9gcSPnoB1YQgHJTgc1cdQJmVhZEtSnk0OV9H6UjBjQK4
C4DBmGnc2xd78+dSkbYfvF/YI7e5lZGFYnDhuiGiZ052caUIfSjnSEqBJ/3wmhgVugdOBhxjclz/
K+TeN4aq7+ODZqO2LYo/SePg80dRsxza8wHkVyyYOnuSmAweRFKtfdWSY88eajHq/0R3gQ1jgg1T
ZBKgP9pOIEnvWUZCz4Ul2VMIRujCuYU3oKMDcMJk5VNlOsxA3JureSPPC1jAmthuRC9UBF8fI2cp
wYz44MUUrW05SYRcwPrBNOz2DW5C0Arf7rZ6DUmTjmNLk50ZP2O6QQfaz4XslTZ5ycQu5E9UEweb
Dg1uNhV7MJ0+P8LpbZ9uFkHMvLg/EtG1ZWCj7HIFm+sdieWnzbpDa1TjWd4gF48TXVFVT3we9mpv
vqwcQITRGE1GMaJXLgKRXqyiKm+MNaN44hJsrEp7iLVOFLPGoDqTph+fHQdg19j78dRmd7Oxiz+y
eEACCacwb3Ih+sRJNzrRTDRjUvCFUly416aMZRunX6wDz8nEE7SibuMVFG0chkRLjObMa+l4SNzQ
eDQJEzkRibGNX1fk0c0Z3HXH6cpcpEXpQit1Z8+vXmqylVVemG+CWiFcN1imK2DppkMnaMS6B4Op
7QHwaHNZaG2vV+WZpQtG+/jCt0sOb9uQsbjRXW4F+2xl89H8rDmWljif0vS2jqXYv4g/fGCuvlMj
JJzqYQtViAIfDO8UK9/992e0oF4YxybjHlSsJAZy4t5Cd3hB+maLNpFFFrT3IwcgTX5+b/kr4kfP
lONBJ4/+VuhA1nme0TWQFi84C3Sx53zNINReDN7VsZ8899a4xhEt0bVKMMFMBy3bDteqYgS7wgQy
mi8dmK8aH7K+5/ybDdUNDHlfUZbK2hPIrYY4VwGoLY1AOqgrOyU6N8hX2cGytSTvG/hzFGa33dCk
B8/EEcF7gTFg4A4MsizfMEedh7Lsot6+v3gvsJbyQv1yMp7VLjPQwy5LB+zgcobsyZt1v96WAF01
Lx0imBPH0fzxH+NVTFjMa1mrk6a4VdYaLw6H9C+JRzKtPKPrmHU0BI8sMvL7izYUNvsw//kaCP+/
8uZHU0SulfjuFiqPgvAJ0Ik3EK408RXgJMrSXILCPKRlLVvsrAYclgTRY0RA9VyQUSYqyyaAxdPe
b5iyqU84ludNvfOBV33lmn0/WWZdN9VG1h5zfJkOWSHc1WNaZKC2/v0TBrrOWW4r2x7r51+g5ieB
7Vd11qjMdxUAs2/Pl/jM/N6zwI5jn1fTIr6N1/XXAP1+7WPXngPfAHbGZCKtZvPwd3TIovBHb+0E
4stJ+Vm3yaibOXlTHlNQ4xBMlLt+FUaUNhE6rhW/8ZNJwGokBgpCiHCgTqPzkqobFVOdwIH/Xz+2
hgBMIcbb8EmpPdXkCjWuU05DufhAMjXVtizXOAYHVCJB+n5O6Yf9O4Zh4MPnzmIDEtI2+mk7k57X
XXLT2Z0s7m+iIRlXV9lFcRdrWO27bSh7SawnZzmomlRd1rl5XJrt2ANhY8llXhm2YOE4dMTiPgL8
5AklpWyBQc/n9whYcD4oRJyhyogm2icKkhL8VYv63i4IefiDmLRyzM/zC9yOCeGjS/oAv2zUqB5S
/DAHTxwC/nox8207h2ONVdP1++I95XO4od/au+fDtO7hP2rAa2V51CKoFwJ5idZYOBWt610mtNbK
aMtxQh2iUR5DR6DzyYhIQYhN7ZGn8gpXH1USo7KyYaypLKeuM0kOKezykffp12eEp+gBjEORfweJ
G+XtC4tviNtSA52rRiMPyI/EKLf8SXo4cZPYeaKFj/P4XeqD5/CSBYR8M0CmLz0dyCnUUsVAJ3MR
ISaB5PgZ6frAJ+/AF164GwXOV2XsSe9miyqg8eILi2tZMuiyAHu1hqoNHDblBExwkr4Ees5aIoF+
9v6CcPalFaHsrrhOvVZl4VF7ay8iZ4I2PwlMRbs3rl5kjL7+0VAeSX+2vdfvtLzB1l2fAKcz2+oV
wSd+5T1S5UX7tP5il3XdW04E7UMHkSzYwJaVOvgcolHXsBTeeH38/ZafZTThNf8rkok9a98vnv7z
8C09Z5YhmjyqnJPwLRmPF/qtjKnFicb3DwSY80+sJDJKz3OscejtZ/SwbBpV3OEAf5I08oKyRLa7
Y6S2hlni03zEnlCHaJE80yeYXIVTcQJrkfTMschal/r/gd29A56dtggpgmuReQ0i2Nd194OtNxKs
HlD5BK5vsTYnMN7BWPGvxVXY0/Up8Ev1ClDCvcwiSSUR1B9kBhPr0JJmgW0Tjwkoexl65CgCkcMQ
AW0pKj2S78+UC5khEVlkUNsSJBx3UWdWimISmJ0p4cQOPa891NTMDKRQ6jYWGFCWkze6/eX1QZjV
0Bcx2YPy8rzJdYffg3BiK6irqQ+a9EUeDMpvb6jkRqZqLNm6Kvnk3jqxEK2l7Dc/YWb/unVyOy8J
UxaAfHYrLdahd9kHthGC/ZnknKzpvZ68RDa/y4Yn1qvrAD8W30i+ig6ioPOJAkxttqQuk1PNv1iF
/3Ll+giWC+7azKVHQcB/fOZm/SPEOVD8h07AtxSVG4qj5iYs4RVexSWtGqe7F7Q+XTzoWRSEsi8q
reXNS49pRBAjdLY2B6WsYo32W0s5NGyuQ7YgOVzE1raFEV1iaq4lmmqtQNgzIDEyoK/kJHPxIS39
+WVLJwXqBzhB1mWHyYxMqhmVP+9YQuKNtTNFgQgXwy87z70UQahJMtqmy0OGGjwNp4W0A0YeMWrs
sMM+9VSAgJh+hTLTEtQF0jJMXfJwVi5WoUbLomfqku2WQOzpupAS3Oxp6/ihvaWBv7AMmtypAnxB
QcsYWkZvML18Xl6ox34OqTFb4Bpf5yj0z4Iv0RJdo9mVAx1BqasT1UGPALc9dbnq1oK2J/u6WL2R
7AVrnqNmErNCStN6XHEb+gdyNkxxEf1fizSewn4vuVLslGMOHWHW5/Er5WhC++UnXCaR0UNCFOwO
E0WYOcABuESVfgPgBf9fd52rIwkP95l0A+eN/Y/S9gEcU3rHdQ11Rcig3CH4xWw3oRUi+wdtaFHu
anTBoDF+EHpQq5/R5+dTozmGg6fIC/j+HZlijy04oqlCAHFYh1JY3wMftflClX1hEZbBIHuKUNiL
ZMZ9dwNGKl5qLmyINr//3Mq/7f2bb7Wla9G4s0HiOAw3oH70MuwBQ74NomKbbA5ut8/F1D8bFmTr
IsFMEnVdFSxaslaAmx1n4AWERojGd/LLCbdbhHpP+y5UqWBJzcMbDwMc0EOD5X04GsmNXr7h4tb3
CR/4Y2PjQPmp2FbLdXRGB8Ee7dL7n+nGRf68TkggMOgJ5YWik4i5kXh0K+qY2QSvLAvHHrOxy++k
dsUgTcFfk1HRec2L3GyNWcni0Cyt26bEL3RYxqCAFoIltz1PWhDejZyXF6cwe3oUao6oMgDwa4fF
3HqGkH86bMqfyIqAksxrpBL0dag9pNSK3TvE81s2KwPk0vtGlbV0OdOLBWhFpYN9IS81UlgzuzzJ
8FR8HN5EDjp855iGidU01p4jUC4aFcqt2rpnixw7W25VD0S1siZSsgg4mKK5hz5llcsXzwrMZDxU
P5M1NL1cDgx0vgQpywTVrUrAiKJs5tenAye19mkF7bz9ntMjP6rK33uBopZLf8FE381wME5QxubF
ust73AtiqcUs6lviDyDYK6bo2R/8fUXBj73trTrx6Ivryb8HTMMVGyDxLJsnv+as/Q/a+LfgfyGc
MUnw7b/YGwvEtkM72Pcs64R7KpXf/3uD1JJwYwmYCTCMvypbR0SRkfgicsDX2yJ7y4/fYrBV4okG
lZv2d5EnWbjSgB2SjBYiMUKvRLlxQqmWajIbONky7DbVRSHpnOLWhn6tRD2BGgd3sgIAO3jh4ry0
WpxDde4kBj2JNmCOxxdrb1F9+BCPq7Bo8wx2C/cq0Kpa3Rh6pL3OKIU6gKaORkifTXTsTPjCOouo
DBsvLZKn8BEw3LAp0ydkQ66TdzGGyXwRQF233i+Y4s76NpDG0rvs/a8c5REgvBodvVvxsCieD5Nq
hHSBANjAcC9CO41ssaj48doXmYDbyxpBTP8LFAZNwJMy7CsjuXC8WfkwkASL4HYFSs/1m/FlQ2WV
NgVFTFEsphwUofeoPJ1N+LZ3mtNXqjwI9GpoK8582ox3eHKoouVNdcRoe8wndJeXrmDewDTl2HV8
8PJhOz4nyt3AjlzoQjx4rNNlCKkCKd1ZYhSCqlyD52p3U88znO3As0T1tNevPmwtPfJ+E97m2boe
Iib3q4o4yaR2cfi2Z82E3FzrQJmaFb/5RuYmOW66gx2UZTy58v+dvacd+VnPo3CPzxLO5BeNVrBN
iOfl95y6PArQ+xDhdChRo4BRsEA2on+DwY6PiJkXAPBpo5ic2vckkkGcHDjo/gZRef4W3CZ21X19
AEdGbPsgIfuzuwIyE2HuhrMQFoItVEgSfdDyA8Ih8OveTyRvXNL+Nk0FYDGaTGRqYucuA/WIRGoQ
S6rgQz8ZAzWAPgVQ3/jbVu3NubjnpEJqYDEN7YLd1QPZhX11t/jgu+hD6hFDhnBpZcXtOg7eZeIm
mqku7j/SSiIQNs0ptPX9BkWx9kLf8/0dcYneD+OivyrkKpg/TJxYQ3Bl6bbuZnMs+9cxPhn/IjzZ
Gs3yhcotjPA3NXyEPCChLrm/XQXsMMwvE8q+2uYe9whq+H64wyZoNnjqUZ0x1RbY0qIx9zSQRJhk
K+FxWoekHgg77tD38JTVcmJQ1shkdRpogKgTAeywVIKFde7dXjEGzV1+yDhj8lBG7TSo8MMD/MrC
B08+6A5CEJBBowUjaMSmjdxh3bueAyhx5UGpNYW7Qq0bWt09MhcHdlwUS3Qpv9eDWkL+5wtrogTk
PjbgXXtUf7Mtwjyiex+Fxms5X95VSxtvE3bSgRZDzAYeucifD+RSrqsJLe5g9Yv+f53nA3enwk0H
mXC/xHPDXgmmtkhcriLkz0hZhZai4JQ8kNefxRJ8Y6rS8MJyC61L1w3ZaqpMsyodckhf/NAWimxA
NszCS/59E4YIOPKGEdW8RESHCvnnOWcOHjxVDhHVv+GSltiHJCO24XVYoB7V8RE42SuA7PNudgCs
ORmK4SfhF4hiYuNk2XJoL1oBGi6ziF2MhdcVNIQBmfbRQLO49kM3kSmQNcbFmDVrAJ8T5KTZ3ejv
7MDqXD+KfHgFvEnUSMTkjouP8ryATZs9pYplz2dHuIDIts4LhkS7uNb4Kdd4tr1dT3z0gVzlE+J8
xl0tP9LKciKWLXsoHTGhXcdN0Vs+f6AYtIta+tNeT+vKYXmTuElz9nOzxXX6aERbd4bPhBHPM8Hu
TJmdZWnZX7MeMN5cb8epBlOkYy3Pgn0xvr1eF/pP8pBceauh3ejswtbpl//3hYuR06HyNTGG02bP
bB3tC+9nqSYV8e2xnpzb+CPKvFkEt5UTCZ5VKBRvU4KGKvi2V1xFK9+dcAK2MH5pr/tjEl+Q1rec
BfEgfghDtlGgbuuVdVde6tOb7Bja0sdvHti/NmIfgsvC94xtAqnjtaVvAcPGwczgaAFb/I+87KDw
rgK7CQKKJZURQvI0HFoRcxPnOmgOfqEsJSrIxSE1FcvWkrn/YlVHHzQw0kKiVZwk8OekXOaJMKbE
zXjfmfa+D8flbXyr3ycbqNk7kTFzD48jdX2veONM80C+yIjfcb5fUz6+wDbR69PCHFYdwGDgk5sr
4MpZjbVuABS/dBNnmkYjIgEzk3fp1cJRRBEVL67NaN3qqixfQszEsw0jhe14Hbs56liAGZZNsEEW
lzJ0hWpkIFVkcVm7Ya3t/PSUN4aKE0OqrRINh5RfbZ3OFsxS9+NRIiSPNxcWLZ3jxiN5iBuxq7UK
SsMQ97vD3bzUz8mivgxLMCJRoxmGryMMUBHj3C3my4MyizMqyQhvIkSIXfHwjs7Jdm77YtiN48ya
wqR6x/HiNGwBy2Y9X74S5CmYvJdCVWBxmQ9CpZWfiBO38XirkT6nokUaTZL2dcq227FT7z2ywA9w
rKHR9cXPTzCtEb68+FzoGO1oHdRMAot04JFwih9NTQmKYOuzK8S4GwnmDCV/2m9AGSZGc7SF828z
X4nRJTmFpoat4zEYwouNezFo1ZoeWV9UBthiFrsKu7Bx1BfF9/yKgQ7Su/okIGjSXo2AhH3eysYo
QIDyi6eB9onIQZFSoT8X0ASLyRGbxyokWmUs9yjc2Jm3kkdKqxxEZttBUpy/yPufTnZM9vbrrmd+
5tC+3dgDqlpFYVQhan1BBpkccjx0XMQj3vK5IJ9hjzGDpmyKeW4FThrdEL44EcAjN2nKONTrMHY4
yhDNV5l/hHEPKVJKhuwfGD3dt6naDdnKut+zRKShOWadnOQhOS5a4pvARV9aECnSnQ4R6spbjLSP
ha/8Yy4VV/yBtcXHttrXsOu0Qk8gleKOsPgQ8i9rIUhu0V0TeaDl4301ECe2xFobq8FzSDo/KsrV
hgruvH2jJ1/0KycXbhorCKGdnInX+TgF9TlHmv1UUWxMoPKEee5i0TApV6l/jnXWMzn9C6esSlgA
4ObvhovFl27KLwao6vt5YAW1X+AO/7nTf8peALwT7l45NoGLUjYozrGT4qr2RhohiZLmuDQ5LJ9K
KuABwJTalK4oRUxdZyVGrgX4vGb86YkDqtZapc+RAc/vCejKpe61XYimhkqC6sjZVRCmPyL5AWm+
0Sgp1LwVpaThEW79u9xLzAWwC57Nl3bNC4qHKQ4+exem7HOMKN29oWHNIta3NxmRlooWpdzsZaLT
2QClhz0jgEG3uUUwqr/NCz354x6f8v5AS9eEjInFI4uLq2v9Ym/TKaISVh+rmBojfeJkos+CPDrn
DzukIHP0/dABgynvYRXXfbM5EIiiYXT/jmZG0+vLPHnCIe/dhbIEengDvL+05GI3IObHFinttSsT
wa37bWaof3qlPxDXubSrVmN2QiQ9O4PrCXr4XCq0PdMD3V9D+QLlRSU+0TQdPfKTdr39Xo9Soq6x
oN1SBoUJ2O/V2QYFNuPXkXT/oiA7ZJCpQh0RVvzbrQWfmYnJ8T76cheT5Clym4fIQ5TSoZceYdap
Jpge9/dp8sEmsKwpcEbNLMYdyWVcr8ZdYkDCFFjkjjSPgVv+/aao/c6AHOJFDpGBPYEw9AzZPjCh
XPQfHtG5cQYJ6gpsnJup/0v+rfKOVBYnb9oZZmA/6JJB7ZJVxfmHXIwREX1iL+Txc3sj+L976N3g
4A2zQ4pXb/CBjf3uamVAdYrjFgnqCri4yo66esKm86j6hbIX1joxyBVbY+yslDY/0rCXSHNJuO2W
UKDp8O/eTxyR0PES9n4v+wB8BAx+BsPoO4slL0l4LuUlNdhzDySeuurdvNE+AIvBBoXwuCeEF6mu
9w3MMYZWi99eSGppwruPRa/cmHQat7piH+9GFUQOzLSdxEvygEUUHqFM5n9AQyf1XLIINsfRoEm1
9RAQTO77qwxtzzfOw/9pvJj3AAIiXIPlrJ3skhRmctKjcpp2Gs1i1MBC/Y3NKrYOPCLxGdls8dVB
49F7DlRIqU0Ja9WF1XJk7vAhEPJ/VLfOGQy+5Y275WDW82eHrVIv7gedbQvfWM1nMjolBqULtRrW
ZBtiByfPyEV/YMlqEFPsu1SELGdmwwROcPzOgilGPN1gkfRoyTBj6bQhiSJ5kmL2xXdepJ6NNjKh
ySdNof9ZnJ77o5eW0tsay2QLBuMg/PW3oo1k1tqRI2czm11hJMZrCn/B/GfkBd1Lc/WEM7xFyeVt
JYwkkZUQCoVWQ1mK6c3GOwY/bsCHxOgel9KGTTgQK6AJEYBniD0NXdzsOwRMyenaB2NTcKcCnHTB
pKHzkRFTA1zLNU4KERvxxt+ikBdbLVdFDdHolafuKYbHO3t7AXs3ZDCWhDsxC5fgBmHltdDVXE8t
G+nh//Ei0IPZagKCdu8OzAzjP+EVIEiTRkiCxebWmoBSVczFXK9D5sM3IYkKRic/7qbOcrB3yiEI
aX2CsuUK+SxREMZXZjkGZxkqNQyqdTEpa13669G3jrDxLgwcRswSg+UhziA4h54tyJ3Uk8FcKeZ2
d3GXWiuQdA/xq83OGVNej1z+5KVN8zlu6amqdh0qQugRYB5nDfMEWjF1Syh7uprMCphGcuOt2q8H
/BS3JmoHKSPt+H/Ja0E4Shqm8Ir9Q97jWiwVPWkWw3tFd6JlM9el6srf0UJWGjPGkF3ghYOfID0Z
3+dxIBJZ+Nh5hJduJFqXCp3hdijaO8t/uCY/rVSqnrToHY5Dhxqo3/Qzsypyx/WCjs+5hXyHVLQO
Nar/LsqVDzMM61tizgE1aQNpO51ztSyT6Uav+CKpVdfz4rcC7LQuSMTKVfB7psqIjwnWz+9FZj51
I/EUtYrT0gEIGUL+vxlLIUvqfX2nNE6tnLaCEp8jAudd0UC1IhfYCDZiCcbpGV624+cN9yyNWx9Z
/sf9DMov+1UcH9OkOQHjNirlv7O7rxOo7C59t+bkUFCnjBoLhnVP8DNSot1yXHYuL6XDPdsqKiKx
QidFylhzhlqgu0cgv+ioQfHtf3C9NzxwW1h9wEHw4QwzZJWSy62s/wD6ofxf1houp3GeHqpy0G5X
mU5tHnBoJbIWudyAV0CHiS1C0WIFcYUPWkiiCqeD0XkUSs9lXWJsMb6iqWXyqAytvGjl7hhXD1LU
uwtEwT+JA7wIsj//rVypazK2NjXRh/2wTiPjFjLvCKuZdOywqvdp1LRaqS9Wg3eb+7emMjbGnJfs
NktMfgejiT4aKncS1oleHxiVRsqWT/XhQ2f+fJqXobkcb0WfiVnnt1aifrQcWrJKw0VlzQC7FTkE
4YTLdbZcbmxUcoBlZC3z1GK3sCh/S60wnOg/c3F7eeD7egIaK5gluLT8b4ZzEvdy+17eSgzY2wt2
DOuWnyStz4X56qz3/NekICjFU3DFG/GYLTwet3svhL03kekOC3pCWsjCm/uKJeeWis8ITy9OqKlX
/bfChAsLsbm9lbY8SG9WcSge6/9bbnrZ/7ActIIAkXKAO7MO/jTuOrMHkBAZh74+nm7qtPxqU7Tf
3Jgqs6st4TzVIfTuUa7RR/jUFPVBRfBE0vSTcLyRwczeV/VoaYnh+eCjCb7sMn9fNNxooBEP3wer
a7wN4W1aMVpioXK2AeQIKAK9TUXlZSdy20I5fTH9knpLowDSoeDVVVTd6PNj79o3WjnbI2Ie91mm
zGBIsbIkId+QENoKEbmzqD9fk0wqI5/OjEmn3wXBc8ul+ypOjtEIlNOAzmQuKKBDCNwhmTiCSiRU
XhogrPzxCmWaUhtLfQagS6yIBGEN8zTezLcc0be/aVX6kquSQnjeZBTGnkaGdgDgac+30GZpF9pC
eYrM6RHuC2p8mKCuOYnVyLotShFQL9WRUbkDO7003PTM1Lklxr0odCRO+9I7+yNqrkiVHPPop1HY
/BmK5awgWCDEOc51f86AFF34GK/ZCGxSRpH42CDC6bHgh+XpmaH3MAiA74aDn5lglxFKgI6KYfD2
As9BreBmu6KjCPA4wuukGVO4svbx7095L1TX5Vf6c9ohQCrM7ysvSST8f1ewdz57AlGdIM/d9/It
Z4tWIvi6iTieon+ktrG10tyaqOje9vAooNoPd0ZML5j2+Ls+3WptosoyvNob0bxYAI6ILCpyFRFf
C/g9ObjgQRMVK8Bt6gPYmccrkps4lQGxEgXY//AybgZ2c24D3+/xu+c4RSHTlomsc/rYC/VQQdr6
Nu2P4h/GI6iAaiGyzk0OtEPNStT9fZJHdkEN+UnbUlMxEGZSNOuScAadoUV83zB77wbrLudtWYqm
hKh/OHufMqE2j/rCypezAdBdaiCUDB2VQCyDySgTJOlwM7ehxJi0OBSPadhn4nz/DQrA61CAuzGG
zgfq10wHZmOKYgNG3/n3ZSn4TazhpTTwex3Gko4kXYefb+uTRnZ6szdDCjQ/g7Poqer1qW4e80pZ
VhOeEkDZI2nYTJWymjF1zyvycZfAdlgjR/vUe/aO8/0N2zxSFyDOc0I7SoxHjkE1bzCRfJuUpByK
gpCuYAS730VPT+yBoHP1cf2EyW0w8YZVdAbeNu2FwCiheAVoBGyuSO47evYCAvSDwXxY19ulJO8L
rWZd+lKAlcTUIwA8oalVeMdIPay/PsA0idM6umTUOtynIYSKeTzLy/QqTZjqiq1ujRFBBy/JGPwS
mKXKvDOltf7bH/Syl92BA7XcqINdQaUO5yQdmjAn65cOIwEDhX7HKUOGnMHc1UZQx2GtB1YC+mMA
ttywlzFOwNnh+oqzF+bTED2WeFgGZDMxW0QFVP8n0ZyQbeUebq/jKaHk3SE76guDE3can6WN79M+
pLZREYg3TnMwXCcKcPF/L0rMeJW7gYBRtNq833mSauHMVaU+fR/q6ikf2dLBvA63PsKzR8ikf6Uw
m9qfei/VZj3dby8G3PXnDmhARNrv7Pz93NcHI+whlr/OEkxihjgxANhpJIDnntm7kIcVV5/hqboW
z6uIZi5Rldg5Oig9aT2LxXdUS+k1/UQ/wc+GBY3CkLuVLNwCrBZ6/rCzDqin4K8LT5zHXj71zIqK
eGNV7QOBPwWaWvUmVR2dYzgMlD1E8KMF6dddy7KCO7CI5+2ndFm1ERQeFfL8hvbdMCJWYvvExmET
v9BLJ8foJiOYf5qs9r4tTQMtkW6ykNbZu0tY6NXDCoCgHiqJz88yIAYkkb0z3JauNFv1t6YwII9+
60a3lD/zlNOukWbljZTZFV8wg953hqaM7GCB++EYNt7oWwKMwl+naO5c2uhSnI4/ACfsP97iX+9T
IWz47iqGeu0yY+kOJeXg/UlayRPIny73Fen5Jsew2mh9XHaz0caaQYO4xdFXDL66SGTFUBebxW6Z
C+MEB7+EjKHbxR3bsEwHTP0wx4svk16bEJ8eMa1aB53Thh4s8cCdwEwIvgz9wnr4owLxTQR0TGKR
Xq+dL/8zqz28EuoBzHRU8JPXlc3uOC1SN0mOQuUFOzq7v4cN+rHMWkfpACx4dhYQjQvFXoeNNQ8Q
bQc5CopNTOTUgkboqRzoheLxf8SWIfjIXlC1VnUHpDyoL87UWGjEpy8z5MUbpwZfQ9BAU3Zfct2v
H7q6c8srhua4uDAFGdZjELJU+qBOzNak4Zb1GmUiRBDUBI+4DiHkHUYrgCAz9TszuZCr6rya7uJY
HYRTusipqD3kQmETdpRB1JyjOywJgrNgCIndEqkAZmQTPX50zhyShtR0ARVEVvnFgAAR2ofIDDaZ
H8yduVHBhMd6bopyHbVAsPhK4zIIEv9XSCNxaiKY+jN/NYkrD0CuOvsZhxa7WITR9aw8dKvMdGvg
G8nVT8Cs1rR8ygSV8iSEy+nR51JySlPCg9qJm5gizUHEdeNBbmfb4GzYlW2wXjTzqrhJPe/VvDo0
v5P2V5d9xBsmU1JQ4OtEvtHcf37R/8zzS4hy3iWJbTWsyE8qZ6Iup3GhrEk7OfmSrGwnuQ4nE4HI
ixcuPUUJCSxlPfqY+G0p46h4p9rxRBxQ19wiGMx1ePicXbKDYsRgoRkenKvjl8t3PA+18dxuH5bk
lmW0+bgowzrWLo8Wk6rCW+xekZBzFxpeJ1rHR68GZXcWotU3is3iIbKgxzoq803FGHgua+1nYExd
G84Gco4ZU0ySB8QyPU1Mf/wNcv2SscNv2tMnvVgIJesBzt3TKCceZervRphYWnutY2t9Ol96l6FH
G6eZDkBCFxAYoQep8+XT0nbyIzwXuBOYLcTNgTsVzSqal4H5D0PEYsGR/UqxuJ0heMcr+dFL2dgB
6fZZRMegUg/2y8icD6hDF9xdturLafaPr+8TZ+M+tVm7VD835T9SZfxK8slOboFR+U9ZBTdz+ui7
Zxf9sP05u4t3FcdsSl6KasZN2LrtbtxHukfLiYq62hGlSbbqVvfVHHqvINmy0Jj0/Gd8WcRdlX6P
1Vp0eBKWzylZOED4gWYXlAh6dOPv5gUhhGTMh7zQDYvyLCearfkAUkJBu6iUByDUq2afpZnzoH2z
y9T3CTUPC/f+ePq+BmjJ2Su5OdudryLILFvbS7nm9cGLSSnvLJlOgUIqLmFb7KeI+XrQNQs7ihC5
rvAMKt3L3TOdv+O8TYBXuiUm4ujQRpUKElggM7oXiYOiqoz/hAhT4WSQi8mtqpgCKTlQ+qE4zd9E
fVGTpElWaWGvUuceXHYVBOu2w5ZNokSOWz3quJYHXfScHBwY64+giyRDwjWL1FBSAZ+dENV7XDOD
vUODpYFnoatb9h6L2htBDO3jGDmqzXjsQlCqomDnNJF5iRy2nacgXwScrq/eJzF+PaqsUpuJWJ6U
hX8OV71pqyrWKiis3JW8u4/uqGHB36NxBJxnJqK8vvlCHchPoL3R2SMSslDprNAkKc07378TrleJ
d+U7rHblC+A7U4Bwm2y+fN85Hew6KC07xGj8/HhENlNVd2KEaDwcNBLYzdwH9pKFS5KM5Y6Wh3Ak
s9kcbjsLuwDEmVk8Hl12CCSoaSYkaVkZ+AvxEQmxZss5qoSBmtZZrZTe8n16Miml3ObDEMZs5FYH
Fdy0CUer9pMqtL7tD6zXt1y9urkdq520c39PdSkYLsu9spsyuhTUJLGBAQaMZrlANDhtNac2IaLt
qc04GkuwdGgT8JbExdWtG1YKeYL2fMNlKcgwc/uroVxKLSabSmOcHooPHJYA35IFH6P9YB4/OlNL
GhyLB0gCubBC/5bNDWEyKcET3Q/rCvHCAIDjhft4Mff6rFdJCyddW1UKcQIt07Zen0tC5iWqEoA8
f2qwaSVAUWlJahCYR9+I6+ibXHcVoj0lTxKHWKuex4jPfRs8vHGh9TjMCF4o1Mw4Jeod5Ok8zsLj
TQYTaVWO/zAOFLrVUnTiEmA21UzCx3zfbyDGrdNsJmVv61Q0G6aF1Ga1vcItf1jwz1X8OqoFTcKI
1iUSdchph3zuwYvDIGhW6A8CkJ3kUmwPxYWP71RaT95kiVjqvDuId7306S/x6K+yd9iezpv2n4HZ
ebAGugHGSsmJBcBWW2LTph2D2l+HGBenhLMYYDMyxIttew7xmkqkkReJMLgZumF3ElZccJCQGieV
fB2itNNS+uNC2IVdRlkf9n4aRNPtPB1y/QjyzJpqtZR1DhQ/UCSHQHfVRj1U/jRPls24aZHs9lWU
C7iCPb0Rp23+UFPm0VQRw+px2DKqAAzPLL5uSKFTLGRitHOH34Djw9wbLeN0d68y3U5ZasVp8Dez
N5/vLjTEGMWyzl2pL3QSl7HQ4ckLMEBE1o7iPAneZxbLMwSeelmCOWMdmWPWxS8eqZt3GV7lY/pi
8hsQEphDeonRtKxz1LrHKFQLS2XLTonwwAh54arzos4NJNNeLw/lxt1hHWaLLcp7FrqulZ3Rpncz
EELSM9/lVTMlSPhZPJRXepvHEQ6dE1IxOFFn+HJNmBNZX5Ycyo8T1N7U5TkFgsIAVHVNRdbv13Wx
qs4j7L6m8yrNRQ5Wss9tZPpFFb/aUTYyKuzwhoa+uKaW+48dIg0bOYtTej35vn+cY3c2MmK9j/7B
CNkCGtUO8DTwRfpzmK5UtRrrFMWAchgdaCP0R0e0Kp+7SBYH8TEfHWsvue7CqyLuCb1RZHzYxcTE
87TZsDDaomJbWMzJF5flz0DbqkrnN7Tj2o+n2ZnBByEO8u6AfEKSapCxLlucgGdIDWeGc6ukjSVs
FbAg7x0BHvW5H+tP9zM33mKXzNHgAyxU51D5ODWL79ZWIMfyRD4EE43MdKMHeKg+Bm1KmdDnYjRK
h0TbiSL4lfc8af7wiHO52ZqJf+LFcBTIMOAAxwHWzawqGmKjh3w+YWc31gzhIMQaIJk9n7FFDNVH
XVQMKxBpZ2HAeCIcccd5X72pjR8BP9y16A/Nr6lnmAYGCTJrwvxIfBG90e+em3eN4EV5eItqtsq9
kpVS9jTwrNW3f8kqzvPqbjNXDNWpmNYChsQVdMPcKmpSJupXf9g05LVqpryn8sa3u6O60+0SOZDb
xyiqOH0aOZJFOviSc9P+f3u/pxr+GnRqorwQVOtTlpI6APPMkm6hPuJZ+tOtlnMh3MxNd+5CPW9T
BFQYToF0meTyzO0cbE2O9ApE2xRlCzAxNobQSLKxqmjwQowX2wYNqIuKfa04teF/Yuoo5QS0k2V9
8OPv4n6UWy9yvEHNIpTWgCKWA5JdcOqTQCyzH+UoRsq6u6ObDtvp0P5BHWa86qRREFOGkC/i+gJ6
dj/XbihPUtLTCutvli6pN4CFUY1V4qVRcyErbpw733SqtfsfQBpNejFT/WU1QZM4fQe0bBjK10r0
77ySZNAS6D/s2IGpuCX/A/9hRq1h0osqbAhswEwaisGkDv9iOPLzUZJPqBtmTeDqBdMk/RuEL9Wa
9wgy5AwIbn8KgD8Vigp0bO1KnliUC0OQAWyjmNjekRzV5KeYSFLWBaBdXjC/8/ZINtR5lBLB9UAO
EZbesb5HViogD89YhFScKXcAmoNib9AQxQ/Lutw3pr8TcOA1ERZUjJHfsxhR5ONWLIv33Dibu8qr
JGd5YymS7TjwOlCHoSX+TBS6iO7yP7FdQyej6tA5qgwYtlO6i3+e9lDhIygb8O0FfEFoAroCqJZ/
iqZO59LerY7y9Y+KUKkLLFU0Iq/DkF7DiUfJpryUyJ2ddI/ztsyxIcMF05JKdSnTUoh9E3Fz4yNg
wO/+DZ3VvErCw/+Lv++38Q2oMufYfZOeKER7M/WJG02KQD3JPQtZt8F9MKYBB/pk4bjKeDfvmfjQ
FY/nQic3xIxRu1RoQpOBx6q2iQDF/QmXIrEXM9+I2Xd9Hb1ZnxExzgCkQym/OT1H0g0F2uypP8Eu
s0L6DUjhdFgDMegyhxqZw49rPgYklzAG7ah1wlTq0tPZ/7LBjJPNC9ozvt0pPqL9Xd8LG+mXxw+l
xJE8HSkYQT0lt4XsUxFeGO8X2jQLSsKlA6SU6NTJcMKCwTsKLpU4WNx2TM+g0GY2S6bRdOLEjYKI
hbhVnrkQiAxrXBGRvhefS1Qq0DKeVZeFothJSxfkV1Vv8auwh9yYQwgy8WJAwyFV5sIuR5nsWCWl
O6+5O+q6YH2DiCPt/MLJpr49ItEOHphu1b9xcERQ8FMx6XGpuJXfw2O4K5IAzATTCuN7qXYh9WT2
fcWMqbt4g/Y+mh+Tg6UtIeVVdnZAQjsIzy4yPk58Zt2DMAzoLVi4tS+lJA5DTXPfY/BWIxu8Y4/v
RqNXkjADmAsY1inTom5Q65vBjAzXrMTWjZZz2xwe9q2e8OOT9b6rtFvKDxHwtRx9LSZAF/CdJFG8
QWu6qk+KBbCl6DKhHAUJYxkYDMolat3q3CcDUXzndOVWgIqptPbj2cDOms6YbIvVjbnoger/6uLC
+qHSTY64e3iDqiwipTbk+wkJARnk09au0PY0KiA82w8Z3H88XKRcLPuutlHQ/Y3O3Zz1t8JQU6kT
g5Z/yvkLsq9/+irJARmEryfsrGkxSYY7n8eo6y3KydFRzv2fWx8Cbkf6x4gJU2EQlaCGhOQ+yDJ3
MVQpHPWWMB7+XlkXww5dnn609T/PoaLhgX/Z4ueuAMUHzXSpBItMziT9e8IciHRS0v2Enf+qg+JB
fh4BXeuHyoy7Ba5SG1QxHBbkTS+cggzaE+R1wQ6Pwk7jc3jMKcNBLHYKLlzRbta1RhHgkf+G2X8z
aC0lLiQazcGHYM3J2q7RDeIFpAu2OB9j9DNCEYnSidS4liJ2S1/FH+AOsw3dTcsg8+E9lJue82gv
H/63AdPdjVshNxKJtYO1jBDrxOFrSQ+RNDWY9Zf1n6lXiFA7HmilNC7kQJ2OYul0qQ7vWtr9g3z4
7tRPuzBPXdXypbL3YC/PjAUGFglIuNDJIO44Xa30EFOTLuS5Xbqbu/cqQMOtEA+2c4LQqcMHqoYK
HHJu98nnJbX6532Xa2WRUy1MVb+9AXlhvusk6tEJNGI65QL2feTIvcBIJDP7iySrIRnRW+3TVUFj
ceJtEzMhpRNmFLTDBTSr0oishcVrwgUarX26Ig3nXiwsXL6uyaSr7PuxbvxhUOFieNxgIjiGrXdA
w+YJznu4uDM5Dxabo838eLJ4RVuFX7ot2E1FaqM/OsyoGkGX6I1FldD4WkwoEY5AsvZE9kUVLElz
r5HzNyY9oCl6Ohl77D2TsZZO9zOdnly5dDgGcwiyyrfzo/07X6hNtKY3hte9ox8cpUb+D4e/u4LN
QfXxVOj5PgCz+oIJCCckV+Jd7/rPh8xFLGMyH0AVi56ZtA49PkG+pmy+7lAsLJN+jNEm15iwiB9L
w4FrveP7dJKXEqdm3jEEatZzxSHyNthT+8oAUJUeylfL8FMDGoPFj41ZYXlfMos7bOMLkWEmzMJF
7FwgiD4gze/OPPSflnA4dEPNIjjg+KNtAQVt7kJvQxbJJPHptRq1vsIWzpSPvDxzsbjHVgEz4R+i
FFQqI712v6cPaZ8p38ID4kqK3fC7KVaKuZYRDEwb/vCjAiUH+tW0vvqZe+C42jnmWDO0tVwlst8w
5NIzVLvfKRGLXDz4NaxvmCSE9ooCsrDohbq5xE7eyji+WONjXbGzzr31tHhdIR8UqPgjJpPjxpye
VdsFMSL0TMKeL0zQBMJ0CwyqeSp6ZmtP9XTdsOdsbboUuG51Dc9vq4FKPlrOysTUizeoM/Ea+reh
Qcyo5MejY41ddWv6PRlUBN54JHZRDbDzJrwwoRQsaeQk5QHfUqjCNkjxmuyZZjz0t5CsbCRvnzXp
nhyh3oaHsX2zIKjrUonLSoGaDCXdFTQ3NGBtV7AykeI5STlZmx/piqJtiIVU1en+lXd4rJggAVXL
93KZrv3Qx4EFZ4U3KGQ4XXgjA7qVoL6iBbzS0eiiO2iq8a8tCV/eHx7sZG0MkzMR76duCgmwQEjd
YyAKqCk+yCp0GyShXI16/Y6gmOu6ua9s/N+ovLarCrxrlb/xUPvsPWvWYWw09yBFVmY6YewTd1XB
zfrj8PKgIo4PQDyPG8JF0T+qD3cRoXNU5qUo59wK76l6sh4ilSaIqmC8OmMg/dhtc9mJNsL67ezq
/Ed8+qGRQBRgOGg3o2lv2jlvBWp8xatSZX7/skYgynCc+44vMgBVOTFQm7v41WDB7CyriSSQ2gWe
s8Q3fXrAYB+1tcBhK+eeCtGBL85oUm52L8WLC8tTrfd00+v10jcEnEkTciB3BT6AFDaQOIT2v4fH
HI9ZRlo+PLtp3QIv7GmIdt73+FYfvTdPcObb71hqwWXljFHc7PZn9mAx5cIsuj+wTiB+GNUxqRjB
PriIUtHsCzOJksEpJCjGEi/WgwHD0WwUSTqNOxfYJP1TVjSQ/iA6eVIgSaJRttdP8atgsHEUsGlh
bzoD6dboruuDgqge6l+zVEXeYbeXv9EyIX2HhGH//N16iqrMLRD/ynDn7hqvwatNN08jgHq168wC
ju3C4xZulHZhW+IWtkQbPZ9nuzJYDTQ9X2pp9zHZ6MhjUawbjLnEkg2W9uRddbEEL6EJS2VpOd6H
y5oeLcZ+bhtJ0AQDyQ3fgWSKQXqLOM4cpx+myGl31q611f/DtLrvfu3sthGbcCxbV9T/VPPzCtVv
5hwuHbtTMeYxe6C/9oAbrZs3cv91y71PlHk6VF9JTlR0NOTl5WnhZfqzrppQ0t6a05Xq3OIixif1
NF47MV5uBO7m5cOvb/eQa8A+vnVAV9JJcMk076JZ8gsu4DnC1arAKDqcBBEaN5EVr1tGe51qT+/3
TjiATpNzDtPPayXln1wNvXRO0HuXtYFk6SzB1XQuLp7ShEu4ACOxALOuGc5DeTVKNO+o/zOSSMKr
t1R682nXulUrsLJwnK69LuWNMXAIRZf2oBR7nbrepqt7zbY8RB97/HZxSnJGREeYjQVGOaBBWhTO
sRaDjf8zmqGVddkYaGzzchCUIBW38kqclmOaXI3l39yBGGx5bdszk7ww9FYwupsXBBFM/PdNpa8i
S/yFiCrIDgopeJCBs9v2b7SroTaN1lqMVGDFV354Tak1eTzvBBHsvjBrZlYkrlweKd0dbtNoFP9J
ffyfw+K3YQY4z2L7gSjkxCX9Vk1+9Pr+EqQjmIwcJJ/FYzVGKypVaLgs4Hkts23+tOSntOblU/BF
olYNLUu/1f6WTfqFZrZKTZCYxxynz0Hz7du5iYCaZE4OYTQ7INsDoRSj6XxUd1h/vrDkVrLv/nQy
zieElIJUim/gpY5/yLjQmAOD28tWQXdBdzgteh+7BwZ1oqDWujfx0LZIvXWtlScw3U6fEbQEEREb
m6XImqSOBMfKq9fuz22iDP8BYAPPva51gVWrzPI6rB+vFUXTAqWrZ0UhgzBOVWKXOjknlnwz2/tP
ztgW+5/cp891vd/JtPzIbniVYJIueztWz0eEhscyHuc5mIoyqTIG1vdZsfwro8PfzAs044WjU2v4
+wg7hUWuYak3LduGvsNIhm3EeUbw82/DO5KqSp4TNizOytTnB7tPNiBjUOtZQFACHHC9fVJTwxUQ
ILJajS+rPwrmLTQYAmv3zhA2SJSAyos2mHI04DcBsAlqFFdWgbOPlh8qqica76HkhYY40VYUqUl+
ndtqjloVXD6ESkqbnp8lVepmCitGm0zVvMvDbs+Rbc79oaB66M32Qc+ZSPmzvBRLVRT3jHKRJzqA
gxq/2xWsrZ/oAFeH4YEzTwOpsFtKpXGvBxAwP9N9kLw+2aUvm3A5uNkR/CgN5sEbG7naODkYyJRO
P/Yek3GNPMtQ8G3aQWjOk3vN+tBYiHuNnWqgj6+yLugrdTRsNDc86uPsdvSnGZJsC6Pl5DVNDp1g
P/OOm9KgNBR63DQBEGw4VCGCVWSDNRQkg70g/x7s9EQoutlDagAhFKDW7uacUTu7Emzvd1vCIkyO
V2/EaSolj2lrq+SOZj34wJw+ucPtUpqjYy0bqCd+BBab7qr8dd+RKCGi+vjhS9Nkn6TYZak1ra14
9ZV8FidcqycCY7WJ/jKd4x5zkEFXbLtQwtmqtPblShCSi4GgHcwiHqakVD1FcUCTueNjcek1vLhj
XRY82rJd7hnfoOusPi7yBwD7cDahvzU0PdcseEHSFTdo4XmXoIBGGw5n0myjg9j20rrJcO+4sRhh
SlBWi8zxtoN9TxP1oPSusBgA+QOM9WWWHmXerySrsTPaO3lZpJo6Wlds2lG1Ed8X+lg60T4F9TiR
rQTtuCJLTq4AaPaHhg2kq1g9YZn8xPRiqbjtP0hRCVLIUHWe89r1uEAExooLDwyEebUOz3e8ML/8
BjVHmIzZoL3uZhKLNFX+gC3GfZfdmfgtrsSfXgXAsuNbHD7+W0L7zYYwaqKwZrBG9c958t0wihJg
jB8L2tZoNmL5gqIji66OBAOcR/NtFK1/Q/q5dghkCd1tXqfl8twll+TXiYBf0kw9J54WyUvOvnPE
XVDwWGTcbJ6kxtK2Ntfuuk4JUwF6RyxIgRlKaUNqp2wDlVxxt1xWLappqQVBONktdKAJwOHqRhpI
MfnUZczQMwwXDcX5utXDGRiDigdyCTu1YDt+ICmiUZhaKKN05d90u8EbxmCe9YZXFlGN59Cex5db
gWhrpcPrxxuJgaXGsXs9e8URGlXA7jQ/fa16pB1wXkNKbdVWpEIaKuk2yvLLC9M0/11kicnsLkfj
wnJU8StrcnIS1kR2h5nNEvm3k5XuKRejcLXjgv/qRby9PdeuDv4nJOgZ2I60K6yx7ixCcEP7Ls6e
oKhq/SJ50h67mlY2AROQ6LXcvUE3zlAU6XJjTqACI7g/COkVswrx4xscOvs1MCCX9ZmlxGzibWfV
zYAt6o8cGYX9TCdv94UXyatBQMUy51i0YUk4Ad+0DcU03gip7omGF5wPvhexLSzMEvCaD5YxUPuk
cnET/2/wklXaBmF+jAbOc1Kmk03qPQKSi0x0Dl87GHSPLGwvFfLZnt0KqQRYR1wzYh9JXbsBjUdz
XuR/W9v1ihI7JABwLaZFVRqsSLNCjA3bqWHLI+z8MR2XcBwCLbgSXtu/XVk3As3uqLQoEHEM1XtG
ctt1+B9YUG2r1cCaW0kDVxUZamIKCoapx3Aeb3XlO0WRzcFNFO3UiaXQER8bqgSws4hFjAj+C5M2
D7wIiExC/1NlHPv09rMveLmwdxeeyCrJ3P/YpBBi/Jt4WM5QuGfTwqePRJu7Gn2OCZ6AnQ+aVeOn
V3GMLYBdgsNIAEz754yHiAYcwbLgHJ6tCkCBU2uDHtJJqe3fthBkiR9xKeRJ1FX2iFArlqzuzDub
V9w0wvK1Nam08WBVAGq/9dHGPEcfNXcLDxkmwUeCv8EJsSvlxaENgl4IXzDswOpSsrLv0ld6Kmcn
gziiwQ9QRwKmjJafp3KeXTo3jVHeeI5BIosAw43hHjxWen/2wtYbx/54KPr1pypuE3dFYQYaMYm2
zsGxnTc4dwKV6DcXW8iP5tRzpDPAZTQ830fwU/dwc+GAVPf21Qj7dzON/nzJcFC0lwD9O06fTJW6
e90XcgzgVsyz+xxzABfPPcVkE5CNu+NUZ1jCoMGv/o6mifTisj3sgZuZSY31fS41thksaoxBns8P
U4Vjytq4VIvRrMkuPVMJ3uSSOF4UJ9+i01bCtRTqLdlG6WRnDwg6NANMSklq1gi0fRCJu0OrU+4a
AmoTgPcrzMIokZNhLU9ngtxruA0UCyxlqTJeb0U/7uvdSCsIvdabuWPuo5nfG+TZnj2wqLhzjAT2
27KRWaxIMoxum2XZvz0bz9sP2gpU3yDdtbgnoy9PQ0ydyZRXSMqu4qDHIo0oU80qH38k0f9c/VWn
cWgVr6i0ZSkGVwA5fwO1EVbGPZ9r72KiI1PItv/893lCI0WPRgSMKGKiKHpLAG3RWEDOevJ0vBdY
KF2SujJ7pskn0irv6gY4tNm28kozIerT9lB+AduWrLiDE+FGDAb3Yiw11A0aPikScd20zu+ERYaX
iGYFVCGkWniJNhv/fg9rq8cFVVEf8fR/c4r6DOcKf5jIHz78IoobeQB+fNmCBqOl9eCkBEgk/EbT
aNO8JcpbzyTtZXvjrkpLHUr4U+aJFyDGtQu8hLiHNW/TukvEewkB7cbLvAGtK5ucDB+dTX2gb6kT
mvG5JfMLUYuen9WnfZYVS7k8SiRkcIL9XEZ1FDUQqay2rYWBwYsyOY98baUlzs6IuzUu3mkBea8N
yaYs9paR1lV0Q3HxbDGKAHQyv5w7uPkqL/Y381+O61rG62Tjbzut9uhy8CId1eIS8wr2lPcJ29/B
jaOwcLruDiVCtsGkv+d7XNnG3v8AJz7OyX16reSJo/89LwcxiPNxyB+RMNGNJdCTMKqXSgPUDyoM
S31nEbD+AdEPysoTg2oH+m9i5fnwENg355J/9Gz5zKz4xYtDqeiCxNMoNl+bsz2I8o5sGZUrfAhG
4stflNzUMdlgHY6YV+/nkfHHXGDNG0vM1K/Q1uIglYWhk8TsbxNaGZdSQj4SZin9y/Lo2Xi0Vf5L
86no+BHQZllghfUIQ2FxV4xzxKdvRgUkgeK3GxR2A+da6AkQwEO/CyXQhY6JUhYCgoC2bB2eyamy
li/zfGPQQf46eEMhKGCN0oO6YUBt5rB27SuzBKkGm3cBKJ1yhax1r1Hqdwq8x0oG84N7hwLzHL6y
kn+B7bob+9GXb7mgpwj7uQjx/1njDBaQoC2WQcyQQ3yFq1+plk2x6vJfj3Fo+vA/2SCK3LosjBCY
3h+S0A2qnQ7gt7us9epyDaAs07kkYgFRO1npM5UQj1VnZfQVuTdb79SyuutggcP0sGZzVQIqKjPt
MP/knQk/O3oSCOUv+ZDNL6IY0EBtUSMyN2LjHd3CevN/Z4tpJw64OOPRSrehQxGtEDlRBLKA0Ire
6utnjPTZU/TQsivQVrrgmrnswWVaf6TUE54l5MKAlUi8yQWyWOGRiqLOMOCOEwVL8sXtIrESBnN0
P58lwtoSrYF8nkADsZrxd1v3tCQQ6rVuu+bNjijskA2yqUeDyejXfkp7Qhvvu7e+GdyPeiSXSxhU
tqpMdt1mz+Mx9qUGI2L4AIkLakcBT57dMmrFLN+MFav2CEejtNMXXH5t2DGsmQvLUjX4ctJfhcfy
scfLpxnOJWVotAUgHKceHz3KoOs+yr1ifjQHnVdRzYrw3zeyJMQkZGX4U3kLD9QUU3PHnVoxczTQ
CVSP5kD+Ccv4j2uXKHgBBZsgG+US4afyfShZMSbK7B4u4Hi8Iy7yN36hwZNW4IRGqyRzAYoMhGiM
mhiCH2ZosjA98HHivkFknKLi32/Q2YxozVepA5uJtTH/Bnh1oKgdKG0KSm4BTUu3z8pLH5iDXYls
xK6RV14ldaIlw2maYBIcBrQi3oqBFILm0tTBV91QnzIjjD0Gn+KtAro60g32qFg00+ABUE69m6a6
EUDe4Tfr8OjqWONnHqWHRYRGa7TJm6DdHePalpnzKmDy+UhDxqC5LGeVkTywTq/pWllmFBpMblRs
y8WphmD5W671pjoYZ9gE0eknoxZDOEZyWy/tSavelFNCpOXsPlJqMjeOstiIaQVljZvW02rNyyFs
n45FFpRASR8NSGhOadc1JklN1pubwKQjYC33Ejj0spvbxhOFMHQtXE22r5hs58itQZCcbSzLy4i/
hgY5Rf3EEcfpJJEgyEvJyHWKkNPpHkhwoniAee5B3yLKlih0xT0SmDWRbCLi4NK1qTWIvLfei423
yEhl95Kb1QuPbBe8fT/0m97MPH8U1WfyfiQjkCgSTXM/v+aie7x7JOO8WDYYBaFIrUs4ERlgITT/
WqUajD83tegsXpUkggkTXrW8YQQ3PynYz2R7/nKZ55E3+p7GOQ9evwVlEDlRHHPxUGzatf9ZGvmK
0xs23IoiaMJJgr3lSP+iKvgLWAtNsgRUjGSatFMBsHnxKNHXgGZUHy1Sa+u8z5zB/35sOAAwPEex
7oKUepiehm3MnxsNMURQO0k28/2FUt5lKpCR/zacxrTvXrYXzT3eo3tOzEzaMLClo1S9RKKwO5US
XuqMO7ulJd6vTCpX8BmKFfVNaAahHY7mfKEGvG/jjI+R/49CLuTwyhX2VCbZ54drT3DCMWCzvjxT
wdpjprL69CcEGjjW1gJxKxXEurb8ax0QUgCAWgf2pBQMdOJRmL56sKy9Zy8VF55b/hqFLJPMp57C
mIRSdiAGd3OeOomoVEg5nLLTXPelE967Uv/wShgzn6Rv2dm2ChEVVqRMAuRXD43tG8lNjpJnnN0D
wM5NF40M3bUMphQKNMftbMfE/uYaxZ04u7wCLkbg89mnhlI87doiiokaQddsM8u2FcuW7cx/YK7+
4BaaYvtyr6/FY/83je686b2YsxWwmuTpTSvCI5P5bS1BurlaNGIsaO14fHmvuVXmvonvj7gwifO7
uYXr5CdASoCh+Va4icVhULD2G5NjsbOOe1vSbtoGqVc0NAlN6HZ+8MwsxoydDpCWjORZ09zSFCMi
flUpf0MzJ1G4phYGZUILlzcpFMnkbaXDnHeQzyPFZLgcCAssdYGF+KZLU7ns3Zywh8+MHuymGOKu
zW6WIYaguKUFPIWEF43HOJNmz/THEuQ0VgJ5IWJ9wt3WoClCpBRSq69zrUArcynSRKewFiLFyIE3
cEcrexlGdhYiO1AShn3fMGITdzkrX0fGIrDtVFa8Q5qa+eBVh0fu4ZqFVyTMdDYq5zsz0Ol6ny8N
ajvzufRYTa/q6vyVgUJ+kUvidAoZ0yj5Eyh3yVaSjxsWwjOjfqv1O/htrgnmcydaqNdGiHOAITal
VNnW17GRWyPPmMQ0cetP21ErpNP2VtO5qG5pbyf+H3V/a5jC1db6RoKstTJINhD64ftw/TekE56A
YLT11yUJofqYxr1b7mM18AsdQ7j/kVKdXkj2m+8Y8iKFu31jgwWb5bywPyjxnGGiyuLFoEhT+XWR
El8vjOLm3FW+SGAq9xeDds4K6blNr4dKhUqLhzlhwwNHRzyBL5KY0TEK3on0AJZJ7xckLi4XdQCO
5EbHbAoGBaRnsnTYK9cR9dQpJ8Qz5I6Ys+WDetH4rv2yEZ/Fr4VCOFxf81MzySv2yYOcEDK+S/Ap
elqEaC+Upx1WVAxJTumgGvhotJTlEmV3dnuN9UtdvFqiWEYvEMCiBMna6vX21YRMR3gvQpfMWJ6j
0osqUM+UYn0TYc+v9BzSTssWYyYEzcfCn2S7N9Bsrgleb7+lBO5eeavGZKqIWJqQM2TsKkA+PZrP
YkLLzTgTLKXU0G5mXd0Y2Qgzb/ipPjSsK/+ZpDlk/RbD1Hc5gmZoX4FCT5hZiV4YEWBIbSGn5KKL
rMdSL/A9tHY86+K1za6hbP2yxLCPNw3HcpWq9WCPTZbiMX0i71m9Mmz8BTko1evyVsrkQ9ERlU3P
lwCrvyCaCjwwye3B4Uq0PWqSYVVuFfHFTvS/0kuF4Lc4lJ9yO7gvc59EoC5N9QLpoT7Q4LkOKjGF
ty25Wjauw7jsq9v0+v0Gvsd//e1dMDyVDT6n1mfhchXWv/GEewIC5aKTnOWzsSW6e1DbsZxJWosL
1S59QfFVJoiORBdNWnvc1THVcHgu4E8pRMAepVx2J38OmwJ/uuBwBXCEbc8GvtoMYLNo70vAl52y
aC5nvglvZiL/Q8JtZ4rhjqquE/Qjm4dlQeDom8SegtpTnohysPWamEEZdHY1PzAWNtH7TZkXLfJL
DR/3k75ltWkAQSFAAxIbltRCqADM93VZhCZNXHHaR5HWnBd0bOAqF2y2F3pHDjGPQOz78fms474+
3rCZUVQk2u5qgVmBkH2biitsl0cnebkeCSGtFz8pj3ZSzTk7dd3Vsvs08yxBSCf/Wau5tVR682Dx
IoAwY7jVnFnji1ntLO/A1bMlnJsPrGF9Wp+0uj1FC84tmzCXWclzynphiIhOaqEUqp442ekaMYz6
Id8EQnrD9KjgiibrCyPEfnne4Z8valcmZozWu+TuHEw3t0VsAGv9Mj9NGJXYRaRz7VoMDmOtqGVk
3a4XwYX6f2pDdU7J1W2E8djiEwDLoIuulvZLN0BvGHhjuhyYs12Ol8H+X1JsM+4SCDQ2YyhqGbcT
kg8JXGy+LVwtBX2AAhUJiE678oysZ0nVU+vW3n6FuYTkRgTpGe48E2G24LeP8lxSZJ8nVdNVDee5
MYfR5IM1v8G0EaoFYjbbJORpym+uslhCouB3FePP2N/ffG7bEcCJb+LiyOUdxfPLg7FkvQG5rAzq
cNUxlPfB7+l5IU+jPDhCQGV7CEx5C+v2whOEYsYsdLT6lWo7fbrmyRNiQ4YRmABTD+Xj3XG7X8Dp
qyslvvMxx03rSpxT4eo6ulA5AD09VpzAEvkWosBud8sEvDlCtzk5ZrxREX6wT2vFxA2ko0WlZi6m
GRcxmCDpCHmzao9yqd069X4fbYYXkVV05lRYllSYEnAJVbdWMpEb/a0ooV2dmg98EXE/SGhaqI/h
bXwO2tpCSj1IFV5GdbkckOr3BgxrqSbIYG5hnU7PDnofkP+ywGZl3vV4iEOmBTBOPKV3+bqwxlgr
d6bBCn9BwvUCJyZkk8T8X5plaMoUz7aFZ6PN6/j7ONZiX35HFmZxnvOQ5WjzWUPG4SkrfmMCPZam
ZhI5FLMlrwhVBCpEXEgMJdA2EXS2pslnheJXQGCnQnWh2sJbSk+2RmQ9L6MCMhebrfJBuz6FvzZU
L29JB2/nuFPMVRJntSR2WezMIvZE1DG949MInkwOAKqbY7PhAsRGW/M1/nLlZqHFlWN0bTtTeTqV
x6aNOUf0cYkaOIHLlCSxjifh1w9wmOqsNmO2Gj79zIoTt1oYBuIYUj7LEsyZyIBnGvquOBy/7Lni
BMzEp7sVtbyUlgq8wKmWMJLRM9oS1rgz06Mu8/NvJtXN8f3UFk3pok5dWkwPaGER3zUIhy8v8+4b
IkBjp39VOCxkv8Vw4jDJFFwzzKbgwdkpxkZ2eNa9Kqv9CiOm3g2AOw1CaQpsZpmLgF2xsRB2yWm9
kQE3b5TsLO7rA6YH3vZO2KenWqTglf4WOLkyZwWS++jEgbopFuUpeuHDNiKukd94IEK/1qhIeCxC
y+qOXEpKaaUNVPzwsygOgbArElT9bW2XG0sorqeeDDTwoRA7EUh7rEABsyzFFScxMp00GCF3m4UR
+bHgblaem72HjGDkph3i0EnmvjOVx1Zd8OKhTkOhkbPIZUK29yU8kYA0BwphG1aHrBP9JotusiBZ
hEQ3h+5X92vHYd/nLPoBKZR1peddzeYN6L2pvSCqL3cBwp1czm5uYKQO4odK82ULzSDWQdB+5TdP
MMjENk5P+SW85Wb0YLbxKaV28SJ7GJ3gCDISw2btpVNLm2OxaehI3JHc14z1HjxdRYzz5f/t0imh
bm84IgIn9pTRy0+x4NSi1gkMPQiWOXYy5v7LTTAEHFigfCdfiAvBRNh+li/QifJ0DLB7KMSfITfv
r/ZYR57OQcyXREFiWvmGRxMUaLBWAjkvREdLpNR3Ghu06Cqz2Hkc8L4d9rGb647QGXEv2xJdGV+i
2mrPJtiBzcD5M2EMYJ6s7mXpl+zh1VVG+h7J6kBrwtQ8nPpyxDExTkSMItVw6CYjPeZxBEeiNY9m
Wi3TRz1WiJBy/n9AFAfpcQLMp/vjbj9tmcFzmBi8iV3xG6NwfUFqcKMVLihg6gVlcTExk6XaGlDk
pPSNZWbvrVrhMR8zliqqynn2xk0gw4iUe+odghYeUtSDg4rqoSLyJ8U/QmbrcxXzoKDo4buI1Mvx
cBMPshQnLupq9KaeoOv2+3gnLStBtGPyW8oXHXjy9ciJUyp2+uRUakzP99YAic1DDqSrf3/Un1U8
kM24dL4Hj0cot6JqbRaXPzy6Mo6/vyQ/zN0wh2DZ7HICCS2l05jEUf07Ywkc1NtKInz588W4yVin
xQufvggWFdbOzCyCVCA4ynlRP8dhDBRRuakxNMQfDJ8SaUlzwYIWWGpP8QmZ9wFZVdww2QfFnUbk
UeTa9EFaXqVuTsoSHRWj8clKac612qVOc50Ll9c5PNBA7Id6Urc7XZqQOT5H7lY2zUla64W+5uyJ
h6UwfQoILHXGSwYFKgF5pzeyj/lEebjzRULY7tczluqvJEKwPB9gj7VflO94Llj15jEFE2f+f3gJ
1K08l0W7HewjY9h92Xvh6J4mLurinM13b5glu1YxH6IRnaHoSOXysV5O44hwBY1bJU9GeH75BQ+I
h9EtES3RhzzVDdGItLQLfKZJ/fxiJBR7GtElLvYPfuCP+mTDsaRfUxSise6cj8JUqDHybZZMAIBR
yPitJPMbOsY8NhUO+kI5BlZU6XQi7AupEFvRKPTJzm6HMnBuRp2uF+L7eXzydp+vclokOLjLT8Um
sps4C+hduo1lmVHn1r1kYT9KWvRKrXT6MBexOGN87yq7SRLPl96lqlVHjMP2Czks9BymMlIdXqxg
GVHyqxUQUHSiU1ST2xzHBCB6oN0Ygdx5QaT1zCkBnL+KF6AI/ZEv7aD9A9O1q5NPpGIgbbrshsSd
FKoF6wIG+cj3QBRUOa4BGJpPsPUxwhHrpHqRI1nEJx61NQZX/64IAg+NIftu2tluDM4ExAwiCheY
F0AHRaFgXdIeQriW4jVcCqpRe/H05yqcLtavKDTep7Sj1sJqISBWhEAdfSxfaOJrKoGDDU7DuY2m
3nNrUrPZbpqkjO3PvNpa/sSrbEZlpqx39fCtJSJeSoXjmscDoSQCht36PbjNVK15LVC/oVUnw8Er
cGxvvPGIuRSc6LI9rZb48PMPXt9CG6dFvGHMBsbNob+XDVlQrHZKp53R902oMZONIvXzn/U2Qcec
pl5dY1mRHAKt4oBsan+E1NzsNHrpCpQ8ipOfYA/SEoCHVzQQEF+Nq/RJke9lgthoonu7kUfeV9Uj
ZWHtrgaZkaCucXTXs8gPRZoVPah/SVCu/LgX+mFP9XLsYmqgEcdz5aGQXxcEZCKwVxCoio6l+M2L
NwgysXgex9Tp4Bc9KNnu42QBfgM7iU21erjGkyNCZWMHOYdbw0pA+8Foqho1nulED/G6BmZR4TlF
tn0HwHltjy9xW/ZKhOKDhcBStoqSiE4opQSI87deds4D0iuTUNIw1rReYAGDjA4Z7l92r7HfGQ42
QHwMIAUPIMiuVZ4wLIXBX7A/pnzHrKrIaiZjhZLYPs5E1AIJb5s7sIQCcokVfzJMumN48qtNBTbk
QcSaAn5t+23VBSS4Yc1x1x1qhsknsSR6hTOPPa5ll+7ie39t3tFOjfDPfolXgsQ5W8fneWNbIps9
24Hf13eh45AFYFZujC9A4FKRRgN4ePi++lluKQhGiK0NfpzZGM1EdfNdRMtwTKm9nAvP0RPt1eHx
ZeLigly/aUq7Ez81vSnvD7yOBiomtvgcX2J4cG05IyKu5DXo0FWXJo/ErfrBG6FAbeb1LzoK7Lg1
IPNP7Z0RKjUP0aTe15hCWM9sDAArFVK2006EM8HUA30Zge4vSngw/JTRCIMcYy4WrQnaeMRImynj
2gxLgZjpbVLTJyyoUR4HK+qwgNQ8poxHi1heYPaAD9KnAkycbPYELMzVrPK/Yi05r13Wspvo/LMs
1/yS+Pe6HOPpA2Bu+Jw91s/KvaRBt5wy/BfdIe7Ob096QZ+4eoSfbFaNyu8SJtb+r2bvbrphsZvO
eHSyIiqbf1AWcDMQmHQQxvcR4Lzda9IkL/P1SqrqbkqYkzpgzmkoy48cqg98/m6am8f3zKPkGHhn
PYAIiZbsPkhKRoSXJPmm23cl40laszoMMkKjzCb8GdU5y2QOILMMi6FPhi0ciUaUGY+Na3t/DeHU
rIniKe+osvWHtZkOJ69m7TmMS0Xg4AOGZyxpiVsoYnaf+QLZRbZJJoTxHUzrWMKGkDemzzcysFIS
U5x3kc2NJNbHEfepaW6TuT7fcHQsjG5S/VTq3wnZzvSiAeCauaUZU5RSQG/WLSvXPTXz7uMAwGjW
kkAmB70bwto8wRp83hywSUIPBI2YRH4eDI1gOulBgKxb4YagQXQFR/9Ua7lYd7yz5f4ho+GTfPbV
NK2+UHs8j8C6h/fG4deIKRPKsoSt3RcQugKFZ/vBBmWIy2v5mp8cdAbouaaAy4DxcY+/jSInl6ct
HNk9sQk7mOiktVhnlzXeiv/UYSU9pwt5hRd+4Hp/adMAt8zDMWqYgSfwO3zbfJkRCTJv3g20jIde
youhdxQi4DmKlF7tkZRUXU58gzSS4svzQwd8NSm0MubbuCSoNoH5ssi610INJlOGSYEPyhQYsH+2
IciawV0DjFjqgUsLfjvHe5j2Ji+fPxiSxdxeYwge+UoLDI0Xp39MR0lNvnthFARfQFQRo75crp8z
yfQVpxi9YYAJpc/ta+Hy0Q5B3hxQPecPDXAvepWf9zNeGzKpuRDCO2jb0H7okgnHBQyEOlhjnjga
wI/wN9paYBWFXcXBZwBYuNRdixgHeimt7VW/IwbqtCf9zPW1+coD7ZxEk9l9DNQiKhJ6v5Ctz50o
RN5YPPSoRKoZ4NwpvJ1Kco6RCzKJTkT+ZcYLOttbK0cmXhgtsuX+YQ5PDQ7V8Gwb7b8V9ZnWQDbk
zzQr4pBQ+GcwrhKPCqFY4QlZfqjPh3Be9v8oSMKBB/yUG4DVdAsm4JFKfRU81q3dG+XLwtMLImpN
0PwaNe8aVJ0oqinpVMtfaqLL1s83UxyJaWA30/1lG/Dtvfv/8+8dtZfjVGJqJ1pijcW8jro/a3rH
XXq5Ww5O30dD0Ohqitx5ykCos7Fue22h34z/lw9RSIAhC7b9M2Djzm2OJqwp6r9kWtI/LM7plsob
0oMqunbr8/DllIxBngKj5vSc0BUmQb8tM3vRhQWNSQIZ+a8ZJJMY1sg8FoROEhZKoN2qMPHijZkK
9p1k1DPOauzsTLp53SMvRBXoods4NnVFV9XacHireSNsjh4DRiMAZ+ehy7DNf5JI5cQA5m6wU9bI
+YOLMjrhd282B1yqzCreUJvclLaywz2RTZd7sL5N8hhPa9EqJa3UAvCc8wXxqWbYcuL9pAu6iqd8
8A05X4nLm6GyvxPSGdZzzm1eCY88n3F0jyejrrvDUERDmN86oMYkIyrBGe0ifpbTAEWXVEndIEse
j3UcmCYpyktJIrVTY51gmeJCQVvdOXpeZ7M7HCvI4imwA2BJTvDnvAcs132NHspgJan4XCW6KQBp
R9K3CeY4pT5krEKOAtipfeVxxTo82UIL366tVUUaIBGS4pEJ0TSkSdBHR6AYA+tEQCVez25iVrj5
zAfBGteVJdCMWCqvc9VaW4ExagAcPPc47r3s2GbWlxiWEWjsSeBe4GtV9pBiKRvV31ETAhiCw9CV
OE+AUH2uhNXEqG2LLV0j2H1QPBAntYVqNWhSdQEFUOk/smeyO6t0ZOY1phau4t1tOe8wiSlb70PF
gsd7IZFIRRGmaesOZtNdAXUZMOdEioJuAQbHdn79n87ah9z3Tgs1GQvycxgml9Scszp0n6BQ61XW
bpsQV6qxe1OToDxrnkVejD4vnApE2XbJmLjQrCbYvLth9Lhf7v25qCHj/wepMCDDXN9K9pPQcQjd
GLj48XMse5DL/WpJl54sG6nxCTka5K07Pobfdm+IUBZR+aTIqxWLWyFSihrbXOVPcCpIvKv0psjl
aVLithE28uDcEvXcAWTdaeamz/3bbuPIhP67vuzb937hopXEJAYzfDOx6RFgpmKyoBHv4fnN/igR
wohHD+3yXYoPySFHfmjNtRe1sjx5SZoaPSKFdjIOUDEniz+FL75rHKGYUZ//wq7LMC1//JGrZY9o
qWL8USg5zwU9RrKTUi8iyNgzCco3PNZ0Zc31AGrLmLARmOgXFSftuFags2z7lv/WBW/PrA4H7WaY
eI7AB/DImdVNfM0R+KSe7jVFahlINXICRMvwtJ72q/IvBuvOnit4LwBRiYIDNU7cNBwW+p8Hyvmx
JNDH7d2oj2sBBD5yYWIcZ/7c9KffvUFvxqcVQuKdCIpkWQ3gxYBeaHA6DhjVZ/LTU3z2dh5PbU8E
nREaiTMGY9bRTOOwCbX6X97vwSluPTyqdaRsXz1XXILy7xOexWDN6EvwRsK7VLQGPaUHpmCv/PnU
Vxmbo3KlHGNSUpN6f31PGdiKOheRbaqNorMOb2FrRU7neJfD0G+ZP0N5KcDoFl3QLjKY/HpmXO29
T72LBawaV2pz91R3/0VQiAapWOTx5+2nH5cuNSXIDpPIA0nkbOFBQUB51Mg4HZc/caaPnDPEXsFQ
Vrme8b+Qu8BwBvoZfU3jyL4oU4TH9zvJCDnn3wrKU1mQVqlCuSKsAXpgrLzNHR/c8yWelBqVr/J3
uG20UbgO3N4u7nDn46Vz8oAuMHoMGexGBrIlQhzBZzMa7ACfMi3uU6X1+weAo5tCXk+2P4k2BqIE
UFnoCUbIUAP42NAI6g3Ztr5fsD4wKeMFNk4r5nX8h0Q0XvGqgrxHxoBxr3PNDlxihu+R8l2FuRA5
ZyU+Xu0tlVwv0JSx0qGABgc7xhcwjm4GAfWGIjQltgeKpRyR6sNLEVEmHRzzHIy/pvwAF/YlCSge
A7mEbo9+9++INA4HJdSNkyry8bmDjyICTk/kYcg3JCGAUR1/a9Bfb4UwCUHZis4SMJCUBbn/T/HA
wYXtuMLomC0xo7wsx7xF7Cru/LucJBFMu2PLOzIjqSZrgFaXMYru2pAkEZhwIBf90p9Tzbdv77VD
I3v6J9MsXQpbCSHsNrLCZtcf8THXqGsxELhzQYL6tCskoRzEbnUQcLh8qoErXYtHefGz2HumudD9
/YiRE6ORGs2wd82PFEi18302gxkRJ4CLy99DI7a0svVt997Sz1T+vWfaSgUXDbyrn+J8nOUTREIN
0zS0HtDhHW20uEh/aiB5RyE9dvXtGQnTgHX4d0xw8p075J21elgEZeA2CG+sJ4YvssUifSn3UZXx
D2yqfU73OmtgIycBseOJGb3ACzNHqtg28Jo3EAmb3utzb5NwCoihvPYG06GoDs3johIL9jxIoj5E
VcvYDbW6hcF6no0nhd9CwXKMHR1MZkTzOCK5BKMsGiiTipO/exb8WpoEJE+3omu40qiIDlvrtO9S
1WNuOD7dvWz/DdLY19YcD8yS4H+spMiRd/oazJkGnxCMilxqDNFwpMsgnUVDHgePfyj27zccPwhm
Ksm4ZrXhtY2lC7eXvCB/WYMtugGWX480/2bE0k6Ipc/n0wRMwTkr1yLxPqYgs6SGeptGMm0S0k1Y
JBxByAREHSF44r0s0csgBOz/m+AUX86rxygsYRotHV342rNpjW/Ihjl9qeXsqIgDpny/f1WwQIAD
n+T0g5Lh8cg0WGWkjltt+T3zS+dbwnPkXf8tFVBg/SA6hnM7uzai2N8oxde0z388ejMWx/ZWXVFg
2/8uYNcteSzTJpFrmeqWFmibb3PEwsxLSQm4IRZVamjXW1osVviC7ZiDPaKcWFKuE/faQ1T5mkzh
YzeDPbwg4jCGHE573L7yorj7J76Docs2bEqQ4eieCEQPXHZnoKLdO2MlJBBn02vxAQYaJ2CEqnOQ
GQ4bV7c8W4zOOYwA0l6JrEzzNzD1yxTm8Zk2JzASgVvkTN811X02YC9uB9GjshgnqPVsuqsKlxTt
lAA1WCnWmTFmiLY9IvVG1coOIiJg0H90FmLuqF9C+ofUdK18qgzAFXyA/Ft95hw6zezgURsqkIm2
ROhAWDlAZM+3I6zV0yCLijXVthL8mE5XdIrvENCZvLZr4MmzIOQRM+3m1xqd4S2PwhLkpWxKJq8J
Q6z8tFHM6R2kHK0PsJP9VrdH+xjT0a6WWQU67i0/1nwIKobmwpz4cSyL0I1HSr1yvK81alESzMrQ
iP3MLChCrWIkiZ5kR6L8ZMlx2Oxbr7zGvebb9YCJzlY/yc8mPJSRAmiwQQ6SLECBrHeiwBjhNnLm
GCX2lUpjMmYwyck3RJVBcLLJ1S3/221aSImu3GEDjCFMndlXrOBQ6SWRtRqouZlLMYQKT4AcTP9l
iSkl59UIVq9IqO//dMxNn8qWvFvCcyVbdLM6xEr3QsVQLJXsMZcSIBPog6WdyqyMAKCwMBvDO7Dk
xOduPEpFmPo+0ShYAgVvkGRm3a/CBdsavijb5uy087BmKGWX+2F8b+9pRMNW7DoWBDIsFbpy6jh2
ocd6MhrQEuwHJG7Knf2LuECTx7b5ftH1gw0lf357I8n1hg48+1Q0qtTiiaWIeAOcoInaogK4q5dX
2MnFhkO4kvgabDUTyXrSkDP5cM0xl36HrvlR+vT4HduaMHLiPHzuIab+DyPNmzxwi9ohk2h9VM44
WW189GwdM6249psHtlRCgwASn3Z1AbVxAxdV6JJbF2yVkbX7EWo6TkEYU30dodTxEdngrZf6HUvn
ewkq8hqIttdEyUiFazA952xgi6FJwnQ1OkPAqRnFAuOg/iO3epy/usOr4mryUt2hL4Pz2g0m73GG
DdfJBgtp231rxYTSTJF0aOMJfgplmSzncWfepmAFPO2o4OpqLtUiyBwJiO846+EQsKdTJORnEvoJ
/3yiv7Bw0t9YSDwB+Vh2yafxZp0KeSVF3+7Q8cyy3ztDp090wDNfVcdFV+XE0HQHgq576mtUdLYv
k2tMoR1uidYSbznxZRx0cJ3MBqClq5ukJ0cgMDC7Fm5QNsFMAkPHFxIHnz9VtA022ZoIR0cOKBrN
UhDc1ot1BHhTZ8lZ8Y1NCFtAzxj3wtuP7hMmVCz4FzG3qJFJvBA4CxZaUtg4g6XU+I35pE1epLak
vZEwsuE7ioHin459aNOkkB43DimYCITw6YodWwcGGtAG9XW6AJ4G/cCv/r1CLHgpJkRaaxeMqRF4
3ICS1p717Vn7nTzk14+hJfhLvjQwiKFbdUCTuqr34aTRnvj1Ft3s94PdEO+w9m+IG5vV/dwUB3bp
oaKyB34VYD9Vdgg1iQqi3vvIdnJUs06bkyaR6wik92KStea7TEhsVkAL6hBQJDJZifqa4/QmGnoh
aYsyTOIRnxxSCoFXvaEbJEMchklMrz6QZDCeizWA6sedIe3qA+PggK52cFgQR/GuHy4cQHCFCnnK
BtquGX2scNJ5VsdMo7shVr4HOgBuPTMskGajJI6QIo+Fha4irYi3ZbGBAY+7A1vkw+pTBJKJkY1L
WrMsATN/IAEqybOOEKMDnqvEpOWQBhI2SGazlTiSC7ioR9nXFn311eagd05hxRC2mlRFaSX30K2s
WRdS27inAfvh5hkkRb6rGSPCo8r065APNcDyDKL/tii8zyrqSyVmJ9oKb3iyWQh+2xke5lgrqB3k
lYmp2/t4ubpcUDRh1wpkgeU0NTUKR14VQVDX8urG8w6h5+wuyidasB1QPGn30Yvrf8u4dvnRH270
DPlOUmAFYBx+dA/7wnSOY4bdTpQN8CIzWhrQL1sWvmUuVm8XEWJCfAb+BUf6Xr6k9pInuURTI5EP
XUQSomNxSHewkQAWFi1PoC1wWG5PXUVHBLEMahdpRh9w2gGNu4UUGe8PKT0YsnAcV0RqMp9Sk5Jo
SI8sQkG2XjEOUxw6fG3oUQA3F7Ms4C/FqdA2BzUI6obM8vwNwJay/srfYu/ysJZq0Y5jfVjxUYqx
Gy+E8uBod0RjrsSEIMt9yPVDIvTBpyNIypTQcXnFNKtCa6N+nbMTgoEptXTHRHc4+g6gDuPSPpel
q2Qgd6aVkgYjEEjnPSOrFnC/9oHyKRYF7LV7dghPlPm9UzOaASo3k7nC78RT0+Ox+WX/YAra/7jZ
ium0ii2hpl6qIMPFRkAFTJEj4SVakmaDAYMOuQre1/P1L1MCihQq0DrWQPupJMKVdgOy9Rg2YaoV
CsSvSOVOMHcdl2V6x+K8H0qdhMFx7PU/k27p1U4poHZwBV0TSHjgGSGfrbMdJgYTN5xMjQPCoEaj
WkSwutBlC9075ZeyuoacqEXAE6XLhNMY80DlPBfSD1zruwLBxOfBpmnnRi9t8+Wu6FKQsTfH+ksG
83eWqSQDBoJZnL0EoMN/ngZ8m/vE07K1MdDEi0JhEZLI5xDYvvJAjIpEr9rLhSXdJdj0S57e/GaE
OrY+LP09yUtEvoP1A4+b0bbTUyRr2TSmCgP8uBIN2quFGZsLGE2g549faBCwm8c4GACoebD++OuS
nTMyVGJSnggMy5iO8MUSK+TO/uxioAZRi7azGek7LlS9MONJ10QvF7aetRJqlBUCRfoR7nbXQ1Kj
4Ocrn9DuMzVtbrIctf1wU8bZcQFRi/2hbyTYThvCne6V2iVtg9O/c9LqVuwShw7aV7qphMjJzgCg
yQnvLH7tMx6j7peQHWDFiHQcKcTH++tc9Kz8YYo7dknYyedCY82TZuU+miiqRgf7102x1KuSo8Ty
rm2WQihhMnihG6q37nl/OV3uVDCt8a3Nes/KX3wareFoyo/JHTmDlXbpJ6DDXaIODxh7VjN7HmKZ
b7HN895swRWkmoGHmDGiC9knWYBeeNrvhbiqy/QDYnU1KJYeO2erITI2nyTHH8fQsLT6ib6QBLtP
urw2j/gfCPYstv1YpSL3Sa/LmqKd6w/eizbtmcTTmrCgOOVImg6svk8eUSu7t6gTLQMSY5FOu0Sj
QSYFeviJyF1XPmLzWd2C15fa16aP72KMcDAM2Vk8Oz6ZddCoJk3EKKFCOvPHzZOX0M8DdMChH6Gu
Xv8wuiZBeaC8kmRxkPgVCUm/GMRxOC9ZNXssL+WOC6igrDHeK/wbcjwjPt966hTcWYQcBrZM54PY
j0BaUfJTWeoO/g1ANJygf2ilKIByOd3EgsaXHiYkejwWcrmRURul8Va/sdhqB690ADxRwV20+8Jf
xdZziL0ShHIo7XLPAoC0zMKXO2tP2z3lcDIiecsJTXrFLj1FL9SPqxc01tuvoNWu6bhlQEh+SyhZ
Ev+kR36nz4dO9Sad3e9O7ZNh0+0rMuCNhpSwxHc8jyWbryn4Z7SL/uMew1DetNS7QL+HE7Jo0Tkw
oii3dCxfbxmq1aUcsCDg/4dKQY8LT+gxuhH4EJPs7VVtSOJxLnI/9a5X1ayp4LlfRXzkILGlgvOH
2fHdUEgg2nq0Muju0auPtLvgQBjS/PjgUMLLOSAWy4Z8odAhZQCKR16/X+K+0/upav5tXksoApNe
m01b3eH9nGnenwZAm6kt2qlqoHZnKNmlRI7J/uxkueu/vQW800sEUN2ilWuPYnZf3oaWl9npQdB3
Ax59ill6mkbUZNO+z3OlqCCwzx1wiG9eaUEH66j/2A2DE3cMTqkRoBcRQ9km75ph+o1TssHRpAfv
qVMcr4TEyC7WmRpuaFSbqAuyUz70DW+WXs6mfYAKD0Ld27ctfDjH5X9e/hUrLUIRQRvMZ6gEjgaM
fcd5zMKsYcsefO8P1L12tTWRTD/zp2PRZw7RNexeQuRBN+YLiHCIv5wx0yy/nbHGOWNNb9c9hQTw
zaGDie9oLx6Th4EhuWRsLEIURk+WHdTYz30EI5kQ2aWgUy4fwiyV/jVkUmhQIFABrbgjl3rgP9SF
sH0IUwMoJwV3GPaiIY0Tkfq1MeKk0VLt+krXAd5bPhcHQHhzGjYzXbU2XPRHTlENHfTw0ksqXElo
Dly1qZsWqgKC9VGW58ZENr7szMF5M4MOB4mJ27UjTD09OLRzJk2WyYbHclCYvE8WmZfUIGtRBjDG
+BA4oDBU1i+Ux6pnROnZSCg6D8pyAC0vb0ZKyeBH1WggICmyEHl9+Ie7Hsh0pyMwV/gTTXzoqsFN
eZjosQQLOciOoBock33vIw8eBudwTj8Tlo9Mq9279VdtZisepDQhJLvtyvXIkl3aV775z2WbxjKM
YZqdWQ20DEnnCyy5XfstjlhQLdUJ/8tfKXAvCSwCI88EEmQ7NG+G7y1i6pTM10C0FsRxgel+kAtY
4suXALHpg1ciAwHxSgE/cl6SveZvur/ha0pqPsSbOo8eATeA8ZK3PDATS1meW/CEwc1PBLShjwUv
pQtFC4tAIkUjimuKuoiExFFOMT7sKoDVH+Y15qLdYWqLB6T3N7tEWdlJsMvWM060wAZmj0VFH0id
cExU5lBmGs2a9qV2KPtNEXH9uCc1Oss8b0mli2tV4E3a28LCoZae3/H8FY9THpg1vrMwy1G1flcu
8VoqOsjV+R8a6hCclK/brSEuF+cb27iSDIIkWdEDGIoMsHlhbzWMRlsvZO+8+2OScoo3Y6aleUfW
X0FdsyvCQfvvpQljOBtWo+mgJSTBxQjiCmpiByHtRroTloZq/jmyTfDWbf5O0LWXt6pyfPjWzolA
pBCwxegIdJQaQOlbCXDUXsgt4Vx0dkq2U9Q/jlLIO9zOf3xc2t8sDe6Vyj90I5d0rLYXwABa21he
4BR3n/t1jr9cIS4baDsLChHHCV6W2yN6KXQXHB820HW3k3LyT6JyHIYPxfx5RCJvjcdUxXGUejJT
/GQJcXQ0HAfMLvknXyMJTw+lVpWGsebI7fUy7i2msGJyoid0hCjZ3KPrXMVHgQzXnD6v+e2cEoZu
atmGZbsc3+r1CFEueasoOHN0SCHKwFdtr7Gr0mqKLhnBX9dEpFWZIiNjGaBGeMCs6/7QvfStrDlb
o2JAj7nFPyyuCk35aB6SS9OWrYrc00y6J92AObnJLZamEKiQWnZVdYJh84gLmqyn5EyYgv4/XeiT
1aXPggUlxi4l/lbs9s2lacw9bHw/nAYOGbbT10ijlKzPb7KJ5jRiFXlEoV8fW0SAnkgEr6xB08rd
jxYHmsE+uDnHp4vRG51b+Zkh8ND5+RcYXi+3hS5u79Z2mYWRFbqmPFID0Vo1fVk9GNWFdxDib0hi
CKWmPZL4MPT056g4TmoWew9HycP4FAFnoc2H6OoiPCg0Jo/6JTixlUWV189J7T4dCcZKXjkznZy0
zDIAJXP0574GcIxk5STJQNh6lxPNayknhaXo8Pjs0R0b0giKp73xpnWMS7bZPhJTNQFMtGpUVXhi
JEMADXCIVjJk0Ex4PlhEI/9Kz13+OrAD+tGTYGr8+RuUq3BArFQmEmnwQVjuw0oW+urtweKWDmUq
EDboCbX+uOH8yTDMFU/NHSZUix0oJLgPBRIqgQnfAZgJKp4sqMJr3TQ6IEi4mCAavfK50q8owzT4
ZnQ9qIxWIJCSaj7GRIjXcfew0QK5vhZC1CkHnq/etTCDJrT/lBUl5orrh7dQ2k6pZU9nkTwX5WJt
Ry3SmkDS9+aGlTM2JbKRrhQP78u8TMCxEHSd+nxwPER2UDlyOdAHqlZU6aOeWkSqQAfwp7wBL8JY
97mHTDpHRUqvHdw+s80WIuc/Uu5ORkJEtBWfZ3D0uwlJD5iKCmFdotdk3xSfYB6GYMMMBoi2OQWR
/unTCfNYzJglfEZfYvfsd6eq5TnjHsoBJJMbX3+0CzcxF4Ia3bH6d+yFHv3OIpKju5tppAWafjK8
TbAyZ45KYob2x+LUlKnJdBjGXlrRFSLHnEB06xBaLClp7TRT5SskdQurnzjwF4jcu54hYKSf7vdO
5oAYJTGZJRf42oajRMATPx6vlOHXB5uOexpH2hi8Mdm9ZMxqkH8CnvPP0/HLctneJNLTBmpNX/CF
SUQApoW4EfIJ9pnTv8RqWvVk5VN1tnEirbKwruhGRG8c2CHoz2ujXmxgEAOjgjh+cNdNHQ1vBx6W
1rOWuRMNMxpnU1jdQhNnBWTTJrsJsKZJNMktygwflg/unSMIeX8KpSt6qGi9pkCR9sMQUWk3zajA
tGPDBBeB7bLq86WQJYtErnGrgcV1H+C+qAsFjGgHpBtdU7DnWI164s6PDY6AUHRKhsDX5etCokt2
0roK3exs2CgsJLpfMPxOoknVIbm2L18C980aLO16EBJ88Wtd8wAm25SVZfH6iWcUXSxLTsBuPRb+
+49X4Bggezdg2jkrQrV+cGr+BIzIw0ZfItyoxB1oM6jutwTT3sxVT+mz6uzxhYO8cMdAB3jvNv2s
aw35HjRiVsU+Qlj/vGmFxPtZRrBX6zHj40DQOVGoOlawbmlsQtv9dtnrB++Bcdzqw00V4I7NmOhY
GJYtvy9cUvuEALFuzlv4PnZ1CjPnlxFTv5VJ4aoiq+5Vx78RPcmU6sB9otYEXBrh2fyPtBzK6u1D
VnJaSol5gadvUzr08eu04r6FG5frjedrocc6T6N1mJTGCqZRUCfRuD/WX05PR9qSs3EKkXfJMbIH
ExA1OiHfFCcyOlk2mOrDlphN/fo7uBjtHANdmOJisHNcLPrYaZ7zmjoH72zguhaNpOfcycacqR95
OFFOLGcgdK6150PqmhbRqMvj4zLhcKlpClF/4CGNoRiClwRdL9pUPtdstjh5ahfctAHQ947rpuRK
JLZFL2Ur38DxHBzulinAzpg8MyuV465y0Q/z1lPk9drQ7rvmUIXRLY2gv1i7+TlN/DiUh50LTbH+
pktZnH0mqWz+Sg2YzjM/EON4HGLAPOOkn+7YByP0Wet3126+J4IAW9WAxMmyDSg+e+/7+cfAgZY1
i/XPnH34rQxhTnD6DDSQ+ADXEAh06NLkwq1Mj8pr7D1gYMWpsfEiZGG32oyxJZSk0o5szRS7GdEV
9/5T0grbfG/Ad1ehpdoxNWpu8Hwg+y/HZubYgQdKFtlmmgVKN6OTy+Ol1+9Vva0ypS9ak3ivoBQN
FPZZJDjxDx+K1KdPya8DL64jZZ2Y1FR6my1/L61zPhUxlEzdKyF/xOO9NzsEnwZr6zT8OV3g0jwi
lZmnPWuwG2RlaTilwqrOi42gUm5+Jwz/8R1S6ZcMA8a7w+QXzDAhAqbncawSnbhOo93/4n0LISzX
qUZHHbG2PX9LccD78Y43bs2DuWvEgDorfgjAdunshYZFNaOKtOUgeEzaJ+pvojkalJ76V1xAL9AU
LRdwZBWiUiQQBzVPcir6BkjDKHqyEIttZad98IbwOtxDaAga0cO1S8UaVs2cKXTIV/2SgcZdEb8M
6KR7jxc76hhKrn/TZTG0Es6dsFRLLn83fh/oOlFDHolfacZOs0/0zQ6r9SS67RQJ4nUgZ6ukFnyv
J5TbB8x0OFK6eOCnLsfEYLEMluQmT9tPFqVuWZtE+OE9F26YMGPJXG6ivxia8ZvXMqy00/D/Kx0n
30boYJv89+5oSAQ+Nj7i3+3EqAFGlY4YXxSXCuMrpqkMIgJUfVeERZj4fhvsd7sAh8CHIRW85F8l
+pHYPaxmH2SmBYhsGcm13dSkrk6EfBGnTX6jXAdMdCvSiHdkSKuqjfDosMoP1jO+6HZKJVzl0s/L
icRlbzFhbF+SIWc6JN1Pk3U4ySCkfzGbNpqxGMIeEZKF9AnpSkU1FVA7m+FutwVI8eEzrZHM5lCo
6EbxDIdnGy2/cuzX5lh8Ezr3Ahzos30bjlSN1bH2AAH+moOCKchuVeIbC3LOZKdS9mU55XgazPeH
d0xvDMRwRIN5Q43xEMB/oMGoApCQIGMuqiDXRW6Sx8PtnG825uTGFkGUnngkDmfO6gdVjSbVrAfk
vLrng+06PlYW4SvgBykMOmancPIxYjMrLRpfMtDPam4Gc/LssruN7swDkotfsF/U5+qNROpEsiXY
6LBSfK/g5t8wjh9LQevNI+GESaCOdcgkp+DEq3A/jd+oI8RWxVWRpbZnnGvSBCLBeKjkNQsOtCBa
gKIbj5n4W9hapJc8DGbLEHc1D0h/JyVoZ453wKcc89k2R8RMrQ6jb9/IM0V2e2/ZYf/6UYLukZw4
TSwR0fqwu6tUJgG4Hgl8rYp7sWh0ZH9MrDZMqF1iimbsJ+mHMMB3pXZXpCmPaVsFQJHQnkqrp7sM
+zS7X3vee4Cj5IvB9dona6lcqAaqJBqmZrnXCrq6L5gSCOsVBUytUlMYJbsY2Jjr978IGDSsx5X8
Kl5JaQEJwCXfTgiq+a2j7+lXYcWaGHtr2LDxgn6R13KAlezTOmrjcqRapmXdoOiOMIib2s1ThzBs
XLxEAJy2TuKWG0jk4T5srGlzsfWI1hYsk0l3580TiBJCoxKsafyg5PmQBSfU8PExy2zGbWt2LqzR
g+UCjG5UoRZ0sokovOzfHtLMyvP8k5HRiiexIYmkZPPibSX5SIrWKRQMgd7wIcFsa+WAwUWDTC6m
DwpOuf5DiBgtkSEAfOFwvqFWLK53zvI/gbC2LwXP3iIuLQRdvRSScTdNWvkg9klD5YDlOX7rQ2Nl
EbKWpiqU/bG5r9QTSeXcP2q8f07oTadHWWsxDIkpj4CwIylNtZAm9zQ9YK7dMroNlstmMjidrh2e
Sjtl3XMXqX01V3WTEknnNjZ5syGAlBD7vKsx5IHD/6c3AeZRylIs/31UJBjaBEk9G/eI8Ox3U68E
2vc0EO6kC1/N0W/cJdYMt9JwdScduuuKzr99XeaXqteLIRLcbRJOPn9YobhpTDYL2xX1orH9Dzo2
cayXq3aufuHaE3kE8LIoMsxLCxTjZQAuKeXHJQer08AnQ/26ugOHK/rMy+LMEX4KsZTrH6khfoN9
bJ9HBiIT8P6ugzHyjGmmBzi6yDt5bszREgFr8lBPNme0EChzypxddf2lQkxtVq8Hl8K8A7pw5OCY
Z0UFm4u9C2HOCyOLt0qe9GupwDJ8dm54d7pk68sJDB/nDpd2Z+B28HuQ3ehHBawM98IE1qcWSj2v
ARzNn+Jj950S1umsJLLf16+VxNQnIzWwx9xdpZ6P67eOavqHMiIvfdNHIz8y6h23Xg81DwyJPSt1
DkqngoXJdDl5EBb6Y2SSdWNdSgUNI0J7drrTJv4KRONAJ1/JFLJxc7C53wx1yXrsKZ6EYa1gbKdV
7IP8ul+T7ilevY+2NUEqd7Xqc1ZEjN/pIRWj8qbfMdzER1aLjh2xk+CH0VDW84cYt1JLrBH+Jawd
TOfIFH5tRE2RZEv1sTxgh8SE6KOetxw99N9h+g1OD+BX3yUWf+pFfrfPQKjacYmQbcARFcSAca3m
akDu7ce60S1rMpB+P46U1hSvAUPDrlbxZwUVlRm4Y/hmhygz7z1p3SLSN7qUH01rthm8Qr1gg5Yi
KQ50CwuWEus466GnL2+B2iyTBEsWdtgJzUOK8l+EHqQxO0UMt2Pxp/pnPXov7JGl/PByCR4ryvr/
4UnQ0b2/iJ85itQgEdD5iB8IFl4UsWKgXWYthXA/NfB1MJHoF7+DIkuq7+GF4kr2Ifulsk4ozhGm
KTc+UGQugYvnMnZsw/jQDxnSqr3yC9bXUNqaMLOIqawcpvmEzt3OPyFe6F3GBR8iwUKHMY/ioBge
WzjNYdK/4+n/hTSU3XmxmoUVAOY24sCkNxQTHe/cyMja1N9YogJygcmd7dd6ZthFoAecjGeqaj52
dWkCz3oU7fVoJo2Ixk9SQQbFi1fVP9sJtLlpc7zzvUQx/fqxrCdi8MZwBLx7R8l4ODNv4Vql9doQ
qhoAw2VLtkwWZsJcsegXRhxjSxkB945povQ63+3k9Nd/xqIbYR9m5jcwDkdRlWJ3PoIYnbcu0y7r
HJkYyiScsKkMed6yoOKzEx5jZposPxbmWE087yuxCWiFu30eShAM7Sa2nl1fXooY2AWsFLc0sJZU
J5vACYafWf1ULKb/at6+ri6nqor/GFYFH5BYx4oS1ArUWizftuo2VfEYeSh8nG7ddUqwmfK1yMZO
QB8qqAKXtP58yAAPRVBrLHXaGlM+4jpptjO2Cg/V1JRbP3W6z06lyWjNBOzDU14rFppblEKqwP4+
+kmNKm54zpuWZxCnYAv/u7TF8AO3VTRTCkbBjrl2f19VysL3zT2O7TxLlxUuRaVd2RQsXm1pb+Lv
hFEC04ZNHmSHEBVUeKRTFgTo0k7fvY+DGRmqECZV8WYJsDv5FWZJ5aEk1LI68rHQ4OsChtdykJI+
NdmCxIhFf/WAUptAi/LZyJmg9Zx2BKIosKUTtoJ67OVKWqdxRBtwvRBFXDy6O+BnZbiNNphn9QuZ
c1dAYBjhYaCMuTDhG/3T1lhOyvDUAeuDHaWsWHQqebjMKoT2r1Vd/jcQmJY4aeVtXGQxzRv6Ug/9
MGbJL4fUSxHQughnyMwufbXJGCOvSBZb21XvB5tyh3988KJdY8HOfHcnkhzoMEUhPkGmfzZi7osB
XttvYJsZgyiSJzJujPYDL+1L1WE/bxW3AfWtWIJBowJG9SnHqpyqRMFzzYQDMeFkpEBmiRIGlfea
4yoAzXdTcFg5nbbXwh44cdS/de/L2wjhm3ZhkqVzuTMHWSFFHQZbNdil8jEvGlLidDrdv41MPV23
Q5nyRrZJncU3f3bRyoUksidawPvFhobD67b8+NaNyNi8Zy9d8O8PROg8heSiLeqSRAJdTpwn9DEO
74Gr/Twomi1oWrlA1lQKiJqiJUf+NtLkjeJCgKoL5d2cXhyBTgp3QTQrG3qy+2TfdW2LQQVwOAmZ
T/peyXPHneokki98HqCmyK1nvCqxZsh16nwVOcMeEjo8/1pt3QDb26juTJLRQ3x/L4YbI2eZv6Ah
utseoTJJSS+9TWUcqT30hn30arIk0o4MGldvDVn39k6j+TaSta/+aDkX0nc9GxDuG6hgGyvvIDvt
PW1ZSPo38r7mVwpbMgl6C41Y/o63PIWssv7UaGY9YGEx8jfxC+tXws+Q0bLPTGpZO7prt3nx/O7T
mMO8fszopFsrNkxq0XLFW9PMwWY//LgJjJHRIzM8GcfVFnHnv3tf45UYwlW2KpRUl+dMnpWIYloi
e90+zFJODVUJRi4A/7/+JYbiAmpWIPmislyATRJ9OEiVdjLB7O8a/fN7FPUKNhjfNpBJ8GeoP7J3
dA1k67XT4rXMOs+hKJ1sGtQWXvePpBVTx2ND31cQkIqo+PG7NFmK3M/8psQFUbwzo/hG8R3QhjYI
2k2Y9pyvTN2527Ibi7P2A/VYX600NyGL1HFMaEZIEhpb8hMuocgEusYet0oQ7EamxyrcXbWoWejA
6MlCcnBpQumde4HrvLXQPAibYhvOoXc3r27Fc6Lw6T/hIwYlSj9aLP9sL8TMEnOCKKH9JcGPLWAs
Op8Tf9HuEloxuNImLVYu6JlEEV9ba0pE1+DWpY4tk75xMaNSS3GwSzLl3IgYqzGPfYq1bf4c9Nwl
SW7aNOjTaPrVlRIucLavkszCPrw+auInT2drGWarm9CBMW58cobbne5ToUYywYF101gtgmr+6L3W
aKQZe/uJy8ncQzt19+lw8g/qdBOcEnFzwsVkDADzVcv6NVmT5lwz9026rQNb0dH1sA4aqgsl8BIU
leojmXyNNpmZW+eoeDXRqh2ytaDRzUIJ5pw/E5v8wqZ7ZJ9SPkF/rtzQqUg9fkQW+JmMOAaokk20
G84g+gnJ0GZvdKxIXtMGrs/YTkRwFL47r626ZYr4X6yACW7qrB6zam5jI0Y0I56uZxoq7KF5wtJY
1zRHclqrJvwLoj7y4hVwd467odm6EP/7X7+sh+3WDMCP8xeucDcH7fXTcZ9Za2ki6feiUIlMdIxA
/ZyYHFQmQHl4xutoswddWmp542DuUHrd6zKsBy6OvePHCSCZYafiIfhB+c+KaCnB5lSs0PXtdajt
WdDcg8bkkl0V5JT/UtgV4k3vJKF8+DE7attHf6gb8BgMY26TJJ/aWGddptdlBuHyDYMvwe+BWeIc
pQ86ohIxnrwYKUJRzkmCQ9vWUCnM+kCXicG9T7I7nS6a11aDaXM7Gq79QzQgZyt+Fx0jWOXCtRAU
N/ijeEBfcd5i6W/RHRRrZaDvKMpvP8VCieWXTHyrL8pMRZ3+Z+9kQGljjdDdYFgPSkJMc9XrHLJF
sWWDFlyznBeuAHb0XQCXg6UWuJiJiA7SwVDwWKVB2QrOTy4nC46d0X+u9I3o2CdNykIyo63L634R
rBp8jKAXXjRKgBdPd7fDvFkRTAmmJOa6sPGNxUP/LM/b86s8fqOv+Um5i8Y5KEwbTGKliXeQvOwL
5nUsw6axyvV3WcXP2PhetRlAzD/muE5MqLh46yPXR1AjE8Utm8wSqHBoq/939J7XlWrzliYLO0ou
s7YK39QoOcQ/YyNf9KZJpazLPaMTGvDHoTVYZsNOZ3/cagCmLfklBhFE/oGPvqsI8MBUDIP/nfXb
r/rfE9yVNN9UZ2dxPOqvV3sFh1wsKhOajcQG2y77JzPzcyHv4L7F6He7oabV36ZwtlXTRWOQmor/
NNwpZk+rkGpyZIPzOFaasm5XvSZ8J86OAHo+pTVffU4nH4gG3GTcT1KWX4Vwu4m1ifCGuM0bqnMv
D9raB5+mC1R9gITl3TCEqjKzw7yjcxPI9brJSWMcy+dLdA63pqHm2K4rL2n4fMEIbttm1M6+rVxN
M/rdSRMT38kPnAC3ylUNyUCMHC7yslVYh9jQVhdPjvEzUOddYkqXvyCOWxJZX9VJAXo8AV67PPQV
TaiO5JMGy9EOw6lgvZ1OcyAJAFneyL2s7cI8icj4feBbu0kecfUPBIYb8jMFi5KSD2maS0hsCZ/N
lKg9m7PJme3Zx5C1vajOT61XQb1fTavfRntBL2LYv346ptveYqMPGZemnLu2jFMEGMU6LLGU1txj
7d53jecE2hiv9bU6dNhC03IY9g2R5zZVx3h1yWCIPHx4jlq7P2gyHPGrQrJOPV8mGcNwSCr/Kurf
bpts4wx1qdDRq/5MfljplGWJi2+WpnsIwvvQaZ7etp2ZRox3NxMRpjvfPQ222MTpqqOlrsR8B8D0
Z3jkEhKq6sIQ5m9nSFz5Q8GOFh0SZlErZH+BUevxujqHpR2TbJAQCyyICkatZIsNtQTQ8QDtJykX
5ATgR4Y/9r4s+seXTpC0iICI8vIiHhMqFHrg1ROnxfI0AZh9LJIO+f3HHtvDQ1CWFP7Q1NHBcAEw
1pBQ9Y+0SMAtkMfwTWkmEnwSQ+68SUXNj1lkVlr7hylCzoR09osdniEBKvnvazK+149LGYZSKy2u
ZDDKYrczhqE1RL9M7qbh9pNFSEYNYr4O2oQuqeCWNv3lfcy88LYJr9gqlownS7nbCz1z+lCuO/gw
yp9ZyXEjErkjoeDwL2ptYGFk5UrpLhjWuP64LHfLpWel+lpunWvl1DVcgLgVucEY0utuqzYzHWz7
O5z1GVSxPaDoNBNLOGuOBzlj9Nvuib2NVT6FoMDogkFjwuLF5SqB4Gnc100Jy8GyUMEXym6ArqI8
tIN3f/0hkfvHtMzCCoWTrWYOy0PsDj2tiohlv5V9kmoz+cZ7lVRkVTD45BstgR3GAct9MW4UMKRk
z5gxenkqpVGsMdoSARPyDG2h4W8DAWm151+dvOoZLsuwDmLK+ZW09EuC/RkKv5jPubqJxsRtTeAI
mnsO5NTw8tl07JLIBhIf0WMq0JLkFIkmPmxfkD422tpf4RjJ3MLD6dBFgCFndcqcnVc8rg5Ythan
2dNxKbukbykRMkj7Q2Xt+yBf0wF5ItnxKO8n7esIXOFmc5fjbnps91qQgmszxmEB7LuZ49v+KCjU
+RSIex8yRFPLk66quHNdtjTNgLASxGT6P8TiXxs7YbxjRhoWci53K558A4ffE8etMi6cXZxBZ+Ay
u1SxE3N7QO7CX7L8nm0WhlLtyDiyz8Dw62tMn2oCZzCiu241NSKuFk8mUYou0wGqhjuxYVeHD+bK
z3vCsb7DGlnL4nIXNT6Ie/E98w+fuiCo4xpIdpfF5lURiqENgMoPow1xESWaVrjyHjI8iYq61x7v
dt2j3Jo7rmb3Zdfa5qEelwC+yUb0AYlVQVl8cPKDdjKtBDLSKLqKAtyqs1K0eIym3Zi97acZd1u7
oETxSpN3z/k9bysy7pW1KbeAiSfIJTx+Jffo2Q+dnPxBOeD5VZ6iO2OM8hlVt5tpKxD7y5Ra/knZ
r7MIdtrt7mNttArtflEdclGyKTiDU0SmeiZvGfBmWrZEELYlEZQZRX4iL+tYAgURXNbcSekghlte
g4fVD0AFhtRixSYVsfv8IuY39fmXrlXupUVy4MxsCknI6CG9UaMfJQM9bFFUWOhp8PPeH9J5Sifj
FWR6JT68we2uZK4to5rzaUupPXybC+wFWnVHGNVI4pITkk34PjsosqAAfbvu+MWknN/rg4BktrcI
OmaFf2STpRfMkBNSG1rmrkr05MO44Jk09Ta1zn4rDIJ8Ta0WCd2sdIvMThYe5VOjL0kjBQwBSj7h
XoNJhxRfOPiwSRRodc5A9KYbLde+VhN2kq877oe5v9KRTozxHN/2V4e7ys6HudKPtmBl+6ARpA/8
5gqTPYj8lD/GSl5ElnOlRiyjdW1JuBFo8fjQhLHNpatkPHcGc2q6Fzykey7W6CNP7xQAoH9MdgNU
PGPedIiCme2C1DlqFeIvFDVaW4rYM9hbQQXjDTsvyc7+2Ym1P+dRtcddOHd5z5+/O9Z0bRaAfVZU
x+GMOTBazNmi4Oy6lnDQpa7nK5Ij+jcx7lbOEt+LoTHqBJpGQVNlJG0OyoHKSZOwM8XwE0eLcxke
JH+/rkx3DgjSX5GEoH056fidcZjRTVgomzs3tVW68uc7UU1a1HhYflUNbBwh4RsdoO50/hk+3BB5
vaidm5yTG1XfU4eC8hgzc96g/iJO0K1jx+1Qa9bC81BfDY5nw/6Pt/GXhvcP/YHP8NC+ngIuNRrb
waAtXzbUFWzyZpfnsGKer2xDXXRhcglrNSs+EBwYh556dZgC6woHgu7wxBOHSxICQXo5cj2Y3vzi
ibzg8czFR66/mkydCm2TcOjco21Cptswu2l5zm3xvkoLU7porvLUolnWtT6NvEXO4p1nG+jH9T+H
RrZUuGLFxLpp5eiG65esE8vrjUCS08DymDZFYLjJjqX1L1svV+l7pmb0Wx76sMJhDdIIRgvsYfwH
eQ8svx91iy2172N4lMS34HjW8xGQ7AnRbxoPDXxWQNdQx8HDHKWW13eWLBkrlqI1rZYBBPeHBnXQ
Gf7DBHYgG8kXYDTV3nCVlfD8QvQ4FlCygsXkfDBM6IhGMU1FXTMcB8yE/7iAWkEOEMVFdl2RhEdH
TBPnzbvRAPnzNpaAEJaPQHCIxFncjjqa2Q0UUc1y9r8JgEfv+iTz6FLZxSSyZUPZSK+euvdlGbDv
5KGRCS+vau+H7Bq7ShEYBp2lFNezDZyDEunMt1HG1mM7s0hNa3dECLTYsmU6FUYJ9eXVGbPr0KUZ
UDV+hTJlnXsci3H0P/md5vgzzNcjwXkfza6RIYXRG21uY4pQ0A1KBzMYlNVmpzSQuMmUkl6WV35y
AiDO9e4zgwc/R9oQ9PeoKb68+jiyWfKLjaIUNRduPRoEZwvwms6WS4xzqJHfM5vtiYKI/bgnId9C
TYxZzJJPuBb0PYYx242zasPDmu5hYwnU0UF91JkaWnr8DMM99LXbFp09LY3oTZ8BLYMzGB6Vzv7v
rDm980/eQ2rPFmDIuw19LI3IVi8V5m6lmy+v//GtDMinHv4mfBre1aFMByku29v4Vyu09IU+NUMy
bKaS9/EuEMINM+s893zSg4Qfg6W3ZVY89QCjNoQPhQjfsNe/8aAn0/IeZ6jMlwqIN81pneAnJ7SV
J8QsTwqlWflKBGrLXMnm0fi/wUw/tB0c9S8EJfjjIevjFuj2bBTk26wDS81DF24zy4Hc9HWJBdcl
BB5Wf51si1hGPlJs3KKwbswnMfrlZijyaeqttzUVIFc5Da/YgA8XmlN+w5hPJ7S+xV/f2KdxlMKZ
3ieKs1807s54j+ux2ARUimyjNJ9F8uAnGsLreZuZwbIN6gv7Rh8xEsgBI0uniAqlwagD9bnBNI0Y
7AAYhQSbOGJ2JP1jVKQ0HJEadCsYO6Vv9muClb+mUTlkDYgtiMQ7r5WAG+43yl0l9F7veWck9aDc
MDdGW6askXBPSpWWruM7ubVhlqkkGGkB6V0ipjtF4CdmPj04IkryvphBjVFpjHC2jADpQFCFZ9a4
CUrR5fXiYOzcSgKh1Bq1dnvKEN+xHgQdpn35C2mw2XNdri1MiFFDIpt/yNENG6Eg14hjCYoLlpH6
mI3Vnohz3bZWAKfEQHwhvdrqf7Iv92Gh9JYDrhWSHpeh65sScQr5qItI6uM6bQyA6+LpOmWsaR+i
ZtCduSPTKRpPiV46s2D/sxXFxOO7OMxSbDEouYkvpN7O7UAcjINfeP5xQfi67zRR6YD7C26jD2UM
YTN1BXH0Linj/FAPpuG5u3ohsWvr3CTDmpF0VrP1ZmDVc2w9dH8wFhg3eL6FyRkP2c790hJVo2wT
4Ri0mkf3coaXIfgTbIlKRmUwklar3HkXjfDrnPqsZ08/iZc8s4ScYRPM6i3UX+DdvTqWpZoQLH3X
K0e/b4isoZ6UyJLLSFGk/hvfyic0aHRi3gbyq6Xdoem1qek4ybCzYZsPiBwBZpZOYtrw/T74Bmht
bfDoRNz0q2jIgVFG+KdUZuE5SI9sQ6oncqFYdbjxmkClps9V8TAnOKKEefWGi+Ves0COjtIRuuSl
JYVtMcU5l4Bb2KQ5Vg5jIwoiReSdQBY7j/NRT9MrdLgEMJmjEN0JUDMYPHOMW/BHgCcD4ncpMpYY
+VWtYnj3QvzlOlAUer7kZioyg/4RaS80sBdZhyNTsb2PhUtK5upplTqWiqRtmR5nGsOkjp7gdHXN
y67hgOaFvzaQFgSfk/U1x007WimNErDtkGG5dw3bg7d37Mb79RJVDHGhIBVTAI1eRLBRDBU8dGAl
BslarT9ONfWQRUvTtCih59riOjUlhwUddYw+Z1/wDt/HMVZ+6tfyF4anN/3XuEcV7AjOe81NY4eR
SwCYRUTWgXEz1AG5Zh9QxMq5MdKG7V0Z9z2L1ixLPEgk5x5KDfgQ6XXcbIn40QlR2N/RV6M831Pz
HHTret76jwl4B8VkAYV9bUxI+CnexVO1//2eRQ+nw8ie1BiNsxooSNwPS/g12gsp25XR0xSD2jYd
jjNy+TQU2Vp+jB4nLVWF2pDRjqfG2Xy84xkF09Pg8687L4MvqRAIRa7/8UmTqKjFOowBVaGXIxnD
XQGh2gpcQzegLcTDLFXfu152VjxS8sv1PjQEKho0feqcwC0FAadRqHlUoBdr+sA5JMZGzcq6yBmk
qHFR7o0GS/gxAjkpg1u5652NDniOvRED4cIKMm/kg/C3e7nZf/tQvP82nIii8fsdUAeRAjYNYbeU
mu4JOBMjtwC67RuOMwX3B7oR7XbLJTOllPfE1tBXZrNk1MjRyb9aDg5zKcC1Zcu91dyAzWAnKBIJ
5z6w+Z642awDWo0aNVTaBcKLwOB7KnQ2kQt/jTpOPUjsxEsnA8JYnLx47ispc+uRkBUmiocN7Ygg
PShpiMa15xZ85F3G9JLTCA973NuffYLm52FSIQ3Vc4UweYOsrofbkrGn76QVXz2/tEYhTGzbXb16
9ztDlLZ64rztNng4IuNj2Ebnee0AaR7HQM0kzSSccXmRfjaRdHeYfy6I8TXGPNWjUhJ4A+hS1aXw
9gQLFeq4EjjvO28BlCplYotF1b2LCZi/mVSqDstnUYp3qKXXbc1iFdm2UPibPRe9E47ea91Uzdyv
Y5+/H6DXPm0cxw4S2IZAcFEQQYpJaVTGN5Tb+BeAlg859j19seD3FRdxOuixMSPzQb+lNRGIS3jF
2J0V8ROLdo4RssrB1YwVKkKhyqurmyFMepZrf0NjO4MKBaOiZMMVvjlAKqHvo1bzNb0s58Yfb8c/
gAY1c6jbG+I3s9w/BAbnzwAVKa3COS1HrHg0cWDgbfPil4+SwpSwWXwqRG5t57Uh5V0uHgihXL3u
lRNR88p+OiAphApUYp2RzzSM7Q3mkBul0uxlbMZcxjq6QSMfW4szwwK6ojuZ1YPRmKwIy/KVv+F/
QA9RoJS9AaYeOA4hqnNhx0lcYMOf4+PLWxIwAVOPJP0lkMUxIB5zobbIF3d7BYvlteNqZlzp32e9
pJdmJanv9zdHVmRmeQhGfvcT+18ewlHrZUyGyjeUDyUNH+pZkz2yxDQPEuCoKaGxDic7bbaw4Egi
gWv4rijxs8WoKQBhnIY6eRFgs8l/r9J2DAWK117WiTyBmSVj9jVAQzTi9n9irpV8pE7oA3YUL+Cf
GDmbq+y68RgnLWH+qg2xggrYtvoUNYA/7z3q2Uwd0F9dpfAbsQOdIBOH5d4JFn9fWda+X/N37/1o
vp1qf+G0vxEhwaJshPyt/qGHvbdMvqjCkmvPkHmPGtAjGnSRbekp1oKmhZYUVdWivnBfQpH1EeWB
799vC3NbNGdKXuk3DXDqVT6eqkSkwEfqXUgqAGWzmzSj7qMy+pWruIgjxnmo0a3yq8UJ7kQwx+Gy
9WvW/0NBJxkwl8x0zd2jmtaabXb+XkShoIqFIBucGjdZJmjXbnLAYI27c5FgZRHw768t28G0sNXN
sPQWk4iiuydVpktpiJV9vYzZfdEBMP0jTeRRNMjjlqnSfPXqkdbr6XRGDtxrnI4xAlNrcWDSaUTb
9Ow6s8nmOIfKgZ43335j+oWCeHV3teEsOzSmT5uojkNSWgnocDZOLV3iq1JVFhmYS5rvlxU3DfjR
YCvirtwnfGbIaWG6a93DJI8nV+Y9muRZDOabJd1lvvIkCHuw/1OxJoHX9ftSzvWzx9rwbbnRNfGv
SL/PUvVHcYg7O6yx/0iOc5mGh/dv7wUiwqMLlqHIroPohus3XYaBcOPnkiYXsnztv3YcxXk7NXFD
hdVFGHTUcL6ZtQiLyN4vN+ntJbcWPkX90sozZvr9LrI9hNl+u6eHQ/dnulC+jkDDDIqcqCmrxNQv
Ia1RNMr++DzdM9yqn1uSKN+uht509gdh2NG/6TZ8gvJJ4s8e+LPCUFQ+kTmIBQCfzF+sI3rzO9I5
8SGP9LstBEGoj9jmeZ1AjbPfscfiuAWTOp1UPNXZtlvl+hiMBx7QAxg/BvmS9lNZDx8AXcWCJyh5
Jw7lrTLhS1bu8GtSOMgTdgfXBGE/ywsZnZfaKs+2YPxl0xqYxRvxv4snhs2Jub1LRdAbUTmImzXp
SHjYBpd4XZE7YmGQEB03t+7zkHz61Hl4zi+rp/JPQakjM9Yiv36E2wzwKERFooNW6CgspYCUI7bI
VGYUm5KG8ol+zKmPByoiL5at1OjJs3bz1WJUiChWwX9Um4Dj/SdVtB2sSQ+QoiKExQvN8xDlX57o
BUW+09M5WKS9UaWsM0VTOB58mfl8sEOAla0QpsfYbZ6s45aiAVKuOuiI6Gg3TWPNcpD+IdfDYk8n
wBQxl9g3zT66xr17pJwlOAyCf+LQ6V2Dt/vGthHlkdyspVaxVNu33U3O4L+yoHrIeJBwUlWyPlM1
SyMGLbaBLQCjPwOhDDBH3k3gIqRH/GyjBFQ9eOYh1olYNcqw12FG+6fDgFHWkMWt/sb/dEMGfCVF
kgVtWU9BvrMR39tZ3a7eYGHA2Pq3aky+dmz5i15DKUXZtxmv26NYcmPtLuE7lvl1wySl4QorkeDG
yR+wwMp1SWe9O1qVudhvyl3Qmsf9oJvomBG6+z+6Bpq/qqdcG5tgHrZs/LSAjRslDEXuHwkDDvsV
VoFhzLNRjoRZxlg0S+/tPRi7whALe7GSiwfQi8xOZiUry9EahmrERMO8UNjFcezdR5Q7lyOtCwT7
qAB67+Ndx6P9kcuGXlyJfKv23FDn/I2n3NiivncT4ROhqO/8Qt7MlPM21+qf9yHONYa2KkPEPLqc
OpSlS10LIVNkec/5GylJOBeHWkO7ZA50hA8oV2/QyT9+kBnY+n3wOKvvzpJZ6yOWSSk1Zee6kt0r
tPoKUuqxvTJC+0HVeBAMEPZqefOPiq0ckbuc08Tv/BI9Y46q+ZfRr3A/J/hkBY7Lx8j/V8tCR/oT
4d+Mnoj1tEPy8YAH4I2cTh6wdaUFRXmgGPpmKc/HKjeCV8Pt3ah2QOOnalq/Yu6r5LyZY5Ocl7TQ
Hjtkjj4G+YycOnozECXvgHO+u1fk4ikcDyVmHT15Cp/FBIlhtP1TsMONMoWlxA8Amc9X9XWZWgrY
DTHanW3o4mEomVtETrTpyGarErjiw4a/yFkrZW2qe7gVY2ADrEFSb0ev39qQt+0tWO1IEdDoIpCm
RHBLdBN2W9Gh/dcNr+Rh0FE3fjUl6rJ8NmalBoGXfvpKx9LYnorhfA5uKovrk/TbpmCIPlemHDkC
rZxUVnAPkTPEYVmfypIMimheYOxdWntEstYUndw03VPlC6W0dHiE17f+GdAfe+dJCVzGd/wD9BVT
oHnkH+G96f6c4leaMDfhhKOUOA1C2nqHduqnhCh7HWUBdo2/dD7FrlHpRuxmNsJS9pXOyym5u8cg
8IUsFUadwBpXBneZOcXcv7Vf6w9uiVNDRAStuawTaNu2GsWa7lN+CG7C6WCPvs/49uLM4a1QthqG
MxUS3A6FxaKf6Qj1FrQ/+j60n2EIZ146WTp6XWmSFPUczRATMO4kALlQn+dRLmP6QAzGrRWdIvVT
VxHI+yQaKyYduYMedMyVbRghYPZaqYZyYT0Zwxooj36e9VAcb4pWNP9skHOaqEj9lK3AI9RYuDVf
GnwqCqTo73VT0RMAxeD1dvGhyJejNGDlHqVuONd18muO0lWimyJoo7b6OXpsXUl+HlOJcoqEpqXJ
w3esPUtaz6Ig1KQLb2DypluAkwxGJB6+dw/sAsk0FkwJNLi0fFwzMXNM49NQy6nEsYFt2ZbQ/K4o
xY4D2t7LlTO4kreOdjCMxzubVne1y11cVPxRAtLaGjr2LaKMVzhp45WCltAl7ahBHQfkVtV9+VVc
rPYqIeApa8Ppv/KFVx2JD0FELLGp5LRyUN45NjfIQHotyYehoDFTjqG1cZdGGOgeFvKhi7GdqfEW
bHKLLKL3czc7tMpEWIAsJWh34GOr7WleFpw1QbCta1NZDerZ9o/1KECW+83tPopUErtZ8sAh/9oo
ZBX+9VcF6qldlMGN1TtRl5aLV6BwVQAE1ZD2Mtq2RZr+Xno9rHq9mL8HQtZR+dGRxgT1GzhcvrUH
e39H9ac9wvp/O7Kyw0vGTscWp1bfyP5YL+uHGwfPwcdwsfZYFF9ex5sHou5x0bTuBauWiE44CK8F
HrlcKiKQLh+YVkaM0e1iwRRIdUX2Z/ftwc03dp0bAB2d3wq6EYk51Ixl8K34vCXyNbXFfEbLEeiM
mkxVZ8hKqHT5nJCvAR1Ibm4uSIN5ihEsc1hpOsBK1o3SaI4mxEcprssR2Ct1IG9L4Up5Nx48cdsW
AyK5fX19OUYVfeocHj/+bOOcODu3h+ZIl+Om6PSOxhOrOCdfPVL/RYIQ4bZgL061Pcg27GCkrwM3
uP/xnb7O+Zdy0QtBP8yPHrr9E+/ixxyXafy8+W5OrobJKO09MIjLd+tJ2AlEm0MFTCOtdXmVEG8l
6ENQf6GBSjFbtuGYx0Vk0Eqfhwnvo6tpqOGE8qSt6+CPzAsik+BZ+x3Kf0YCxexjZdrKuCYVA2L2
2lN/a468E8pI+btj+UuGhj6YUHKORtqGDzzPOxd/dIfNkwSuNVkjQz3d2kIanhCKVVTKA09bQNzH
CT0DKp2ex5Dg+RY9cXEJoOqyp7/YDcsO/uWKe9oS4b1E7tMR3qnJKruSRQilriKBoIsp7ABAyQKY
rUkGaHadFObpefEkUi78FjWFCMfa0WzFArviFKU16fqHFPSLw7vhYSwjnzxxQDS3wsJzyYL2BFRQ
kAbciIloQbW7fp5QhABbncA5fpiSGYGYiTD31s6YsQ3c4XeRwVVaP5lfAFnBwWhpUuWnkZkiwWaq
q3yWKHBPhqXxH7ZKqniAG0/R/6+ElHLsBrxs1ldNl8klbjlv6vICf8UPxXip3kwtpGv6FIDbNg0/
SSZxpmCQGrBVY/B89OniKpZLDIKfP+GYf3E1pA0IOyVg4w2L9Vlt6/j3qOUKZ7IFEYVJW1anUjKV
Pqvxkei8TPi0JpveiIxpMFqLgWWNEpqOua4mqLOvUZ6eHsxTnNJpXDXZUXztr6YlwJCwIe8rHfd0
vzkO+oWacnG3kpk305n2f3S0EpD4jOtWyuHK2eyBlU3kEvXveqg+0pDOXQhhAIS5G1WuNry0CXxl
p5Ak01lUL2+z+hLXwkX/0FCCxvdJGRt+Fphudr210ry6rf96lA2hFts+jZxe+Sr+rzHEasbq5Zn4
nqPgcex/DFpoYGd9cfFaWm4WWF6PWyLoXK8v9UII7+HKgo6r6PM8gBkOBcgpYW2YPkn8qfR9+GvD
Gebe+C+SgYe9ykyc9cEttfu7RKejK6MaOD2y1Bpy3mBIqZQqT79jIrbm5o4ScWdEO1g+pl+uTZrV
qWFvY8gFkCUYs1AeDRiP24m5F3lHYcAKLnvZ8tFOK/GemHmPe3gL13wMlQbZNFKM6bJ0lTEtDICF
MUDGLMXSTYgxCjNYLqCVXwowEHcqaP2Hb5UIcOKf3p2neJ9U8iCW8tIMTxHPbdbVvhUsfSPeogMU
mjsl3mYKZh6jEDecEZm7676zOAweFWP6kD5BVsD1uJ1WRC1idguxwWq8eBX31kE5SVWINLE0CwpJ
5EOS3BB2rscQPgJwU5u3TFV8a84H5YZ4vs9LhDv3X8lw0/Ghe55sEd2saXBrplH4niVWGTy21/lV
rzFeqGxj8/aZJjeHIS4HG/onFNlcb1wSi0hAn+Yj7H/YsvpMEpiNPP/w4XBMXU8YUDPo2u/7WWNW
c49sXrSR9sWSKa6O1Jxq9AYWM7jveY30w/iSYN0+7pEnVqwFfJMdAhpFf+3bO+oBf0qRCyZvkEZl
HP8+zvEuCvGbP+c3JBS0Jl1y0P/RRrCHoOCYy1/4x8doDHMIlk3Gj/XWPKKk7CgnwOpTw+XwTqAP
EF+y3RRX7ECj0bG6K49QieW7gbRg/RZBdboaxrEoMfzdsBcHzy9wA/k1ly/2Mh90Gyyw3jWAQdHc
j1wCp997cWxsBc2uenb5VRsg3uI1PHbY4q8iMLqNUtP1xU8556TwGVZjG/sCbcaHx3Q8v2HydAxX
LGmihf+NxW2k1NgkLd92lxl9PVV8v4hTfNJ5A/l4gKaKeTVTG5KREsHi2Z/rtC9doDcLyJlPnxU7
CWwlH6t1N3/snlm1/S97wqz06hgJa0tHXTkduK5s2oY2SQxBuc4kgYvNWOyGacZosoP2Atvd6OYl
RrF80S6/Jd9M/H8jMgPAsLLNGCa9co/NPLSoJ/mblieuw4qr17ZLhqBueJN97odSD/9M3T/e8hLV
pQDtkIZZnnVK32/M2ZCuwj0YMt9B9FZqzP8byDKjWvRI/JuQMNctcyvKpg77wPD44DWHcJ5N2bY1
m1KtK3+xoriV5rCC4D3vwypdmOjLIvpltUjzeDBoqWaQj/53mjzaTFroZYbOT/JhV8Lj037kLdBp
6HOG18nQU5CEcLlM3F35nSFwoHlqY0JtwN+XqDae3kl7QgDgfc17J7uE1YHE1b3qQe52lqOt1xPm
2Xsyg5oEJkFUBAbnDcFRw67KCcRZgiqygh/DOIxpc/UWULxVkCOBe6NxQilWj0ha0yhxLxZzGDt7
KpZ347+7uk8WMCcvbI2wn3ZnvqGiO1GF7x3IiDVHygQLT6VAAEYzo/n2cklBU9OwHbfoV+Bf1x7T
TDW5fu0ma0wdDXNaS4gK1Vb1p0SmG4E0dt34ehFlB6Uo8IOkW/XvJKrJcG24JaP5vNqiUN6QTJKn
qKr40gSOFwwWfIbe4oq9LebsyFWBIZW7r6Pi1S//zXieTReiv3oFm6jFexYd5Xbxkn7cdJ9K/M5U
W5mlah/T+Eq+DeP2yZDuQiXKcGjuF1dGb7g2trKgmnY8c4ACJYR3PR+Qa5qhCeTK2lL2tIatkymu
YK1XH4bRc7AhCfv0WEa2KCrW3ybeJlPi7W8ccA4ZiZ1tiHp0TUa+JQWFYD3sbCiBIkozIQyJb3CT
9H3j5DfogTHfUwTChG8hY7HuQLyPBMSVvS82x+40laX9Sk0YUctzthq8+Xk2MUcZjGJMoA/USjSV
OWG5NFmOiNCAtXittZE7L8M23NHZdbRce1BY6xZYYS0U98o6huWxcjT4c3Ku0nGcMHvxt+fxMmss
uPRFGhJqwKqv7K9UX8twFWWE1FEyv2NcoxLchMQiZauUAOUBZcHk48UIKJdA+DdfEkyR57I0jlaS
wjuGrxZCMXrhP0dx+QS6pnp91uEMiHvZy9Gv0A94QJXN0bHtHQQeLjvvFf37tAAGXZ24Z6FXerZ8
b9cvYmxJoh5xb9gpamVKhLkdoXKnqA6IFZigVM1Xf5HaR6dtvtEw63PnaF0iuF6MtmUCAjiKTk60
K6ZQVbDWmkw0nQ75ODvrC09FW8b0kGQEM86N0gh79AAI42JqJB31jeJmKKiwB+bDGDE2kNzOGP4t
+Wx92eAUm+BSyR8SaJn7i3Su68SwhoiY5Qq7wdmvRXWoq7mT7xstlaJXtMH1LfGAkicAB9FTASVA
0iD1ztco3B+aADTQjAbRd7VoMd+xJ3cWrU6VZsMLsGo55I/ysGp84+4kv69grXb4I37uXoDF5V8t
gI8UqEKJtLKjwj2bVyrHoaujzmCHfVQhRhK+AHS3g02Sr5lXZWolvT68x0Huf1WBXI+cZ9bVMGXt
xylZkPFXMEMHxmfG00uI+PXr/5qXVCk1336NnABnHA+Otm9Cl9UXZvnZHN0j0ocEl0kLnDr18Qvn
4pKgEMp3Zti55rV7cJp0816q3PXjOZVEEaI+NyU46FHFVluF7EfjXMi6dtlYXHrFzpwdlbWppWjG
xa4W6GR/8KFzSX0KW8/LCOfK117L9rZYm8Gjds9ASjfmcNLy4FEfleZoE11Y6zF/7pjrBZlE468b
noAjHCFZ1g5swbEcKbXHn0Y+cmF5J28In8NeTWfVUMzD70P364+KDmsIasmx3RBCpcDKZISbITrL
nUeSUSc5u8tWADXg83X4GoYbhU4WHYgqHD++C2DUeeDMAM4pwBn7muoI6eK0VEbt3v+mhgu3kONh
PnVl2vTAsfupLYYnnXYx7LxikBMbmqGmzoFq0kVnpSvgJZhjVqW8UFex6cTLNKoc02HxP2h8LSZK
UIssonm5zjm6RrAO35OBq0hZkOfz2tIhT1gzeOpO4eBSRMtM8oFyyjY0zifDE44qq1qYeSAem3m1
85nGkyvrijQNXhGMc15/gC5cfMZh49j6wKmvYBr3dvMfHfPSK0v3NboOQJkXcDZAADsRxFUSsGGS
IsNdikRt2g2cVZ7L3hbbeP3dDuRq7pFe/yE+VEllpV7cEA6w61uXYdaqOlkH2aeI9833f5x+9XZz
EILjNv0Me/ZBlDTpyOcWp8drhTRJX13hsANdXB/9U9Mf55WF1idJcJWCXtjZSJQ3TxapePjibSB8
Sf3gxzo1VGgJEFRb5H8NoyONjUWme9rsVcngfgta+RjH1L/KXoqRyxBgy56r72+tJ3SvgHwEds1D
PiqkZuEPN83PGF+RFzyi5WINENUiR53nNFOuhDNe2qxytpcVcYXRr9cNdtbknPJbUk7Wkx4IU3Nk
AC74cW3S/W6gMMWrpkmVlzLi9iU+iwxj+CZH4eKI0WnexOCIZPFMaDXxTHgohXRvdLWY0tGDVZ0E
WhjkKWovRb7l9uKu9QrnGTNF+sEPI/uuL/w+XKaOW1lsgO2M9v10HuNtEk75qqFL8EN9jqv2wDZC
Rof4pvtaRfshF1AuNNiLMGFo5G1bavk8QogxEKl/ja610uULgwoEL5BK/pP98XBK+fMJeTzLJ/fX
aOd1NCaODnm7geheXkHhlcGoqVSr0Gmbx5u0k8ujkL/rEe/41VOf70yNGOJl4L/hd/mCB/EDFvjd
AGSA4qBUuB//2ENYv/sPCJdbVIe3YlKeHXOurg66Jt6YJ6oQzlTzwfbVpyDogBdQme9O4ZBCCj+W
7R1s5OPQVVCRQXYfQkkDFWZOjU2GsII/ylcxZPFFccqCWoJkkFVJMPfRziVUhKyRGq7Fsq7hCoRc
a8tfR93Zf7xVx6n6yB5ZMAYV1QsoleeH6WkCY4BjoXk51zi4OdFQEa6sZkSj4K24uUO3lxs3fIRr
VHeOqWykUq/FJRyVTjH9Gp531NlgdDK6iI/Wb6dwhndrM7YUPzM405C9KPItf7ZuOwWD/0JgDm4d
XTsdlfNCKGjXwbXD0MPhLTvnEbrxFfglQGtlHPKXq/dd52fsA33p02Rto1hF2+8gel2nz5NVoymD
djyCk4Ao4qHjv8pgLfBlh8HqSUoc8Wg159fG9EMAbuMdPEpkPGtZlMlH8k1rVRzBMOp7P4ELZ8gr
L+IIQPAI6A7nUmeBlWhNJONb2zIvm89w77xzjZG6LocFkW3fCnRYRr1QORT7jeyu29WofvRpUdoT
A7KONXtgpr+JMXI2ggQSUsTma1f8ZgiyA6B8jTHTpspZz01joFX42qcDW1PuxWwJElH7lxfJPFP/
9GU2kBOGS3EXJO6/LKxcf8WwiUl21ym4d6d/q5sLQOoD9viFfGkL9xXzvSpYNlAl1/zkH9t0FPaL
FQRNpHN21Q+uQbnSBV80RqmTsamv1vKa6U8W0f1IEH1SksXqIm7tPmIJ5ZvnZtBJrDulwVjie0Cz
ZQ6bqKIjxT9OILEua7UpI7HgDQtrYUyfw2GUCZeSEaqYWh52fThqcFcLgCg9shdpV7Tc/e8v4/pM
HEfH8U1DKrZnDCBL4Sfn+t4OViZnm4eoCxuxduaLfcPYEJ7Nc2r1/NFYjF2n8AsiibVz8y7FrKrb
CjVCioRIrszx/LNIPZGtARMby7zca6+LNP+ZpKQFVyYeYb6ktHxNSkYBZnJrLKj0gbCMVvdCna6t
wNqT6Z9rBA6kvGUtijKA6VnzuJJ5pVUvgCClTYMc60gIChHEH0B9kp+yRampJkh8pCJwLKn8NGcj
H6GRLyscYgBX7Ms8cvxkIPziPk/3MYPPQnj1NkI010Vr0NyrCFbb2CQjs//G4cg76yPUlsHDLrzu
EctztLoDnt1isXNlAMrFOwotzfPddjhwTO9uzHBu3nhkpf228b5sBecl5TILS5I8ykF994lk94RH
FdL46S0/Fp9NifDUgjCJ5fngVpHi8MNz5veRkxBq3rXWZQb+IbrvNL/83nVfXypECb5f+flJi3In
xeVaScJG3k7WZVFwiktBYdF7I0A24Ns7p3Wc2Ad5AcoYyPCWTD5kBjetNp5aUKKZjt2VUlpLyWcb
yOjh6ERbN97C6sd/KaFS//czj5I9PDuwxaR/fKsv2iHj/fJ8Tmme07eHY2wuC5McG+YdZKsrcrKK
Wrx006iEe4XkXj//Q10sVcv227BkeQGDJ6akMaQt9hyh3+WgDlXrE2QXQplE9MPeUtzKnu1m4CVQ
0IHmQdQcDN69R04px9JLqjWDVidjLTsmDkuRw+Hn+y+JzSwMmbZWvzhKcUSeQkVGvU5XMsrPkrCv
n8p0Jyhnl96IAfZ8ol0GJ4HWCwvM0wxXD30zA5R4SSI9v8rcHlI9LX1uZHz3HrknKPl3htpotvpL
oe+bQKicEJREoj8oHtC2/XzNuvO++D668GO1M8Tpb3W8zhW37NUuqAAiMoR3KilUPaep5mLJx96i
nfym/pqFT840PMYy0PlNhzybiyWlqQ1v7gPToj1LH2CMeQ7BecQYyeBZYNPReUpz8z4XSYbeDy4t
E9AhyT4V6JzQMFZRRz8OqiVUaSxRsJSaQWmf6CjT9eRw9ROn4DeOSZQOz2cBcQJ3d74a0q1EVWDh
vDhjdOihd14/M6ZKRnlXCYVZbMVRWrc2hXr1velCg4uSyx67C9LFH7PXL1QhDYniNNTOEbiVAg3g
NCmEkH/q/h3blzHxHkHqiSaDNlcg7zlly6gWbX6DiW2oN5NyLu29+XaMlIQ2VqLvlXIMSwEUPj1q
/1aGv5FxgoHI839ITAoyOhJTiYf5GIbPPLFqkCcU589AJZZrRFt5VZWQCt8+yWq3GYwKCMeLYjc6
d61yPb8oZDqpw2h+7/+SID1fUmHNEhYFi4JLd1TlsMvzhOqYO5RGSZwRxEiSbbL8tuoc8lUVN7l1
5uQDxS2+tT0dftmZy7d2vxLVH3N8yyWA2Jz2S4FGKU8KUNLc0fR0dqznVzJf3khhxYzpjDmEtwRc
zvgG2/bpSIDAj8hYkee3S6TKkxMdNBrZikK4kJpdoyB2Mq0Um6diJfkcf2Eb1rJ1QAW9qwKeO5xY
fSw1q2kL02labKFhegGs3qcH0YNgV/LI2qIJY3Ix65+XgInrpsL4M2L6Uxy0V5jmXlkZwCd1TsbN
lJAsfvzS0pK1kwQKDLkgghe5ZssHbHZRKg1PID5EQQTfzf5cIeJlSk86xLHZOGzqikeeJ1et3oEv
moR4PpdoZXFRbPD+fewEADNRFtuL0dfIXsgp4Nlb1Ghl3bJfvPBqFc7AufWyMqaQzXbkxF9Hh1fc
0BcRETTYyPYkXfB+LlsqbaaUv6LOgYzAohMYp798a45a0fpBoLR/UXl6lDv5Ot6a5oNajxTpjelZ
j/ButE9ljZ4ZTzvnHcDddr8oagdC2LY8HrxGskC3fkys5fQn42WX118uboPxjQ2lAviUNrtkgfa2
FMkI2Vk6j5pN6ws3zBeHo93WNHd4sJyGJ/q58Wq7mI0xg2NNw/1idEYDOJwn4jI5VDzWxYiEQPNr
u7aJrHmQLOHu4gMjO1KFoOQ+zlLQw8l4MneJLMvNC91rtrdXEjNLQ4M4vvfmDfHERjrPJVMKfiCg
CmqHWqWkrX3lZkxLXLSWLJ3p1EfrtV8Wra9V8saNSkmYcIbra9v8hrRw4v9WZiglO1g/1z3AomFD
IQM64H5pVuJP971qTNUeEB3eYc2lr0p0bjqhhh5utlDdxHJQRjQMEp1ZvjT6Xn9nMoQGsG23DjU3
1oU9tzrMqBkonhNAFgTd4N0mY4PkypcJ9E8IYCv4J/CfDWKA829wNjz3zZsSZ9CKtzUxD9PbYLJ0
aQTUOlj7Uut9eFfRKD7B8tK4WKTBwGfZ0T1x+PbP2HFb26wFWKoEZOGE5O+jVLdJzBpEUUgPQOLa
yXXDkVJml0q5prVmPlkqtX8+hKxmZV8hiBHXSX5YTtbRgaDdm74OwyPAd+hrWlA4cRloDof5zpLx
T9vVlIs/VV6fGTgS2IVBrfs86J3v/2gUH8F5ymOpaLKDHYXxk8roDqVDvNAxBbGUXUtk8uYViaV8
Cd52wpbf9cuhE8j5yidi8g377xvpDx+fcqXGN+EMi7BR3L6Um5GbulBQmyekAozBSxVnDe+fkc6R
+abvGHLxiTrYuVxmeukfzvNnFVHdgYSlmlWveE32wQ0QkBMAvQC+bbbSxmjIey3m1/A2ACTeLcnQ
8jhWLh0kofHql9ZiT9HDERq+FjJ3Wjf4SQ89ZP8NJeHGsOElS1BbX7+FkBa92ggTHvmAO7oMEfaf
EcH1QsW2gJrSOYLouTBTzhAEvLwcg5XUelPBDkwDL5E8hQ06Ne7y+lE+Q6y4LTJcGaxONrSM71Q3
KVoVtU4d3PkNBeBJgmFmPTC/8kOqkgQEfyXqAS4FklruO7+4r99whKhlbnhYih6RsRpOewIq1RNP
JdQgNxVZO6Z9U0u1ph1BwRKcET+Dow1nw67SV9xrcRvhhq7F5Q+6JegIliUeJp5+t1ABToNopqHq
DF14W5XwZ7652kheD7MBPwa29QCZTM5VSei8B1xLGKbBe9or73W+c99L7sVEFZgROVxD14daOJUU
G37Juq8KHdoceJiDirWDMEaY7iThP1NbiCJ/H0oY5LIQzYfKze/szYUJ27Emcdq2Tbn3Yq8FHN6S
Od826cscYNKzOmZFGgeou4m2CLWmnnQ5hzhWPAtORcm7BFaxnd8Y6ZPahL3cVnemKoZc6V9AwQCl
2Drg66Yj5e5zXbRxBgcv9J9YFK/RSwIiHrOac7RKeecQ/eTMCOKiA6TCqfQ+IDpzWAFwEIdVnJI0
BR3QFpdAcFI6e9Q0F+mXlGrAlKNtb9G9DbYSNk1oTfvZjhu6ap1L3L4KYC89hXQilgLgIVPV/7FD
UgzVZimLBn5i1R5m9u0pIOvPn0QpmczqIgBm9Yx1/sJJWgKqIbill3tYPA3DfkDRWksHS5psyZEE
+rRbHy1sQRyG+HH2yCHMYlGDPgDz9SXirWrchhJbeJR4YXf/TXNOfzFA3Kw9K8ZGyikUxpade+7t
jFkWJyx4BVidf85TODFkQn5VyDq+21Gv76VbQn1ELIV2Sjw6m+9+LcFXyyJElTndhnpyS08I4ruW
KvunACwVeC23BjEy2BjC+9o8kAGJ5aA5hyRIvfivTbZJYuLih6FSuf617X30mil8hgdVd3RDsFme
6TBxsIxmeeEE5zU7tOu5gEsMklHCovRW1ej7Zcm2daIMG4+k7RLxYP3Qu/QhqQ5aQH9IKAB1pMZx
UsOlppcEYHeUAbUM0aMbrapvgnJiWUGNF1UpzFxgzAnU/CxGsoxspifBjnWot63MywpRBwY1iGPt
hWzwnhkkDLVmou8EapJEjIvFf573+lcXuqe1ekSR7InDpdRVgetDotQ2WiF8fTlSh4lTU4tor2Wx
bbfBuVvpA6IaZzZFYgA7RDYWQ9DfDkM+2ab2V0XRBqioYwTqsKz50o8y5V2mwdpZYCgARNl8ptDY
sBkNBMKVXSET0fbcVQgXIekTZZ6Tgaloa+3rOqsC6xffQFlB4O+QsnYrhpddhPoZAtv6qnBYWnrg
JYII4/IXrx5F5tlZfK2rwvygxWHquRZMDzK1d3mjf9iuisEUxAPlks9UpuEFFqYUrm2p/rYpTBF0
7I7D4ea7oRoGejmGYyJV9IPWFpeLTp5tr65n3kH5tcZMUJKmnH/btkn52e8wqqnHAs52LHPZDqsD
QCGfjfqrxzfI70J+qcAddWdEjYBjOX74BnDMx3L+e+Y3FI+SUIlAddimZq9j7Ief9w3/Iyz+Ywqv
hWbnx+nkHTMmIA/VIBLB1h4Bi9MKQQwE6IJRbQIhj4/UGp2yX4jLtUg+XRMJmCgz6QmfDCyGVTVm
ANnUMbd6Q0fftGaOYTZz6nCr960DTDav6rvs9XX33exW2pZloTWgjoBD8QpxnFbOMSsVsOxnHQOT
S0HqGwHjvuPkp40jkQQHmLQXvpHWJVME4jj1xNRfvsLfpG9hscEfffhzYRd0A1ZAROgOcNSfoxIl
hErh9RViMg6/l/p4DHDxIM3V9lWrvIdM3MuPwqRFsCj0LQaIfSNjAuMAC+uzMpyEDCd1U41B+vhy
SqcoDOtFYD2pkl41Qzv2A9d/u4PULOsGRcWN9n4/y+2iX8fM3nWelFmu3U5KlJPwBhR03Q6KF5xu
vSqgSOLwTswMd7qg9cDwk0l1haGG0YEv3jTqQqHGpcPCYVziuZerd2mFSjunPWd01MjQDnCczcGj
TOyXQa4+Z60UNtd5wH1Aj8efjnnFpwQ91L7+AbqSc3Sr4/Y0A9VdHtncSnF4+UGEe7lkmp4y6LZh
LrI9vKep+rA9rwhx6zMQMzptYUG3fU4XlQDugSP/G5XULMdDDJwhERnK2N7XfQ7IHab3a2+J2BXi
Ld+EjTOPIKZ0sFg/G0gLDNJJN5JDHGEJY7EyH/78FMmEQxRTjU+lNQ4jkW7uPQd0I9tBi2XKXvTO
EBvrEa5oezvOhPOtmiARCGFcL8zeqCw94M6bQEy4NNaiI0FrcL0JyfX6oMPmjhza5TfsS2ZmDmc6
BYeBPOsmtPR4WYe71MPu2d2zmDD/0h9BCi/gfQx0DS2iJ4Ye8tK2Pl01HFiLsl+Oa5xzJMqu5lO0
fyMjwdX+3YjvTc/SpBTtno+RY25ZitM3YocRW/56aKPvj3WFA9PBO2I/u1q/kllSrCI2mpSzOAn8
Z1RC/uxNdAljn0sfRs1k5BT0QmTqIBBkmWGEqZM6M0b9BVugQFtd1Fx83nHTzc80oCdYWum9R8TU
lBTHFjQM6+CinC7JlfjgQyS7aufcLTwxil068vP2nvYy+Z3Lqe6+6zGbmR5A+BXmZn2luG8Lpn5G
meBhY6xL98ma6A7NX4koJg0A55TgcLhQi6NDeVizpbkGRvCt/y2P70FrzrQ1qwSJ/tbw1vTSQwGW
kTAHRN7RxI4jwrx+2Cl4Y9TGpw3ik7F9O6LQCiellRKE8XswZ0cKumk0O3y3AoHXqWR95DydfOUN
Bt8uaDlFJktvqGSFEKY6gA60WKw74XhfcNjmbu59Etkz8I9HPS6Xseg0yOwe0ikp9sZWvgXEV/+D
w9kH3W1fSmMSm+HhZO+OeIop049STGguKgj7DwoHrnL7Bn86gwnvRO55M4nLRY3Y1F8Aj1w0JTQ2
i94PEEpsLgovRNsmFNhdnkeXZJw8ZjApyw9RxzjBwQfWTU1gYFgR94iMgnq3Ho3T9jBcBBY38o0F
DcLdKfCIh0FYTheBKsFXgzjch1uBnXo6kOhCAFCRPCvQDIb2baoEzry4LPjApaLP/LDHynNUowmV
mAUxOyqwM1DIM9nV6TXa4crFM2Yl/J3PzInPwbF0kCkvQjQPlOSPp4OBiERG7/N90DDu/PVnEqkY
+giDaObhDW8nV/FVU3yl0AMWWY0jS9YsrUGki9CAXfHCzih7Uivb8HYltAP4DVkn/2PLYFNcaytz
ZAzQZSmzj5kDTZBn6Ntla1SdlWcguV7jkh4mdlXuGZtsjJYchwkPz/laXOgqR00kuuH5imaqYg7z
vcAs01d30F0oMHWg0Y2sPO3BbUEhtZKmTbmJjqEkz3kzc3jRgXiiv4Z4h4mAtoYvRvHiYAOAm4T2
3JdVk1VH+xn2mc5zcmcCQqTp3K9V6qN7l0t9QkHIvd/3R5kDJfWVRJjWXZnLFsnYDR5EKdce7Fpu
0PutoZwLhBaBqqM2mIZRFzh8f7eaxKfvuxUgZL5HAYWbPlnmKuyAGWAd4ICv1l04hPGuX5smDhjI
yQhYiObMY2PcQU4ejrBS/VNokhwMVOlyQ+XEwKOND36TdqPyoU/MHQA8oJAZMw7v6PoaAxA2XKXC
Ykce/pVnPyHhYgSL/7fBkGeW8ogV9SgCa7gORImzBNXtjzFv+eFwBni5p4mFffr6Gb/9M/v0j5Vw
7y1ie4InqrwvTCdMvTB1BM89URuW6R35Z6xKz9qIWZLlrfL/hvGBXKe/X6JGu2M5edwDG6mp/Jp4
DXcWYxxE0sYQTDa/Ic9rmIT3jQ5NyAdwsGS6N3byYxPJJiXVpiCC0ZFgUs02NCBQTfbIVPbkUqPe
clQEkhvf/GtOp9Fh0J7yKE6vy00u2tCw/wtExba82Kz5UUK3NnBJLxFj9V3QxivRGLH10yNaBNin
5TXiOHEXD//8sCQBZ2aiJ3NasObVIlT5bol604QPzdBZX8BdLtwJrT0Nc8juXWsnKOfNFGVzwV/D
ZGFBerU+9oMf+5udzJvzzINGzC5o+bzxaOqAtKbmhRWtyJniwsXTJ8aTFObXDJi+r87zH4UToDO7
5nQUS3R0oVrGXwxpBgtSy3ZkRJUbWroIMqrBM5kJB3VRxvvEf9FNn8IG58Bw3gBf6IdVfTGIGn52
ZWzdJPmDTlvnE6eWnt1QXCNhxmffREZICxMh/ZDdk6tYxCgbzG213uVR2VAVKvoKLUH3XG27Ofis
xrL5kwMhoWR61yFDztxmKamCPYFUwRDK7RQE53JhdqPRny8wxF9gXlbR4Zc8nxDw0IT/0bgwBlhM
inraMYtC1C3TCGnm+82yzWyHZAFTu08M9JZcg/Mm4gw5xG8X02/3ZhYqNJoajyO5YHbvh/1GrJde
otsiSiel3gaGfjZQiVqxwDyDufmdpxZNpjxSAE/4ZWzxyMBxGl38LnHJ4y+C8Dmc+1pAA6waqmGZ
dTf/WcbWmlfxa0cwXa+djs+qYh0U0s0I2NSpizJu4BSTC+x+6DSyj7hF1SAwrpq+NugF3RlEFTWx
R9c1CGIX+w+xFwWLNePG400tUtCO7SuiphesLzEp86SOfLHnGycXl/D2dmBI7rHq3nTFXg2azkTr
lSkA4ZDT8p+oGAJCa/tFEWQlasqfB5LkHNo+fUJMf1nRYJOa+2Wg9fBtYHql33CBxBuZhsMuNIGP
xb5RejaARWDJD+UEMUI6AecUeDlSNkkj1lDlde8C5N8s/eIOc01kb+ktMNsxghJoZakEPaWhedNR
oDWM9WaF4rHXB53a6XnmeBng+DZvHql+4DWQuXEVlz/Arq66Suxyj5irvQ8vAfTi9/3G5oZkNeSA
rDExC8NLHwPkhetHrkltb4T9rpmXmbum7KQie47bJI0bO6S8xZUJIp2k/I0SOQ1O05MDI82J+XKf
n66vdbAJ7BhLqD0WPlijdQuP7TEYS15aZeHx0vXeb0H85srpbdbp2nJVWM1qR74kCBVAUPFcwrU3
XcVGZk2rCqiiIg3bzVQmwNuEIwZiKJ8zVp+ZjeYxRxbNa2DCmA0Dw0wZg+dPG4NnIWA79uX5s+fW
qbm4KrGsIllUZyYtgAgY1c/ClXsqBH5aO5rtdSksxOJfivCqlJrNqKLYi/nDLwJyCEc/EPRClrSr
gkNuXveM50qb7XyGbdpaEODvHjhwxK9R7IPYLsy6b35YAYTr3vZWIuXnZ6jGe0zxRAvwDYkO4qF1
PXp5G2NTYidy7DrG80YVziNsJFbELP1rjAea9VaU6j69bCTJpcCnYvRRQEKO7Yd5H1YdL2jCtSvj
TFiB0LG8HyuTOCFZVfokQhe8UaI+AlsscwTlxc7sgucd2V2GVf5+7sGK142bNkWb1zcJgNj0GUVS
PKhDEDOrpiinngj85KElWCBNO+BEhd+1qkFX+DIen3PkJXWLOE8p0DcvvyHRF4JjQazX/msbIzbf
zShDFeafThOx0ZHQ+RGSeBpzK3H3pf1LXP2LLBK+c8NhWL0CGBluG7TwusgrM+g8SvI4WHC+emSm
UzH+gtDrfyRrNPUFvu/EIAO7y3UWFO1yPaasysas6lmXbLcBxeAZx8w+abiPoMh2iN6MVYiJDQYO
qUgK/S8B/5rTt1hAVblWViF6LUdtToq3V/r2xx4z5di5Vw6nARtTXrGGAmFzG6OxFmda7qanVeee
ygCRWX9U0jP2B9sNZ2pKYMkMqNMnSytT2hqbrGmREvRn+HZN07DwGhbSYFBfG7qOChwHxmQsdbS3
Q+arXhY3cvBuD07sQe2qCj5g/p7p8Blm/L2sxganCgKe9n/cKg5uepy4u4Kw8S2qeltUxXmWsvrz
YTKa/9f+l+t/gF1NoHU/+s/l9Iepy1Jd76MB8mYwF23eJNz3Z7ZukiJLJFkwzo+YeDeC4TkaxqA+
BUBtKF/TLH0W8F3NP3inYbz7gimOS69nDBeYKYXR+OD6lNryY8sJYa/cDcTJhUkcdkzNAiJtMEUR
TWF4uPQY1KcKFku82bdvtDS0cVE/qEwDIKqv825Puhxr/nLG36Lv6AzrRrIv04GwdCOaLvM46EC3
ns3xTWq4i9Jjog+0wQcDY5pNhJQqz2X+JHTNDwRwujt07EbQQqdnDLoqU04E9OBhkV0POfz8NS7c
DCPdcE+PN/Cv7/q2kwN5ShN7ZCl61kvF2EnjR7r57C72ic3nmFS7x95bFg5QioMHKbl719S0Wd3+
VsT8+zHBNjaWjKCngUTIXQM8XBaEIm2QxzHCB+ftf47t0RCy0eGH/CfiFLZzXoH0oHUwwY3znP7y
IdhFvZf62oL1zy/6aqkwYN1TZGwt4B9boHFAkc5iaHzHXJL7rauom5srvTQm2G8EY5I8Eo5LxAup
/eNLCyzsdzMfamlwjbpqPx97/xJJKhpiWDewD6Gqjo1qjKH6trYoi4pFK5k5Zo1X+pbSa+FwyyAE
IFsR2gRP9dJU4bodKlkliSPwKtZR0luua5Y4jOs1Bzj30+4uxIgvSbiffVAvTi6EH1yhsMbEDN7a
+5g7sTPLaC3JOwHcV/df27NgVsMzBFLsATtlh3OGbwa1rcxTtG+/pRzQVOozPtnHS6Iwy2NYoWcZ
rKwxaCn44RuD/v5JMpxlNsDat2MKp1HE/PQ5P9weyNGqBCS+e4pN1T9YYWxuCjtnvt7tjmdH+hBI
Ov6HodSoW2U32/LB7v/61uKH+SNlN4yPbqjp9LudK5S6E68H/ImwfYRN55/kvfg8oQGjDFIVMEsv
ZvfYyDqsna2VCoul5edM2FuRzocjY6XyURmjBfBVOdO+w+c6+UKMWyv0Fgx6Zl8g0liYC6+c5kHf
TfKn37TZ7bDHCCeXhgfGzrIYnhFv8MifG/oMV43xTuCuhR7S8UfZpKxfY3GSXFG7N+kW1FzmDTRs
QVxL/7ycSnE2wEJs2OFKYgWW/9evheuLN7KZE1VqnS6JKmPsyZXSxay3D9poi9NTj/l4fRoGVq2m
ozSXTVSTz8oK1zyA3QfHtA7zarDdaiJSTR4QjLHPPKjFzieBNxZSoWJAWVd+/nrMIUvuSu17lZRw
LmfT6nf+cRtr0pOTlXcTAHl6VxcMWy2zeKGlkxBbci8Do5iroEAikrknA/NWmCTg9v8AsRnRIc7G
NMaX8xumFkNCDAidjYj7Qpl5u+TXYWKqg5oFg3NQugRsReISs/NLJEvN7J2PHki8zzBW+96fZxOh
Ujg5r1b5JhYvjiPrcTkzv78vqg2zAqy6qfHDis3jM2eTKy2PGTNLdVNmf5q0LYfYCtcxl4wa/IrY
MaiZG4LD6GYMgg4b2gDlXmWRTwkOsBnkmmd7WLoO5/CYbrEiPCu2mUkojzY2eLpeenAtgxeL+A4r
ck/lRwb88Tc6w4Ay9qUKJvPm0D/OLewb1Qa410ZBkSdgLvaMAPE7YW1u7OwZHuG5RorBuANKPWK2
pTBLKcdgWVlNuEH/SIciXfO1JMo/OOzB1+t4LXLcoKNQGUmh1pYZU/jCoKKq3qwQMi4jqp8uMJ7o
iZ9k1R9YBbyM5A3CENM3Fi7SwAMhC7smHY/GiJxuCiTxKfE7vDdwio9HAXLpZA7FC6me2fX8EAEy
KDpq46KyaZx4RI9a+oXKhvThmfgopw1uzFK8G7cXtfXZCYrqueK17ejIef8B4AvYozJRca1Az4fu
/oEw2f2MMV3aQ81T2iR1jkfqVV4DX0x1YNiWbwroXUyz1bypdfVemLySbpbvR2nlv5X32DNJcPhs
d/fc/kAO51PvhLaH8slt/eztOaley2Z2cAhYECNtjwoKbnFJ8j2ByNCwKkhsmiUnrUK0C6YqK521
ZKWLQxMCo2sEDVc7ngS8r1zZxEJsEh07VCYJiVjACTdMAzhWVAvNFC7XrzLjtyeUO502U3dCJ/JE
iLQfmMFX5Z95Q2qOVLBKQNvFUglBs6U25V4co0WBusBmW1AaPhtkgNpsFAnlhNB2OVMBi7gQunm2
DvA+ORw7oatBXPmYYvGpt1xJXr38+vO+HbFyZQKaHkwQSqXaMqT3s7ixGbXORcZz/NasCP1P1Oo7
tYKw5kYxk+N4UVtggyJV82vJ7Km+DF46TRQJPNFxI5+tbyExP+7HeB9RyDzKZF1r/7sYy8/6Ilwp
+qBW3OwwAICaeCdeAZ4yvTKYZaH9gEFNeenRLrhsxrN1WTzLbTSZuxpmCs0hHkRyo1qs1NeBX0fx
8AglyQ1kV3C2R+ap6Tb2L6vZPn0feb50INNVESghnZYnSS0qZV4vlZVIlvokufhjJr/77FMfR+gi
yvAwedA7KmRrbguQ66ZIvcQIQkr0pdj7vymBF0v7pY8YXbOP7rchqa6BjbUhCH0krogAXDom6vu2
/IgodqyiRrzwRlzDl2C9+wQRXPp2Ot6gkB9NXprIhwRCjQhwXl13UFYHDZ8GfZrkjm7rJhgN2YgO
dmrGbHKiOAWktiSR5VQTMyHrASGb7daKiX7Ojx6C5OTI2MUYFYHJIKBRfvj23iFCMLapyrJMiLSE
6UBBme2W6EusGPfiBIK3jOiUS76gs/CN63rjT/vc3+qZwOVV1vErHjZpLJCJ7dILAaeX+ucKyHyy
HAU3y0QN1isTJFc34MxXN3MdDhvj5lb/nMrO6SJ+7vkHDKK/hGW2xZItMwtZ2iu4KWoDQPPPQFxK
00C77cJ4o3wIwowqVDsazlNwbvL7gtvG5awHHVe3cCleXlV2qRdNqVDahnwYF5mlMlv8qW3RbgN2
1feJxQyS2NcQSxWIBlBqChj93MasPL/vUu1OP3RBPMcamH4NS2H3uidKqShGz+a2J/qatrX6DVlK
NVKFTAEqKYwocYiPuul4M7oZg/xWcAAWnCPn4LJlQXx08+BEdCN7dWjSLC5iuitOCB7tdbsS+99n
ld5ezwxFvgFrr9noQ/bc1txwFaBQZZ4JgMh2POQfbGNfxaZIRO7eVQsRemjgEiK+Ke9jxS3hJCGq
DVEkR2Vm2mEd9vn6e3EBWx3eNqD4dR1yGYUOtULEmMp/cl/GhDSO1nUTITEAHN5k3Zxv1XBbv5qT
Te4NebmdE/fzOWxiJEMxzr3Ymm8xZENklT2t2BVZMjwofeo+6O6D8l3Q77M3IJ/tUOnroilAdIAu
qRl+yvXPCj7WqnwjbAuttFo8/gVTBZMKB/DnSsAevGw250xdyRY6d1fTJxl/tT+SeLCH+BMy7fH9
Q0EZiABrSsTs0UXwvhjCSpv3WhUjKh9HYJzKU5rUEMIKVvgShoKbHvjJtkgBzR/IDWS9wMVMXK3N
9t7VEVCnIBKljzJuFplzq9HsKa+MV+jRYrF0w6kiVhocRfKkRtQwuOJSZYAltEcGu6hpgjfc8P82
Xo4c5ldosKmNHclM+Nk7/6FfSgaVK4Wdc39LnY86eTKsX/8rmYJqgxjJqVUUENKXxt1mScFHHNeg
MRisai/cM+vI+SbTcPZA4CiFEpj52FbsoPzYRjmS/zI0Q6/zUVPAbq9BMYg9cydDNRViC9Lg3jHF
go9sb238yOS7aXM3QF+ef6pm4D3UhONAkB7fO4qc3x8ldO6sPDWEJ7J6Du74j3Ci9KRCUTPNK2KZ
SL/DxD0Z4j8RAP62A0nUhBEzJL2L8YXy69ptqxQ4hsbw16VQGerJvDTTRFtAwFXyv5XZN/NTrbgw
ag7VUBwIMPjoqih8VcO5Iw3ovQqf8JT0kH68JKqsH8GXFcHbK6um0xrAxYt0rY0MD6LrtaQKq5zH
eRN/z4FGvEHOdytrc36oHutuGsP4FxufaiRjI3VL2+8VrAd4Zr3O55/iRvNHzW9bHkE2Mw922SLy
HN19efo9aQ/eqLRpHOpmq969DeBS7qaYFbR1Ubfuj8UdE5C8VNZ1ujSnD+v9khIfdGB64I/9D2Kk
nCXSte1JMOkSo2ibC2JPZq5A8E0vLKwB7ojKYqVZuR4Lc6pKsV2dIP7MKQZI3EyCuJ1+xGATRwTE
wCaumpaq7eroztq6ijPuW2Ouc4UaBE0/mcm9XA/WUDac+QQUCWzUEhZrVA5xM3r4ZBwW/g+7fv3e
DmCTSstXdQ25/ueyC/bY7Ip4tidZbMFBMBBJpSSOUIqAbjANAhiaxDotBTyneEyGxYCSn5sJqAdd
5n3b5RjkT4g1vAjquDBa8yGqR94Xee5KDOTBMnF2VebK+rGx5spkhEfFRIEQhknoCs1s5dn8dhE8
Ij+QmVYkm50MWOQudEFIQElprLl4dFQ1NN6JRg6sUKDB9UaOOO4JMOHOyqfrg1PAMfVHgDFL001d
uu6Tru4tSfzKyFp8u0T3jTP/+owGHvr4b/p+dvQaDkFU+S3oyYYJcbZMlBlfHvAydB/yBN4xmLIP
qhp2cbwnvepshXTQIRTwT5yExefyHxz4vvC3eWBWOyE2BKO/ZWvs9+7lLAyhscmqpmVa07yrCSeH
gL00AXdUxmc7RX7OArS0N+8IIYGv4iFi+QsljRdSkakhL/mBsZVVcfBh4L2r1TzAxkGdnZx4+i2p
zcHculKvqXJbM3FTD4YpfMaZx+B/V6ENZPzPCbREYhEYvlXIV3SoMkPS+jdw+gHoUsG6/CZbPK1s
K1BYmseslk+iPjcqZanhZa7w387S1nviUtjF7m0HfIOrNBX8ztVKdjtqak+/wZAoU13u7PJM43iR
j358gsBlsx0bHHkecb1A8JsfensN2aysXIiGEQ9Xcoul4NGbj9kjwCa8dv4f6Q2AtxIbIuljCmxn
SAmbEOQ8DqZyp00LUKJtXy/wBcTAj7XBvTztVf6kp2ynX2gfDaArT33mdl51sRj6wV1QO0CsAKdG
A2oo+1DtRDFUDUpAk3aTkQi29H0dqcjEe77VEb0NcoMLJSxkywGjF8zrX8MagxC6qXUYeuh6bDJ8
DVmhO2i2TkJ144oHeJVwep35W4D711uNuhcN+pzdCdoizoJa+l2p8zUbYWPI3hy3dSsQZESIGSjD
QfDseeoVCqu0IuG5GbU7CHvuP3E9ptKRGFWGuxYxDxRuIL76SvvmUmMAiBQJMhmIThKXF6fFk0TR
/uj5QYDHiSE+imPcZ3I2XKm7u2jz2uo60rHq/m1wsdEiR6MDlu3A4Jv6uRoMhtHlqZ7ZdK/r3Nux
GzpO76fICxaLCO8ZL6t40e/bZzyWwfCLnl659Q0X4nklLRXBipALOUvAHsYBYExQV2ZTlxO0Uow7
OdDkw7B8QKLKfflEpZUrjOvbYiiUsSUoyEDR2PWhAgMHnbeEbWDeNwPUYXURJeaYGbagxOwdrcP2
AoznrChPPmI+wz4iqwdI5hzNsX/H7zI0MG7xSqnLr677GBGdYQN66/uooxbIGePqeTKithBR+Y+s
q1OdG4QvxaBCuUtAfKpMUgQt+Ul3ezSLCuf+FdzzSymLthar/HCaA6ZTQKtqBbtTgAOzgmZPaIeF
Z6QMBQVUdez1r9tWERKSDem0ujz72HGA+ttjTuR+OKkJg8q5dHcc5yJ2jBAEDHb019bXvoNpAPaE
X61rjroYnbPEOWhCPzrpiznGc9+NfDNpI2dNqv8LxAoKni/j/WfPttwv5nKWJbuVEdcEU0G/qsJr
4t+VzH8Q0jxb4C4tSO9Y9JgQzwFqv25dtJ5H4vmrh6RwJa7sxayYDb9pgv4BADfxfG1xBkaMLxBe
WWH8N62kBT7ZYSRBg56K11yZSIAiAOLESwQtrVrs1SN8VlpYsGabnmWyVwil7OsLeA7lvDjMEtrU
80jz5lGkEGE9DAd1XKnFMwAM9lFVhTcYh0YDwFFIBjEAIdZXHvittuJk/lM8C7ESm/Ql4b/9WCD5
w9BzixDk85G2yppssD1oPG+835QIY09GfwsaZX3x8fpes5/FEYC13SYtBZAFw/hDRs6ODhzYEpLC
3n6987QER6/WbmaLu0QcYVfE32lViBjRFMG6MqK9qDqDTW/aBBUOxkwhHcwCCpWYc5XgB0h6IJ1p
Zpdr6cMkNexq809pg5EuRKBH0WBrwox8Weq8jL6HIPqzB/MH7W6LHJQf0ZJwYHVW8c8nG8s+C2NL
BRpgY5Ro10jfc2IamWpwMJ+yr+5rygpeQ5ADhogOSOTD9jfQOkgyBGSHxogp0shBQ16Kknhxef1o
qbh7CD9NtFo1KdLQtMa2AXdUQ/iRJDoxCCxDNmUdBKuYf9F5LZ22IdNCS4O2kkFFRARZvq2ToKof
etaBvwFAZEAhzzvG3Obehsx0tsDuSq9wOcpH9x/4gZkuE9siCmzc6lm533O0/PtPKrudgePMYO7I
3u2pEyC4B1I8nDceRoyQkkaQWI7sc+bS5jX9tH3LtXi68PPyVzhM521FNi6psMStqagBh3HfcPnb
8bRegKVqBR2hjiMTN+I29tGajmOEOF6EYoKjxMLhMnAJom69KB84SRIHX4MZGGA+pQmmLAJ3WHBo
BPOC4q+EzwGQcebmV2X4jjz0Mwk274OOsSCuSM32lAQpgQZpgOuQJgazYVPXgGAJkawfPB11nyIq
8Q37nguEi/xOT1oQ2iXgOPahzwiEpLLPYf9qg7VYqqvyH2je5IqAMsZR3aovvBbfsaWnd8Dt8fkK
QzF0DvL9Xe2021fR9QKLUT/QEHgm9D3aV6wGQOe3GLoteFLFIuChA0Gyo4I+ZIJ2sFRVBpF53DnD
XjJODI8oO5iv7HRJM/qgpF4caRtkdffAUer5zpQc0MOklUBc2HJW/iTda505jfAzKnIl8JKZHIsq
C6muV+VXrp0xnNH+4QyY4ar08dyHk/8Wkvn2XaZQ8WHz0lZdVAq1Q/tlQIT3JBqkfChEDmCisLz2
hIcLCT8f0O++Vy/bnw7KrvX4QCAIMHFdMhgvcabBq0GAUtt9V/kWIgSO0HK9EafRD12WDCGkRHIP
H0l5ynomsANbz5vzYgly6+rZk2rXDNtUosFXIf/sBKdxmWLQwl6rSCPQpmSgz0tWPSImU7snntDq
Pix4vxgZaOqtuZs6MBmyTqLIiKIkvVNNobuIEtLachA6u+Dk+sAHozUbF5E8IQOH98m5kK7H4fcd
h3nvUxJb5Izo0Xb2oM3jF63hvsfMfBDJCj/9XkuhyidfQkWe9Uf+atHWyjs1JlvhCOGJJPAnetXu
Lj+letJ5aTk5rCUUH4bHj+ZP4KU2p7b1OZnDPsplT5Ddc/ka118h6hIVa3QSVHFCp/IRkTkyavRc
Vvz+OMlxWEWHm4zzNEZVG1nIR/VjQkDNYW6uZMKEXcw/EExgzY4Hjz6uwdnOImDyfuEpBarQo7kB
XCbMxmVNYHVjdRsyPo8Nd9mbBGQh4YhqM3B1IZnLUsXh+fu8BIBi0kVdS648gnaj9NSiG8hYqYKA
FWiu8kVPHF1poBXOrKq6RJM6GS1n9wYCuGwA7Yc9ZSgSBSKGEqiEAg+ZogIaZyep5CkSz2EG6IbC
DQC5/QJO2djaXJaLwmL3gfo9cHBXETfRXQ6twM8vy+tqf2e0rAlPvxOgM8psb3GpC2mYswMYgjrY
eutnMno7tte0oVkeuK0PsRQAvMIAx58lzBRyAeYl/6NHeGLOaqMFNNHd9WjkQghCMzGdtXl4uiko
CHNWjuW+3EJKiOdlFWH1nmUSANuJ1s5Zts5yEj1lkK2BnuceLPlw/jVoBb9rGefNaW1hsuG6snZT
1xMg0D5i4hn//QV8QKAdjbZU0KuWDkoDIDT69MfvApapinCfThjCymxpP0GGybFU44+pPQqOLx2Q
sUI0WYDjT/KoOXuVkJXOWKA97MzP+tYD3/OTxdx1Iq1IDrvaOy1e2bbRm7002ADhT3kxcFVgk6R8
9G85a66qEFKmWFZYSXekNSqnTkxh0GZyBTg1yHvGY4DF+4HpI2NANFOQe9Su9lppzCGyw72hT+Av
KZ1RFmClU7jB2t/+wmxzEp/hFStbfatGTGQ6bW+q0KH2gI/ssqS2XDFF3LEeZL3apAHRpI305ZxD
8NS5kurobxD05eaKRriMTS5AHb7CsB9GRwlZbVPRbsBTigLl+hu2RhPyMTdxQfGSR40iG34p37m+
8Z4zqS2KwR4fzsNgl9fr0JiSN8ZLb74sgt7xzk/JRO5OqFyPuo4wmsTWUJPx8jFO57wNSI0e7Joo
4uZBFCUOGm0b0P7xbqSQJr4M9wVyKIXQ/Df5QWPZFT5fiB4tsWnDNeHVdH/23q5fNMI+I/s3Zwo2
wiqWpGB2xeH1CJM4hm0OZXDmWk5HeVxInHXoG1XUcmkO/5487LYdcKoBepj0doLU6mo8i6uvjrxS
20cKRN/XS12yT7koJ64wYPPfJLZc2ZY2sxbxcYZq2Oika8Yax5SyxSdH7yCtGC+0J/xFxQvY1l7f
Q5GxOVEXcVkoFtEV4Z40nQjlkvDvUhj++7jmK173867Y/Ke4SRSTpS4p24jroULqsC45jaV5Vd0n
Yd1iLZE0YXQPVLqJdLFp9xFssoWiTXmSW730ez7s86wRDVFPdUxuGMNrnGFl16BksttKtJcblOPu
pDy3BKkfIjTCAkKpQJ8hARiGrZ29e93ecgkZlEbhAP1upz54lqJ62w6K7kWAZAIXzn1cldFQeXcN
1f7XcuAj/RzdyLlPgDYVbT+MuxPTsrSNdhld+ozcOlooYtP4TF6A+mMcjPL0MLyl2OPcDarK3OD7
g5czU1Gci2KhVLdo329ifeSxNJkeJ4/DfLyn9jH3Sd4DUnRisKw4E17h+OfvGRtdl45nbud2UJTN
L4sWgVPSt7llu18AQMQ/M64KLQNZEAShRgKP16E50V4sj0mMrsRTTVNbtQtWscLPrvod1cVtOsZD
nOZ/L4DQYwWckRn+E1ksL2mW/tABk1n9TCrBKTC+q6h3bKjdEp8GE1uMLVvqkiPn6qDfuXw1QT9/
/bNiS9bRkUbiwW98OHiGlwXo8Dks/LFfpw+EUKnPDH3coUH45tmGW397oAA1BFSVQilLYOkviC3f
xbM6O4i+RsYSD3IUkhtpicYpxC9FmOgjvkOWj9+itBS13HQAkUnNxkqS6aaWYi6qrvMxAUESJlmf
U0Q4uNyPwUWoFR3D8yIX2vn6dNBvi1YBK1zvJlsySD3kIVUOGOpFiBnpgN7I+GNuSByJB/5Pv7A2
LVXNl6tbOQuv43g0xsqBnO7fQWS4CocCFyxKKkdmj45lygSCdysXMf8aShqHjZXkDlUImaqKK6wW
WZ7gow7Ts6w6qYQCk96A2r22OV+XzucR05K5GSLXVtY/1mhcWXMRu9QxswyjstuNmDEq0y2T6L+K
C90ZLiIewl4pDgMaWdM9QCkEarOESkt3QnzJFVGedQsIoXEdUMi+flghunMc+7QXemUltBofxp+I
U0jFJqHhCA5MlkfkxhUX+dnVHvhIL3zgmyC/jB9QVE2gvfeaoajXkyGUWRsfFVTksA3gSjXeZgDf
4O95T3V1v196LiZH8K/eUUW/maUSfJUZg5kwNxLdgC6LnUZLhF9I9dpXsordKpnmRzo4gWYKmxzh
7dGOlQ9sbgwCKtEONXHpox+LlKh/W66vx6HKkb3xXVzFaLrd0kZr2cnbfU7wiyTLXlwFsZ/zEr67
FExltGPsA0mWaouKBs5TA2J5JL/hHEjaEek+bD57eLQsyO/mX2112XERpfVuoMTtYba1qhA331kf
a0vkQYMvr/U4tugeFEGgkbHOdK/cCdJuaUSkDJfN5JWXfMSAJEIWCxPK9dpeDes6Ud1PiCi6xppf
V61f4pu8c8wUjL78FYzNkb1h0NVa0g2bR6eqYo5ba6UUOa2d91h5gjaPgJIDJFNRGKh6JcgsLycW
I4Iw5Ubiqf3FWHPbkOAqMqlDrrjxxG8uHhAl+/5t25bVVxpB7VAEFmtWRvsUo9eqk5isqlnJC7U6
VTRHhtvJE0DCAJvENRGbWbDMWUjlXxmE/4jrd98GF/XL71Fa0hOKu1BDJ68G4Je3+AESLRWfT8Td
S46sv36V91waAxjE97v2WwK65ESIEttiTwfyC8megbO3szQ+S5Q7sJXXzyClJ3Jf9NABnNZuQIfq
lIHiRzXQvE0JnnxYsYjsolP7IwBd1mFkXdDfusiFicybnwCRqvvn5mvuD+eeoPyDBIQOIqzAkU3s
rHhGcLi0i3ce02+1nQCDfXI2sDzsZCtEVGxklpraCtXDD4aMxld1zW8nFh9Fh8eawZuk7qWTthhV
72fPd2/PWTZ06qyaEmjPsYynsYSM2VLbZXV6C9NgJANgjZi39S4TuNDuIN+xZ0G5bVg2Fqikdj3r
NRuIZvJOQyiTqdD+cGx7SSnyLsGPO8u2CirwRWBnuLj/DwQienjpi707ijAQLJDq7Cd8jD9KfAL4
haVvRXrTQ2zKA9DC6ZY65W1loTLqu5F5P0BlcNzU9TJhxLuV0aQu7ps2l/OYjNT1xw3ST5yVfrIF
Y1mi/30Ubaaj94vI5BNs9EtvhkEsBk3ogZSO1vKEEnFxxZouuWZ8Am87OWz1D68AIE1cQg9a96s4
idbGc7IgIWTDLXqyaFobHgZUL4wjFjLhqJJtYKsTY+1CoLCeXJBEfqEniRFgFafWQNGHOm9gsZj/
AH4BuLPBQ3gI5XvztXiDbcUVg8ryvWZTslvZ4T8eylmsvUZuy/PH3WbLNEc9V0m8jJqooCDLmMnf
1CSCgPCEfPYfpA2G+RwThNfauXcNhKiqlOw2dqs42M1rfDJxZOYejkDf3r85IG2Px+ICQMomx7CO
bURY3ixYtdbkd5spqIFa4OSD/8W4ey65GjTPW8gX3QdA+qzbrZ7dfD/4XHzNJUV4qHz7gwZlplvF
wXMVD3Ot/vYZIdfMGB/M8FtIQU7qutR0W6m0LD5tY9mSYlYyNDJky7iXo4pmWbWfiZMgKPFAwxKa
Fdbb3OFZ3aSywRI6hlrQ4cPLt5B49AM0drxwdgtCm72yqlhFTLTp4j9rdbIqxj8AjEDKuvHhHU1V
d4yhPkEwIQXGsiV/vC8fCIvA9hvl6dkgZVjVI8RokVyOLv63mEzXmWDmOLYS/WPuQRrqZeL9veGK
RPg57s/eSiz7FgwVObpRRs9ovJ4tNxb1B5gKr8hTvTf2aWge5dFtePuT3j3obTzTm/YLS+GGcmpx
NYvtQXodtBAqXTFWHc+Iw4DpbHforzASFVr2r04xNEonoRUVcQUIMAI1BanlySV99uJW8E7XHjRh
9aStKinPdlFBiB4bSQ923OqK/PaZJMCUr1hewpkx5YXM97Dz+ODbyByDxYJmuMXnin4qjWAeG1Uc
RwML0OtEAbcmmmUwhf5hHlMadqxzoSqBuq9p0FffyfHPCkxzeS2vPE4Lk00swN6gmNrKbLkmFFTG
ssPISkhEkmLSLukCEOfxZVZm+q43KCUxFMrDzbObf0NdkU/NenS8bAcCo4uOWIey+79Gf3vyf+Xw
CtOrPem08VWEymjC8UIVhFQXiGYdBykDpBWZvCt4qflKsyFZS/S2TRxreXoTvnueQJfaxW0SJ1by
bVZb6CvT4/uYMtBrYV9FdHXsBZodkZOK5L2pp3Vl3rOKz8dCLzqC0Bg9d/5AKlLpiixp4Txh8eaI
rnsUX0DBp7CRNy5DyGVNueSH2B2zPF+/5FvRJgnF13gheSDizPdCIi6r/ef9cVjy2bracxwGEGcu
6mMqZ9opwQ+VqPnscov/OV0rvrC8im+LyjjFCqeY3J4FyhMplD7pjHo3ZDnCfvgOQrU8cbGi8HbK
d7Z7nxHvAVLGlU1GbTgIeZyBXobxgyk7bcBm8aodDPq9AGzH/VqnzdUrmYECprfYwP6ZorerH5e+
4Wo7ypdZ2Z+rP+FZ+oZ3NtC7d1h0Bki0loAenjHAhem+fRtR3VswxsfTvv2twxCof1H7tFwUmwWy
C6tXz5J8neF2AWHS2/3li1rHHQVTlz51faMplkMr96HRhYG5ceBnSv69Tp7Ggo27qeqYA5b1CTvQ
LcWUt4TpYlVyJ+A+H84FYJPmVsljCqPAAZKKY0jdfk41k5SrQJH24Fcwnq7BQKdBusaASwGZtSFz
FwpeFr8QwhVgNnLTOWwJ+3E4/ou/5PqJo+Libdx/ZwEPE0OOQ9u0hC2DOb1WMVytX3IPMJX6WEU3
NFY0oIyIEdxnsLq33vnnGSW/54v4eoPJ3sajkoOCjQXnFe0HarWbRun27SCn71CkuGag1GqXN3mg
m4M8mWA3IPRDF03iB0dieYdzEKlXsNii98tbReMxX6UIZOhBTNfdhA8PzUpTNEd2KqM1Xq3q8Vvp
11foVqMirSohCl0OWV7pze/2YWmOkLEvE0Ti3IHNrs/31F9ffUaB8kfqqYcyVc5Cavum2VuryHmn
vtsvWbnM8T+S8+XAmrx/7MjX6LZLmZqUu+P+w114Clt3oXy6ZgIRbMpvIMB2quCGBmiPrYjr9PSl
nIuxY06HtOBCZQSUVhWjyBIUaQ02+cwE9z4YcNGJyhlX9mtMwe8JswpFJLI8Hao9FdCp7n7r2tij
YJS8fIB5VduBHzUt/e1duK/lq3MEhR1natjlyzy+UxMLcPQNurP1GGWzJvIv6efPhcwb3eyVIYwO
BGYHTB8OEVeUO3qwQLS6LIKf1ETqZQYUr2M8V3/K2sgsjLKFnNNCNdHQ8UDnfxuC4cNyjoTHl3rG
IHxt2083izgR/1yyRsQbX26lFAfLR+v0j2tA4O7PpyjeSW38kVUM3U7UborsieCjdrEt4Bhn33wq
fJQAcYffU/fWynTrc1X6TKEVmeCccpSD+ZTeGGbcoAWS9jzLMCCQKZ2fY2jQ97dC6KXAA9cTIWWs
5dOQVlO1ucFJdybG4ojjG3GBKWCD2BO39OROtqCmLVWA+D9f57NCCretPZS6bZipkJOIuJO2oN16
xo8P4y6hVUknIkKoupF+H3SHA8KSLBi5uVF32XJj03eQICYE5bjqLHSlXyUWjO7Ot4aYmAQFcP2d
OW3b8KLNJWst6EGwqxN4v/ulyIZcGV3tcV3KRP78YMNSUzhIaem0GHmkAzUCXy5CxF63AVBcmUsD
dp5VBDpUdhoRlTepOygghgFyPxnn9XlFZreCM3R0ZSwUDTTInJgJwWx7ibg7iYqJi73ysZ/zJMSE
mnOVUhBeRX7pI+2eDPFaHKSqVgntro9ErFN138GImU0xcQNvnZk6/f5wZMSvwQh8EEVpZRpnVyl7
pYgYZjbEcMIPmOvwgmEscxX5X8cvV3z8aNO7B/i8mSvrmkBFjLX5XPeJDmdIFBlICez3KPYM9a8v
myjNzuAbm5kVITYvCk5/SksE0XYg2tAUM4OIciZuD7T0mJ1eW+zxpBw73PKRKBdOssHCx5nCddQI
NrVm1D+L2RfYDKL4ACf966R7kgH36GozyOQmLQC+j+9LZ/0DdEKSCCi7jKOJebx8LM72y+PzRwTA
ahbU5NzkbT4mUG+H94dOkzYvtRFd/NKky5nnB/Wu/VxFT8D1ih3UYg2ihIcehjeYULb42uVx+KKL
XMFCNzDtChqC7lTDAtjg0LfCeoUsaz6ZHvCQ5SobU1FQe1pTAAEvzi4AUmrkLvaEIqQges7i6VBC
6vjl1T6L4Enms5yUlC9re+5oyHhXRXaAB5lJN/gWaE+LbbkbH+BN34Uui+9HBtgSYIjRUaUy/bU2
sWSdwiMHdOxs6El75+nTOsrEfx+mskVnqUL3VQUdysDyOUDBymlcHMpiN/tJ768teN2jmRBdg0OA
x4LDap5GV1a3/h7rHM5+cp7rJ2zjlByVgCsNfUoT8AiYrmciwr1c71PM9Gs53KzdaZhgfOg1RhXb
FrXIHwOH0HETgEsX5MNuZYkogAJFthoqP7Qtj+/GYk/TY3dSdkFKVYScL4o5JyUbek8WNOEEcuxU
F/C84jLGakIIgLHMdwHQ/A+yqKtNYiePCSYSUCLPPm4sVnKhI37dktyuIpFBy4JMclzqUgMJqtOc
8HPZ3/+K9QpPCr86bMEAQBfc7nq2W78oyxhLeHdlUj34mmJAeUH6E/NtNM3XI7I43mkvylgJ90zk
OPCWdxbRUxZ7Apdf2/NJHVE5HKLdN7cgPaAw/Y6H1E87iZBsi+3MgsakiwGluCYKSDZq2sRBbqC1
ocAKoNWPcbGI2eqQ/uIBcqizQrONMHJXB/EUxyNzuLNJOagDzvkz2EqpQLqg9FnvSMcoOpTAc6nr
u8+chyB1MrBMZWWrjX3qOKBWvMcNLP4MtGhiIVFKWOLyMGn+ZDZRS2XJWxxdjcRV+Gpq+3FtnnPm
st6F3qXlyJqHsH6Z56k07Tq31hdf5jCN0Tb5DKPpQNgKNY+jDDY1MEZ4v5VjIy/k9FoY5gVAcZMt
lVghNRVsK/VRpq8i2NtwKvN0vOo+QVDX85VcadhaJaAWneC60PilOxD93XKOt0pEsareIYrKyzy+
fC4DVxXx7Y7e5ywabYNd23yecwEp75nm7Rou+fX4K7Wb1BLptLsaQs6aoV9iumWnK39yKeVQ2sE8
ilnC2opjWaEF92fKQqPgyoLin4npzups2+/ynp0r+s2hjDVWFFKQPLqZg0zl7yCHzcK4N88Ec9Hf
YYe0HLfnDuiE/qUfQuGfJlIesMYlb8/nKT9loN8T4iSB0Cs5o4PcLdKByQcKBgOJRKGETYDF2KWM
ogCn8wQKNeu1S+Cjlhkigx7xuVd7kSdzgJScAJyjAMo86qC8c771q0b1IX2D3gQ1EhWhAVImKiSj
NEmPXGsRnUsn/nX+Vcfc6Nwzm+cLtG5jnAYqYM8zUbxwu3EmKnH69EfJxQHD6xYMUO1/u5CH1lRp
2++t9iAhPCVDkMKQRgnP4nNO7Eou60U4DTB41slpXGrMksi7Jzawbmx52oDkbnVsDqirj/ALmOP5
sbXK0XphNVW1JFmACgr3ByHQiSCsqaWRK6Nu8wBRCcQmJjX8FPc4may53ixlmkY2rOvH+IZ+5t0c
gLcoI2kDZKX0nlqEhjy8X39e6+wiwRtEAfc8OPKIqZeuWved4EKMouccEHCwKod2puJQ/9pyOG3K
2zvoet4wlwZDRvSshn5pfM+yXUIW1NUdd5zxqAd8etMBa57hCQgbuwIMrhs5Rs/fgHw20lQ+ka4V
uY5tsfw6vEaP9U1MGobKPBBMiykeM1fzZlKNH0DUBkMAHalDEWnuUUnN0PVPcmMSGATJPirTtv2d
Z3FX/Zvq8LHJp8rkHyq57JVI7obrHDKZ38yIWGiSpE0eUWv5MECFX5vU2Q6xRyFEu185xnH9RvgB
3vekAbaqRkMLrvnPJ6PH/5Cr6msZPnCiCDNGeYyXT3uwcbve4by6f/j0buoLyfToq7izBGXZwyGQ
f3DapU75Wj0KY52osC09G6u6kts4SEK+BI1GOn3hfAx2KI/tUlwTFL2U6UVYQ+DDFQBcR6dzwbrD
/Hv/ALnEwGPECJdRDsShD2nuoHHAn3d9CFsltl4ozCjfVLrDVqZUr2Igi2zmQpLzS5I/FefexIlf
yFtobDtOSaEo72RkG1cNQS1vIBJmDduRCTkFNp6JepbSq70ZOWFsW0x9KBdiIh/+FGjoGxjaf+UM
jZvUnKnzr7bj0zXU/fNE7SW7ZXvyfZvMiCh0M4Kro732CpAP5LYXgneSMhvQvU3I8QZk1u4Zk+Mn
KgGx3vu38LIXPpgV9lhLZfCossJncavLSlNxEA99ihAxTiFuljtDC1z814N0SfSeQSywjxd+yuvD
19ML0IwIdMEfgXfksUJgcC7/e59XdYo27FaZa/vbfURBE8iWJdXaGCid79yQ3KaVO4hixDWcglDX
wGBjeGsfW0zuQxbbYal9japYauY6I9Yn5/JUJFfDlJq0+khpT8U+rcBuarJ5xFnG+PiUR8EuCE0G
+XSH0IrnN/I8T0cofJne22npMqGK1DTL/GBIqn/FySpGYaxkxknQwHG86hF2HkpJJIE7WzFfStZQ
H5ib0nbOK7FqnU1UbizjbG8A03Kn12DJOfBm6/j4bUEFKxtIWeYbFCG0oXA6joRiQBPcroX9AA1k
cxskCYA+YQHovMxtnOXaBziacsgTWSkpP1Px2wFuyOpJ9YHSJnHR+6yw4VM0THupDNf9elQEbdTq
yxwda7CIhEVIviP5R8uH9kn67O+o0ydcBLOTzQyL6UiA9BlpBEEszvf9gShNRspTCGNp4gE04pCf
zGK7o740urHkucS4Hm8Xaj4ECUZBDfPGOUvkl851RDAjVKhuzmVzf+Zu1EiVPvVidphJZGMaiatw
l99FKEsIf8t7NgOEuMH3LJltqAHO4ZfKE7+3lg6RuiEx/PkuESrx7fzcnWhKSkDbRskwkundxZ4d
i9kN8aL0+fdy8Wb++nXIxJYCr3V/DLBkCS6YmrlutLweXN5G8sd8D2cV4kFNKR5uNrBuMRsf511p
EFwqED4ublNRf2RRgRtEg9Tpw0U3O+7KxxwdFyrJelbYIdg/BB0tAARQtMs7RzIb5zoSsozMhu/0
Fmv0l5AXDiQrMLf1peEH2cGsfn014+foxvEvpDuAQEY08lSjW9SCuZCKvHwbtd7ulsV+HTHgS6Hu
xcv4xURLpaZHJ938ddDZOIgKK5SkWfOA3oIwC0IMM8dLaX2vv/b620B1uzYHtx939BbmwiXNWhDe
dmCxCmBbpcMU/iJkYmXgr1k4ksDfMuPBQKVIWlvmhrwn6ljBfNJ5GXGDABDrsRUmv1N9Yy9/Nqc5
Zi620/ksAHeSx23/T79N3X5QsBQ76g1DplqfzoEPqRtG7NPnpUyK20N3v5eEEZYWoqYo4TLxrLJ/
7pI9MlygEAsJFvqs3W9HKbS8q+6ZAwKQ5iG++jzylyDekCZ5G0lbQaxX0ZYWQROF0b4AeMA22WXt
9L64GHUJYVqDxXrWhSULGi9cpf1UwLYdZXJl1l7dtBbSAU0r4Ajs3ZQlnfAbZLLbu+RiodRqIMyW
9aTmEJCsrMbutt4CFdf//QtTeJ1+VEymtLdkLNBOF8DXRYw5sCa+snkgRka1SgxXPu5kSBHYec2S
qrdvcwCC0h7bczsCPrVI82cr7noUqceAUhdHbWjSoS77f19enFtxo3jIBIdoMcHlomT6E1/l2jpK
MKKNGUfzN7vHzhx/PUZopf+bxEO5WQXQG3gbUXwe3YjFRGN9eEk7+dENgqeHyuk0PRHZkfY6QWKV
SUDxs+H419s9MjhMPau2IahU7gEZZkA8clKi5CcSikZ3nnRmENWJYjaAym5Lt1CCsH5SXOZGkzxD
xVA1n7rH2mx6n0LyiMMzzMvg01LscNY3nHZaiKcMC3dYgwX2DrufZH/suyNITIPf3pa/L2vtiek7
ay7SOdeGk9f+2fg2+iGTXZV5s3g1d8e4mArEEK3tptYCZMz2FhnvwK3daYCUNxLQgkNGJA5maeu7
l1KSh7pLB36z+Mnm8dIy/iIfDFXwaiMSv7zfkPUiNsqK9lpoeE9hhTIusBtB9QNzwgB7Aob24hJI
o89xwkPycvrwG5DZhGxMDdBSIhpY1Biwzl4z4vkdrGR0+gtMVTHB+z1238ThhdI+E1M7MJrmM6Yw
Cu6uS/rGPvtVkBDaB5Nn1/OxBJcoluGKrW7MnUAbbUidGLVJG0Kg6sxe2nVFIENr1qci2k5O1oTQ
ui6ZBOdCkILOfwufn2EfObbtMYTkqFsj3miny1zm6N59yNSp3ExcmSYepG/Nj8LQUzf6RYnqfQX9
CQYQCmeP+lPYgP8yuJptbtDqrCMpuah3+EMql+5mBLTnppWDzx19fETRcdtRdpq246pG5L2MjCRo
KAAQxWbV3f7O3F5zj5X8CrK9WG72hawW40RmhpCUEgF/S/m0wcNVKKCA9spKGgCTaxru5oZrj3QF
MDpLaN/mVWhGuUDXWAZ/ak5dW8QWYD7/HFYNfjV2g8YLNQmjK9kn5LlXNeCZc5h4whcFDTryz+6M
CclcsbNxK2OMc7RQGMCwtl04zFun0bPoKjmrz7iJULCGvhopqEyLBdC6ti/higPZ9hteFVjKmVLq
vDEwXE5ejIZ3Ig/0QjbFm3E8VRCTfr/fdbmWbnbWovVcpEjeoMjFbGNq1paX+s6I6PCSwOGetZMb
biyUmIFvkudGBksIlT9dLGLUA2REsTyWaS4s1ZdfUoQRNr7XJ2h7J31f0ohGKkeAhhOJfw4AVU0C
Y2qxzeB/5aaYSOovoq5/vKGiGJH3S/+L2rZR+15XosieZVmX+sj2mvk860RNBodjKbHcveiquiAY
IImu2QwSjwCivi88vpOxkGIz56nDqVd9CdE+Igu0N29nzIOim/a2T2Zz2p1KHRQa9Uz6RirQfgQo
x7G25fbRncgWxxd83vosM6x/vyhDP7BfoV7JSmRrFAtVewYLvVRFxFkpocbRT14kZSqZbhRuz9Hc
xIf5tJgM/bGXRQ+kLCGmN0UGXSvNQyff/AkA3fnwgMhvGS49jGDuvkvjn+qZNNbYRn0KfnsUK/hK
G7r+F5BCaZl+ti3XGRd1s0pOz5TJbWG/+xBBace19PTdivfjxfcR2xpeK8pcIsR6CelYRxG/gkju
LfNZann7AJfbf57aXBUtoiZOAHfjrxDRybY/7SiXV3+n+h+a8xGVCNlErZ5eAAzT6GZnDCMjamSW
i8uHuV1L16Iq65eyYhdEa3CdMdXpjf2/ghyePUFai/RQ8yHQE2im//Qzua5440EfkZN2rMzCEI/A
ul3bK4tT/+VorloUYnGXtFX2bq8rhP84Wjp15kMoGz5EFfQIMQebuB8ebG91f8Ettl5tQil/+Zzz
pZPMaFl1o05xGeYXheYQ4zmHExUqna6p/6Fu/ilG+oHboE6r33in7q0RvVBNjPaPssnqWsYQQ2Us
4z+PclYq63NHJJMdbFQY6YdBdi0fZAbHMRuPYJIhkpoii2+zjNVw7ACcOaQpzmFcM1V+wWnXA+Am
bsVGyfu88DPVzTP55ES3s0lJtnZ2YB7mJDwEu4B6xtedLKTi7OYcvYH4aZcMeczERVgft+l0tNUH
81Eh4iIFq3mZ2SAp4K6yVhmK8AX/56Z72lxnrU8t1YyDiNR4QrIo4nhQlRLncawyE9+nJaRwNdvS
PpBoSLwon+ZM6ZjWShzFyManRADS9laR0wkKDkUgh48fN1b0OP+Pcl3B5d/izFQp2CGggw9dZfV2
xwz8WjlrEf5pJemzSm84Vn4FLG3TL/0y4k2OFFbqMebA+87t7UC4eEofLyWS+fsQHnkPmbqZB728
KtT0uANq6a150+XoiRSBTV6uCgKO8KHLtUrTzOsCtHzJDTJBueTWd470ncyDYWjJrTlOL+AH+/Yu
gvE4Ruey3PepFzXtek0BJQh6BhxI+IA7n4SSeeT2mCUwaynQdOitU79sGn0RZ9hCXDYzPRSr5981
u91N5wKSRMlHHrfPc4sNQTaZUUPoV6A4WdVrAi+R+mYvczKbRd9I3m7RdJefJVYrEZ4tEsmu81JL
IEKuhlnsqrvswD/KRg4Xuhg+CUteT4dmE4EnZh0yypBYuvVCk6I0vIR0A80qqjqnv8TYQYvt7MmE
Ua1e5hHGM1b1VerNT/KqXf3q/WCnqX3iZebkBCTEGM29KicuqQmDDwtQhkNX/vZ69mSjLgnQfQuH
I9EFJWyfxXBmppt5rEpjx1aOmPVtTierK1bNBHd5fpqgmMQYFgihPeS9TAC1G71/WVWHuI5bdKXq
9dbdjeBfamVLpkbJTEIVL0uqyXlU0Erxk96euikmipmPQlqptM6Xmw/UAPcGV49hpTEDDWz1fa7O
OHXXup6z3sMFQlOKORuztEtIixFcIk/r6mqyWsvJhZBPXsGfGVJjZNEXvvnWAbvbEA0M9xe464y5
t2gdPFq0C1eLSptmTNmz0gB+JtFBMe3TjBpnoWIai7fBDhEUdhe7gJvIVcLbxFEqX8W5Euevxo9u
RY6Ppfnp2TjRDrg9uvzbBv2FRXAh8isEjXdceYTJr25AFHZmip6I/tbZFwDcDAXLfA/b9550nbzZ
4u+vGgsVn6A8hP5kC6ldE8HwGgVIzMWZaFiC0uXqxG7SMFhO/e0xdiISBtdnk2AToHimJK+Uk25e
qesSOZ1rx3KXkPSKrF/pQsAbAzQ3uas506Ne/RoHKGGEwTgMZ9FQGJDHxUW+iyvbXuG1NqX4zOKf
+1vFaH3OUwEg0NbMKJGJHzFcpp+P0rq84+86RX9NEUyULoWQhWJ1+sFVDoOSTtZOtAAMuT3rRKMF
RYlsL51ZNLOiOLIp2hX271Sxfk40xm3W/miD+OZLXtgm2r6s/0tSwjbNUhB6xse0T/kwssBiN45n
thNWN6Kz/s0yTfi0hcoFdizBqND/qygRKaIg3Ph5hdGXUn5X70qPH0xx1lZmCdcigsL/+0mB7Fzz
cKq1U/g5eQ6Y7ejTS/m22eiuaJDTPMOu8zAfKL1h7MiRzHc3WmSsO1WHRQjH9dWwatBg2Rc2gEmA
d++TFGA3aTVVwWNcgp/o89ebNs7oYpCSe0bOMGrYiuthlOS0ge2gs0HURxpWPT1kmqE1z/Kmzafg
3u4TUeQbXPNjJbfjxK2k9qgIScTIbHi7YSvJAaodWjzuVOL47YK4uA8zqXd3hR8y9U84OU0+enBS
5KqoMNt/1JwjYTKbPWXm6J72KvgPBuieg+LkRp5R8PR5UG7YvlPn+yzGxATFatjojxdbyx9U0p1p
yV1XgNyrMtPU3HtMcZwJ7rgQJ3no4zfcVk/zqCm8bt5pg14vdws+mmDQdRx9YWXlqlz5U895clBJ
AZgwzjiNb3clVf4ohDtKlL1Vk5sh70VaLhwF7mxUu8XIlkHjW1rupbfXuxueGNzF6tdFovfMWeVa
pO+UTFljHVOThxFuO1W0mmQEk27MF5k8GxS+/ed6+kMA5TRhfDEGP4P1ixrcO7Ebn7dEmHnadAtZ
tGqfKxkKTvxx/rylxzQplsn4E8CSOEMttMby83WxMm1t+IR6J992M5GOAW573sWsxN7wUxXLSI9T
J0pKQ9D54TJzvnkG5HwfdYD/X+xEAjZo6IIbKHpP9U7BdfMURzP+oJ071axHUXo7PReB56X4jC1J
7YPMYvT5kMokddSeggdIi0i7VwhIfYIr3tBDoH1o3jNifUHEGsTCEJOmHCkM8G3rNM7dGpK7rrD2
mnkG+Al5755qVRpP/8Xcn6WwPuO+SzPpG7C5KlJ6PMWQ3qJPok+9xcvqEeIoW/34ettEW532mnpZ
LT2r6o0ZSyPa5TiPh+TqdSzZACv8FgjSmt8zH9GhePY4tSpUiAfPY2fZs+Woq5uwKfdL/bepfP5y
dyZqT3l+hZiXzDvA/SlnuYHAXKxXryTIN4iU0GqEhlVnH0EKMb2pMDpak4IpVievNreIr0/lXDkw
lxxr0w7HT4J9CIr8exRBMSIab5WK/IhTum8b1Oel4UAgXVF148p7NcmpCu5dzJcHt1RMEB0vEUWg
T9dEUyaQ327Ukup8lJORWTh7pKMTt7txFdlJfBuUpQrIzVLVxwoY/c5KG8RRIJyHW43XIc9CcMR1
zAINgAqB7ASj6PlHJ1FYcDv7LYem16BZAuCv/3LwQ095knRoWPHUTxpkXLXtftm/q19V+5gyjLTL
CZICMjvXaV63KfzlkCaReQIiIHbh2LiLQO2aIluGUXpiv+DwtFwHG0qPIDiarKy+QRG7Zzs+AI0q
+OzusOK6NyN5Zzl7C61X39o+iAWgzP7mTSPmpZ4ELuDJoOk/uqlEShtp4hcwa/R+4rY81+gJjCqs
OMGOpxKd38TbE+Y/rw+746yD7AaHx8TAbH4nQSv+QkfpqE7O9UN5+v5RSaXTY603Troh9xZkdVZL
9qUyeNFkdcRnDAyI20ffUMS1+yiosfYE3ryIKBIAxKiiDE7P6Qkd3ocpLOP813xqnqfrA3yKHN1t
RuxMsb61pqSmVfzRnHABtTW9XKMCOW+tqlrPQMM6ofwQ/TbBgRF0S7IbTKhwduAn6PE4E80J99Ii
9cpcXXhZ4OiWXAEWrSNt4NH4Pfjan3MUq7I+dzwnVsuFi0paKWjb1LkXSn+4WuBlzq2LbywCA/CN
0vh+l6ywwKnIpN2FqFD+sjf0ZjjxHuLJzVw0UV1RhCQd2Qv8axl+ohOR8d5zAMq4TJ+lfpDe9KSY
pblIQcQClp7PM80UeAGQLAOl1tUyQ0L5jpYkYwPpfoAQBLQA1TzNhxd8rFX8dE6sLAmySOxYVC4+
c2NfjiX5B1R3hKhwyhv6jPmJbACoo2zBKelTUy0kYsJCCo7rLXSiucfIOUhXXKZYsDVQvbDjuIsQ
lhi/zlaaqM5aroPJzrXER5ij0eaOT1jL+Ub+Vvo0wi6NbbjNgOMmb3OBx+QuNtFLZ5HPPU8o7HDi
u0zIxv0f55YvsqPXK62OPqY/CKt5SSmoIk0jIA0JUl6bimBYIHLya48nnDDjlWcdHY+Tm8gruBpG
8hmOi6N39uguipqpf2r0EewRxYWJeYd/XEd3YD9sEcfp+jaOyCdXWcDgHDPSIdZ/jz4cJWdRC9V5
lsWdlU63nRHruXl698J99kHjXUyHbU2G13/+2ZOBXVboNH83fr4+Og3FRt53Yb2d6kHr2JTaLTbu
WCNmUL3OeAcdVFSyUvCFKGtebrm6SkHZ14mtI+i6uyHXPwl3hm5TsgYvA0tbtGYwSPW/X4/KMcYi
igKE0EJbRnzeHrzT0IJpFttXbjcF7YcPinCB0jOOicDzf4fN8YtyAolue0Upgf1do3dOdHsMmWW+
g+vfzlwbkwawasDbz5bNI2P2spHUCxX9xyo2ZrwVNHQ4z4TNewzGy2yCHNfVVTXopMQxK99am59p
bEvsiNM57w8uDgbcAcNmZcUFDCTec2oUyxtzMQSOW5Ora9KEB63R3iqAyZczxDlqEFidpP8X3Y7D
l3p4VP7nfmGh3vPB+dW8vHujmQs/yO+hdhKsUPpZT3QHTPzUgxwaXo/oG3mzXLgju9jTPAz7oMVw
qAXzcjF4e7Q9REY6QSrCxeYE4DgHMmRTTL2y6EqTPdsYSDK/R0l/0CNlGazgB183jhnKedPZWPzC
K/cRMciop10MzhBYPfU5SaEmk2QTfCq5eOGVC/W7JNaNQ3lNqM5ASGcd6d6VwznD+UesTycL+4XX
aVL7+rBadm+ddNtrD1GQLIGhKXRn8ViAuei45/56yebC7mq4whSbCp9wsv7JNkRKbmhnsHojYQWJ
dvY62WRKJbtny9Byp/IDa662COBmk06QQvhgBBPzvWS7Gs+FxjCWvUkJCGIs5GxoQcHS3mOn7sRj
UMyokOo7/ZzoC+4MR2EO0r68z+nyhKFvRHbVv+pT/FZeDS9hPZ+aidKfaeets6E3MSAR2fO3jugU
lKSlHXCAsnOf4z54cxjqpECvl2h+TM0TxKJq/6pKjNFlXB/Cr5O7lpRjKTY5Z4oaZhxmr0EOIfiP
ZHA1fd3l4Ui8IknK9qj/XCfUHnj/OyIqo29cX4CXhfzJnBP7UzgGeLQa0uk+LSxB9GF3XJIziQfZ
GUtu6mfiv0WJKRKtPjY1VlZ+SP4t2gLFFpgo+Lf8Q5JOg2aRdsH2GjjmiNEZhsTd5HpHhcEhqJsN
Xut1CSr3ekT7pE7OSjexbApkWack8SpTI8AdO2sV4VNgyhRXoePRIywPc0NiYnkZUsDN31/NYnJc
fgMJQsqV/e+sBwjxswRCUn2qiDN+tvpNCWRrHGqibNQekTGi7A6OKFtJFb3qmlzR1W2ddNy+aQbC
86IZpAkT57+DycUzfYRD9IRXeSjwfefA9mTjuXqGti0lYXCJgGGRbhhGwuD1mSt07oMppgIk6Ta/
FA549+Pg8lNRwzqjE9AgA8tx6wl3gHBx7CmcSs8rPRMHic1RMYgMFAnQKcI1VPEKN/JE7ID1XnMJ
JDUcl+mXpvamF0d11dWswCOsa1qW4dYqWqW3ThDCubvKOhZvGvQ35c8B3XRVTZFPM6A8cjceX4IJ
I80+BAgmwR5Z/jKBdjn+DhvlZm4fzbeojIuDirr5EgQ7jcuNPiMA8C55kal6N8XD6lac7zsOnDEi
S2qz32ldyfZrQNZZJu/GuOz1vvQDl2xfyL0v4FNKU/BCV+UwmAmhitCrp5b+7W4FHBd1NeC33t/F
IcksOrKcV15HqeYKxtqhgk6eRZj8ahpmdTqx53aQCn/vFTWmeYfpMeSMSq8d7bMphPSkpp/rnd2T
cyaGi19//mkKzpTq7BpOs0MvCDTFUPF5ZLS0TRqGDPYAAt0mRhnR7MRSqgj2/24ea153WDASZ5GA
qBQPcl9fLIRxKzXCpz466guoCnI96+XE3PboRqSzumeBAj3xdvnT7u9FLLwmAfcOo33KfEPo0kqa
D8m3HEo8SOEKEmoXyBcfvcJlgcQeLXcheN+qDllgS/Cg7p04Uq72Ht+AnebzJWr1UN58X2uolKQM
kte2XfhxKiyyFJvMmz+8CMuZbnl39fggYzS2S2/0H/yAtnZOMk7fB45tDH+Xyci1rN3zSly6WZpc
McQDiIXW//9EYFqeY+PY8BDCeM/vQo2o+NMJIT5qsu3smcUcrApxXa+R4SrYjjhygm5j7f9Zilq/
z85mai0QEwUauegarXL9aNk2rwMayb8DSdWyvLJ6TJ1BmPkZTPuP9ifO5XtHrXF6fxJghAxPSt0b
FlBeBBmOXgHZA6flfQ7wDZcXcuTm0dE4FACpUbLbCeg2U772m5OGJMAdrx5b3iGfvt94WMJH6s+n
BhA9YBLWmKc41s/iqtqojcSIaKY1EvULRMLpsf3cB24YKw9DTY27ho7Ce9piu2bbmxleOTJCdfOP
dbFCfzIvPx4m9p+iMgRgKvDsqMENY0EVuDx24lmlpKtuVCT4T+65jhTiPyuEZ9LiSwyjtR/bNuZj
sTxWShbWAbUbenvkhZit0Z//M5MqIP/df6P5E3z8dJxWiXAL9wXXKaK7MAWwMEf7gzaKkyypOJsh
8Ykx2NHUog6U9drfnQcJh879z1WJWXBacQzVl53MO2UOiWG9APObZe47sq279XQSFBiMjZUOKE6X
TNQJFjrTrBCeIj7aGgKwu4rchi0WH7iCVQA0BiH3cOn8Surdmdt7BkidgJ5xlfBvPcaITQOp0omJ
pKccs9A7sd1Sa141Y+5Ovu1IoxHcZu2hdTcy/ShmwjkyRdOyJbcwTFxHTh0zPHZZwvhLwttvPN1p
1tlKuAYPPp+Lka3h6hRL8qfZHYMy+qq3pbVKBDdf6fUQcKgJcFsMkE9pCAsT9CH4oYzByqLyIysw
ExGMZqlImUAXbVbgGcNYRldwd11TqyTZb/V8ofjySE3Nx/obiYUvsO61MHF9PgPjk+qELIDxOjwH
4NBjmHPqecKPr50VMd/lS2hn855D1TDNXxUBQjqNrlW3cGjZTAQS0bjto4EXUaioWyMsWK6YEaWe
PhlSrcV1UHN6ZOHdQpcxLPla4xfMHyGpRGbHEcgVuO2eLjbf5k4xrJxfeNAUQvRMwuvlMNrStMCN
zO+26uWLfEPlGG4Vo0jahcSLvev09oy2q9YHjd72aI7FBb3HwlOR/88qpLpiRZneDhafSLHh2ERS
uY1Or4DhC5gj02NP2D7N/rBmSDUmPYL/golObAbwm1YrIQDrQYKLpMLP9o1ilXmyM2JASO3iVv4b
I7F74SKc+BixbiRWyDSX6pAmixPrqtwFp21oZMfTFITN5Zxq7a8hUgatk8iYJn4kzC+k9TV2v+M5
dvkpdR4QcT6hxVNzzDhavd4pRngBmzkq6pCMcXmXeKQzdMiJIR1ItsEfIkSkhxRJvHoczCeJXi1Z
xIOqkPWv0dxGZx2x5c/8tzVphyhv590RkGWBDEuotAb3hvPFXB3pULmMMbdViqbmcnK9eMoCMHcs
FSvDiO41ur/RwtcX8qGZl/rjwL+twGj8uU++SrrRuRKesjhXD8nI8Cb14rFih4XhiAEMoNpDpAtd
yE7+ZQBbKfj3xMG9+5L7Ecc7I2cozxOtooWlE+3+wrXLCckMURz2G7rWIbomsNi3qY4bPHpgYJG7
GPsIVmup3Ck/MaKyMsCSXwleM7nB2hxOoZRkWgw2MjMJ0WaroCwqkSmtDd6jSQ1BUvBTdB5Ispga
dm+4SG1l2Ehd7COHnHqiS0PVRee2JW67OVckHzXrfxTaCLLlWxh/1JYPppLJa6pnHPbji5WOz1xa
P0belF+mY4Ypkr3wDCRvumsCdqeD0FbX3iC5A9OCy+jkYBpZ1VBtx6JMPdNAWiLyPuEGnKJW/W91
lnrrro9lRRbAoOB0rSRjbLXAdAGiDsoW4qogWd2uDLqhgdx8ZSuiTbE8Ir/maGIcP/ZwJ/9xQk3r
abMyo4qKPhXVk7fNcUGnY6BBass+T1Oe98HEYFjdv6D4HKlzsG68eUcW5zCZ6Y3syIE4LQ+RuXEc
0fwJcVIsK9IIEAc0JzptQgPtrElyyH9JdnaKbji6VAu67k52zWZeuZi2MVRdEEdH7DmopNcJA23N
P0zVdjIaJ/uybBFYjvBOKrvMVvIX+dEAXagzOZ/BhPS1PQF71Sx894UTONVaA9DzLpZbKq3gQdJ6
+uYLokTO7KAQKG+pOrbGjAw667KLs4geXVwqJhQmUNXIWFpHn1/aShzUxVnlOAskiNYGc6ipaxJ2
6/KultGJfDgQm/Z7j7E/JuxAyZZARa8//IW1RN4m15whMAfGp9rmIcD5BNDTm5OhEvv/slE+uEz/
2fQ/v1m6q180VTOfunN1hjA8A4YeNlXK3hvcKGe3Je2CTzes9GVxzCElyPzOoOW8Go+ELOS3Noqg
mIWmrt9lbDogz9oYh+CdFBTduVZgqfRcr0Z8jAusWLRJjTdyhv97+gGmXWQuUkC3l13ehQIiRU1T
JQhkXQ7tGfqAFzukDS4uWJuF3nlNL1Cfk/wUs6KY5hEx1oYVRXKsL+OXdSLlFaDnX6qnFt5v1G5x
ZmYHzaTbgT2Z/Wxw2GUI7tOi98csQDrLa3wHXS2cqtxw068oWSopfGSmax9imOi/KDeHXNw6SE+N
+WKo1EegW+vVCsPgWQMwFkr+H3HixQTPOnpwNbMNecjHO1KRpTXdx3t4dXvqpL6Vh/VK7+mHOQfD
Ng5/kmKKBHznxlvG2eY9ZvMCz5A7AkuvSgXUMThENDVIerjvXP9zjvBNB98+rSyrjk8VH2ciY4Ht
qwXd3Zafv3Ze2y6ri0vQxwFCOdTTDS4pF3JnC5ODD8HfiDG4n0x+atirs+wAv26adYF/9ohWZwuK
wCuDYgQJNgFCkVFE5oC79KgBHo0hjsOYMCOFxqx8EqQNBJ2eFJnkG+8BbTIoOReuESWGOrTQ42IW
r+Myi1EAZqVsVibrUonipLV5MwvwiHpfHhn9SqLiEi1FltNQrfCZaKfX3fiWC7ILBVBrtrVbYWxK
IzPttQMw0uULQuqCl8cZAS4KTnKUsDH4r1317Ov8J/O/7d9szDADhMgQYyNUwR4Fe8grOvLTfDkX
AoJTmpiv2OQp/XEdgLXLBqMsg/c+ssFHsXI+9owTUjsflK6VA1Bs7Ln/z7PRWWv+ncWgC3xBNbYT
+wdLwwHYCyzXeZbwn2HYIj0FtMNrHBinFUuaZlQv+Z+MnDeV0nmAvcD5k0OPeYJX7B49XdY1RsXv
UtycVGschYvyMIfV7zbyLnIMCrpwtuJANhRqEQt71/VyLvrF/UWo33CJuqL1GOWgY63XPnQYNdcf
eH5q4CmxqiWhKJKfCsmBi1KQPpl5vzy6ddfMKVvKm2/GgEGni/5vHFfCHiH/UJT4giA+8GQsQEXc
ocCXQOU+Ln+FeO2sipoHxjUp6Z6kjRech2PzbiCGmM6843Q//8J2PACCOf7I6vKPdMjzoUMu5acD
9NlobXQPEd27/v4IPKMwj7lQZpO8qJXfqsJI2+xg1GBzlFHDdB15N29MFl3s2v7vuUpNYS/qaebq
B3KgUiPW0iHP3IFbxahzzAvsks0woOJUwhOiKQQYMru4I3kGTdy3DYiBNlIfgJKus9HsomNbyStF
KTHY1RQWD6oB/eC6jWCIu9/9dqN4YS4IXV6YXvWTDVkcBgsR45aCJvvNa9+LNFArrtpSgu2B7fxv
7MwHTv4Wvy4GIj4GmgcLIPeGV/0/pioTLAtd2Yx+D6toYEYjjUzrVIOZmj4O4poBDpU0gQ8lcRHb
1C3CigqWILCAlw/17B1jY9mteZlagB6RJU2PSOEgjpRdBCoUKUJiPJppjoPugdjXLuOBad37uE9O
0YnXIHJlzHXS+CQB8rovzqr/DP/Jsj5qQFp3/+UX/ec3Gx1J9Kq7MnAb4izz3SvgTuZ/2gTysjTs
oOhWlEGGh4vhNqT+QPCEKjXD5fOCZFx1GUhAE+vTyzufpL1C+pzePhN9COsKH8x2QtzJ+vCY0YNw
B8OmeOfNwpbHdhjjmkjF1w1xaKgYZDBeg2aTHSLQU+WFfb0sNlJEptgCRBxdhpBwKmkWrx/u/3E2
zyqEaSrx5ijxaTj7+O787XtJ6IF7YH+NTZwbHbqO/6k6EV4wxRSCreEZhtoT88mBaVSRFXWFtWp/
OsUlJzHkSJ7Tl0b2sOb56UVtmgvy/wUhdkf37OmaOdyKBNxAGceF0I/XyQEbu6vtIzEdPK3Qu1Nt
dDbEoLUKH5r1QiEBS8fi6a3SgWd+qOe02S8l3wRONEMJe+XXHTZvBc0dri+83hYYL5jZ0Ee8NkVG
zWREV+sveAZ6cdU5cB1KXrhG9fm9U5tf5MOWzhhES+nR7KstsrHtq0Mkqys1GKy5RsH2OUlnFlSN
8rgAUqhB68vqGPzAHamjniB5wQW/U2bAArXZKHqvixXlXv/89eH3dVLAN9pMJC/3UpWxrpGuP2ET
kZYlbt719omNUBnh+MRhCiMWgnhD290cWC58qHqK45ik5ItAhPLFNWpYu26CwrWCk6301XnZukyb
zF/S4CDCtoRsT1/EYlpfWT/XKTHzCuZaQVvDdoDO+0gCORRF/W4g/KtsJnt0jPgd/N20X8y6iv/m
rY/nsjFl2W7R1EK9Vbt7pXqSMwQUtf3icEUzsl3syCinQbUWvZVHL6VwziutGUVfDRPw4ul4mXfk
zoHg7/dkl9ULYixDc0JZ9K1NvK0/+AOJ8Hexk6DWDfZbO8c9Mo7rAhE6dGDZPd6juoaYxbLQx3GF
dzWrQCx/BRY3IOLKMXBi1YPRhqGRiC9BBUM8/x/Cme0fvGupmbn73oET35/qJOLyqD/faKEHFXtL
aTzSmoWw0+ScQBQIPWKT11Q9blhR6UGy6cVbQVEERQ/QCm73adSXGLmp74vqgGXV1C0KfwsC9YmG
wxYjH1kuReQ1DGulIXaB9dS+xfi2zixqCCPrZfJppF1K5jKCmTW4cV0VLWhjnY0p6IFM0FIMgO8h
g+Vw1bznTG9XiB5Iyo2ewtiWIIVjLuNMGshI3dEgrC6l9S7Lwb5R28hd8rve3+JdCBHoknz/5rLx
eIP4o2+SW/o5yJyJHzXnYVcRVYOAg4fwMZhrr20bc0M3EUC3KwofWlEbOH90jJK0u5mGJDYy2WDU
2bnNIZkz6dVyueZaXeus9T6dIvGUSZVgVKZcDQalI+/4eT+1cOogV4WmnXmbEP5hCmRYEbkW5ajk
jLHXAljxo8zimwOqsBHQxp43sVCU3hovpkXFydt6s6xGOXoCPC7zz2Idyqw5nMOSSOPghe3EnFOR
DRQbj5upl2bjuN8ardLr4JYLMNDhrcDs8dOdXuB4g+D6mL1RNG1H+hoV9o4MaHO/BLXI1IqniAq3
LWTTbwLacQzxGtYjDdvDNvfDR0qwrN/2jznnnSt+NhP672APoQI4ciyDRTg3dtkSxyy7cYy8A3t9
zLPoI22hfBt9AkF0rCi5xDb8zNiy47YTRGxGPGKF6yt2EsdQuszzeF/tlOcMUOm46j7uYPnpNM8c
2bcMlFk7fWxYPI3nfynHPm/PoFien5iOFwlzpt2j7zSA40Vfqji1H4DoqNnFUqWOVbYQZt509Qlf
T9fnPTEMby8hE9WSnm/2Pb3Y8XBCu8e9so0sQtAfxgWjafhtmVzXxKGaRkXW9KFRG0fhwLBblG/S
hvDgTAfbggwpCLJUiSUM/u6uvFByuCHXsyaJDLOS7tvQ050RhpUTF/49UcoGOlNRc4H71Qn2StCG
TQXz6zn9zOzy/7NdbA2DwkzZwkFP4qtamN6P6RFenmZdMJotUBD7p1fe1jCzAsLYWINAPS/FmMQ1
4IUQ9loc8H2B71x2YnKKGUdmcEV/5eCgueioOiSVWPC5AUUCe7y2J7Ml3pRfiFRXMbFJXdZEitZv
1uYVyiwLqCS+8OEhP48/q/0qih8DjSvd/2GJ8xERzh4FwnnkmmuuTyCiK6UKMEt4VdV+inILTVni
WKdI6Px9ap32SsCMe/nvPkfDk91AvCiSsqH1rtSVqjL5vV5Td1gFM8rihEixZ/KaTpLUqYA0regm
iPahVOCYDycU6U79Xj0ULkUD2syOQ2JIOGe0E3aV6RHnSG4qP8JXWyfv0RmuuXhklvVRzo9c8t0g
Dn6Fza6/sWalbNNokx/uSSBpPCrhFfdp8UGyjK4hoApSi0lYamkX0xpX4kuFvft6VdDhcbb8l2cD
DFP1c4SjbX71LwhY+J3Zn1O+RPpR2nwOhY0rMZX5gvFr2+AL8EaFRjpR4ENCvrA8bgY3xAltD/F9
1bDmbHsHaRcAvpCpd+afAHas2EIJ7sXkWD7NTTfPSug1eNZWn0ch47buMSw5M5Z70sKxInR6/fQ8
rm25SIvhHoAImQkCuWOo5v3JcitUXX1DigdwTUv04PVfBWhfhrIiJKpRELn7/yKhHBn+uRx++jJp
yTH8235ZFqFbjfA6et6yffPQKzcEnpVqksTe6z9KoOnI9V7xzx/ajpl7gqmcds1HGdQomins8TxY
vAUQ1htKcYMCCcImtoROn9AbK6R4g2UiZV2XCGz+9w+CW3QPRp18vSzug6p+Kx54XpwAeqNP9Wja
th3OVrsy+tDe2vun6B2g09M8sNuPTY3u1lOSWE4TbhvAYh6W33lVYhVrrczEyY1LHSqvRhp2+yOO
KhdKsuHarr0S40oUMolqKnJfUOKNOEz7FEKcQn4ivrWO7lCF27Yu69KL8zTTEPQ3wUf1Iw7257Wo
11zFKdH7n/J2N13S3st6/f7ub5AWPGS7WFCCLIjkpeIeGFT87B0U1VN+T6IE/ZxP8IOwrpcUrZzH
ikucIK6SLwcK3HbWwXAGm2AlmihKyS2lC4RxOc0iwjjj4nT9jYvuh6zjHH/ttOP6ws3dGP6MOCEi
4LG6xFb3OwiLt7picxhiBDabDJ3KsONVyLwIbLVcr3d5m1lbjv+Hwep1INfYBETZ0ITe1gilzb3d
uW1zu2yp+bPfW5fYjRWJSLoslqRIrC56U9383eNsSaxRZ+EBo3uyf41EEllk9Wm3UhhHEwTglJMf
mXuS3HEZkW2VHOr+C8HBAHuwpyGDgljH5teoRCnLyUEBO80lZb/pTzL5NZTo2ZmK08OjYtjQ2Y9K
TX1PwxDaym8Kc19CcxxCv+Lb0GPvmmhr4eMlFlEo7Q8f5XrmVS9t9o2xxM3IOog6VSEq3+zXg710
6c5Y9MSYf40QTsBL2/SR7LWtutcPqF/45QIAP2HypPRlIgCdEaHgH1Ck91TGt9Pju8sHmHxDv/dC
R6BvW8qRSyAiAhgdEGUDa6XhNemPNzJjCR+ncxq+sHLUSwyOzocEm9liHauWbGtx8WgwSWd3AsFI
wL5HJtoJVFJU/2aPPy4jUxS+ykqkrZ+iuP2LBekhur6Dn5sb3l8M/d42jsaZcFi+CCull027du5A
PC7kX1z66DeDV6PHQsADfkNiXV4ZwH56zswqOCMoNx+rD8aTaazLFf7QjWzRqCWZWX4+zzHXmURI
RNv1CGHgyaS60VHac9iTg3dYqAywL8Gpm+CCTKJkRlVF/9w4ujaskbWIs+HVnbC89M26zeMuCPSq
3g3PDcGyLBQx62KKgAbo7CaOsSfygCZ48vITuduK6iVl1YMNwo+UUOKluQGlKCT1jpCxxOoUJrI0
VPSv2t5OMSWkKPew5/cXwFaZr7siv3o6tm/gkpvxowSqUL9Y1xua0BNkek4zOzxlMhl96Yfw6tTI
Kw8OHTE6/WWIXGAnKnpqwqKs1lq6uRWG/Upd7IHBWiqnsu5qTZ9kYsKKxOWgvWXAyAm/uUUH4r0a
5C+DaHQzRVZ9iXuld5bF/nJseiv1s3lRI8F6uEu7rDZgK9yHTsi2e2wrCuTMEJtr4Sb+Sj8vDUqG
qb5h4v/+CsZ9kPgLD/3ItICUNc6fecncOgbPjl97WwJVNbUgj+v2CrTkCS5K8GaEBw6J3jBZtI4P
rCqQwHyK7s0tNtt9mwHdCQrie+MVRczTaC1JvCZWMSPSvcKbjzgzDLiRORVC0rzBy4uRe+U3lf2r
XI26lYvbvt5sV1x4x6jjyaE0j2dnZmE/+DER+WocyqIA91PreijjZV3wVp8ndk20fDgXBS9jlNaq
i9CvLteqHHD3JHWSFWqbV3o3HmGBZbCWAamhEQ+e9xoXX/ukZUDflLHXvbaawAykIDmAM/BKXIes
qtgVKFo/GMP1TuQpdR8y6bE1JGcWXeXO+Vg5Gp5q5v8/DEZgbYTc770sB9hYl8yGQH2JS54xTB+e
/rFnFHzlYU+EcJ4LzThPwgjXBdDIYNO4pjyudGkg3eijwgxW1rdKgE4CDRi+lfFeJzBmAQLouiJ4
F1/ozz9ZOg2B5xgctabhZIwFOvcqQXfDbuS67sAv/oXO5nUq2g4/BoYhcU7s+BJyZ7j0K+3/8EM0
DJq1+cDslz1Ibc3anmZBx7G7kj7XZNf5QE5QjY5C6cGnyLI0gcEEo2herBE9U5Z2m5NrPnpIqe5e
7LlTZob70emHSoqM6votYHy3+mMO5jNlhY7gNaQyuH0w0Fx5uEaij9gA890Y0cHUdBAgXpxKRGvz
ak5yTbMMCHgXNX4NA5sv4zpkxRsajQQ19jwgOR04ZOmYgcz/FGeQQbbN9V2Bo9lPQ/pUex1KutIG
LqwIwL9Q/Tdpwi1nnhe0ejDDJHl4UD3FeK2xPUX5ruC9uBIJnyyNqq0afdMf6ADhXXpcbynCHgNL
wWeNFISB5WO1ixn6+waFbWP1nLJ2hpMwxMFw1kPIGSR1CjL/eNrjNI7aAWIdWcs2vjvZoVSSiWGf
Svi+w6IylcDFaSvej8fb1thiwmoVm5eyaoXGck1QV/24GqVQyl9/SB1XuCVmCwJuImHzSBcc98Q+
ilcn3WWhazQIzPs+U0SOAPxFimdhbQwK8IoocqgqFzHnHW531QAeRE2aW8YyqU0YDmRNrLlYDIB/
5cAJvJdWZm8gz9ERiOfH4Z9vX5C56ai5ckMjGxljNFHYh3TSnrjk4WhRs2SzJoIE1qTUJ6+wiklF
e2DL/Ig2TqsKRCOATRsItzRTvpb2BpnQb0UXrt9KAP2B6+Ti11JDpw56bgcwzIFUOXn8qZtpyrdQ
+FYYQI3FrWWv9AZw1nHgw4jjikKrAs6ijZUF4YkuIkw5T1Do8K/OzjxvUZXzsoIzYurH0gfBpLMN
SqzPO0fEF+H0NoP1JT3BUdJARxvnShVt8aDez06iwPpn1fnTv4b00dTqXuJ2Q0vSqmBsY9hwQLRm
kAW1xPHNAZAt/CYJ85XJCsGWScJH7Ec89i4cpgGLFAt0zocrXrDjAKEsuXxwEsjUB4whVmPQ8Adf
AUZ2Uz0aI4ByZuiDafjc83dIVbu27dqfi7J3NpSPjXGgvQ2xp3yswF4wQbAmv1CqmtamrT07RE8p
CfjQZ7Me/ZtXGK6xUopWzle0B/j61j/SzcuxFkXGxCwM4lq5s4eXizYGRAB6mu230n7EScuVOpX7
kPUKtB1ekm8aBheTVNFXRFO/nv5ckknvhY81WA2YqpoHdYOx718T8yhy3m46Dntey1Ql9S+sNQF6
GzQGvZqFjZpxyHt3BKc3wV6hk8SMcyLTJj5u2Qst1SlijnHTmaXbSeor3gTcPZdEsxC15zu1cOoH
3/3G2PBL/BLj6Y9ZGTh3sWscv19TRIGyBKTiFDGzlvvfn4kQUDbfiKH9Ymw5jN+CdT3+xKBzRTDH
dgEcyp95J1efKsSU3WsFh0yB5hwEdQ20jjJfCVwn+OoaLqZHKIl7+66Mpoxz0EfBH2KZD0QTfSaa
abof/4Ghz/v+1AF8kkRq3ev95qhZrUPMyA/jKzpIPB+I84TsQZMcOV5Bp3nXhoEfDMLP5jokY6JP
/E9aMP1ryN36g5isYrh93457xrYySXxHeQmucicHXFLzlpozNa7tJtX0MEsMP7YU1wL0bC5GmaIg
ZKkyvNuQbVGH2rdAgov0N0Le8tGrUjXFuydTCBRgL3kh5tskjVdaNwUCdgZEru23+9e0tLEPWAfz
Mf/E48IZn6NPpeGvEBv5p5V4TQzBFstm0mWDmIY+GN7mC9GNCgy+fI8ZMNQ3++b1SIP3SlAC1hBi
Oj+gPlj0F1zuRiq8ThsRJcDVycdV3SMyJTHzKAel+X0v5bEcpMpnYFSn4z2haE3LPrDn6WKbeYb1
uy2emVCvRjAoYDNkEeTLgpXnljinYpX6DNhtH2LDM5w9o4JIKtAnHhJsBzzHTulSwsNIdRDSDHXY
PR0gD7XMWEZTlgRpVJSOBptk23lf1Mb+k83+NOlgTtIiSsHzKI31NNMedmMhUnOj9VTC2CSH87Rw
T+rArd5wXTzHOruQUusaCRztCMYCcfBRR2ayn5o17KwLuFvbjd7w3NXcr06O/mRWL7/XDtbR1ctT
aLieqFoX9MrwzK7wi935ZAZ7ge321DebBlmm8EcTbf1GYXuKulyM4Hccgebf0F17zO6Ql30gobR7
HoU8NRuuPWjNHLJ7/UJ6fLOYgiLEPZJHqeK+NrW1G8NuJyjrCj18om4U1fxk2r1Y1xbu1bkHsFtw
81d5fwl3UB+xLRkxACdQaPgH7djKnWF0bRm2h4vDCo2K5Hcv6uP53ZPXBXati71YSHaX0oM9LVfx
+guptxf+PCqBkZHCwkX+lxL+lAe4pW9ZN00Zo2zPuytrNdQQ+fdPjl1rfzTm3SrQm1gzs2NIdd3I
oQGsVRu7X5tqp3jtXYTViyWMf0uWRdGLIwZVhLndKCvBkV08L7kzpaxrK8EVDnsI7Wx+IaGv3Xif
MXRpvtu/BNbiEZdNTddGldnrNhBF6plUQi0OaLVkfA3otg9vxRYtwVkNMmZanzf/ua2hVPxYkWu3
k/56OV+u8xRMJHNd/GPyzaFKKwrAV2bCE2lQfe6WWVvqgRVJVFANUJH37zxbUHmlrlRfPIxZpDC4
uzLyIpGC9mDD3H5tddFwfIs94Dh/L2R6nAH7cwscxFXbC2ujWCRB5uc+9Lk15syAMDU/oGeXuHX4
JvbLuDsp8zAFgIHa59E0m8706oij1T1br5G7jxX5iHc+DFsiE6SfUapVZS32pMJJ8yhdN2FCv1Eo
qFEUcmYwpYh7aXPs41bzRBODm+SOCttxL97rE7wO4CDYrl/n6bYhHKCIQtVgGiXMZbpmBCS2NdGz
qnrwljHKKLvDbIscGMRnLqWaXefaGdKlZwh9QiDGbswuAF90VnheDG3+ambJIdJJiBNRn60+3Jb4
5oMY76ppbd5B9WhKHMomx5+NAND9KQuYzZDdgoUvFtbP/qTeVB8f5RePdHeRJMRESjef+xZwNKuZ
/0Y2oMwuDpn22seUy2X357FTlMx2rvcEh2oyltWMp5HOBKLovALQ1br0J6apEJdDuHh2sOW37SH3
i1WHz5bRNN3cwvV158SuT6GBidAV2On1JdStSrP/K/c969T2h9tOzXEabcWl8C6WTQM1QpAMwpB9
qhowcs+/0sPiiaEDG29opAr/XvDMX+RaNGtLLFIw7hGIbUvc97pi4LmM7rTrDtWVPffIL81qkIVW
nw/iEj0WHNqk5jeHm7j76m+kZVB3Yc2oDG4/x0LUkjPf6Orsld+ygqUZRcIQ8veHaYCFFTzoyFJ3
2FQAluLZ45Rkr7Dc5pJwnhVUTfK2nOicIiZwF9SxtM8SUUcYfx8cMigeXCt/q+Pnm426/Q7h/Jvj
I+YQ3rW0ACgpL2mLofwlnykoNMkXD10k7gcydmnT1mPCw7N0EEAsYLCYGg46GRet777e3J9VM0Lb
hcYBTMO3seIAZgX8JpgX43w55FoNRRgnlvenbdPWwP+02OFN50Ks8c5CWMfUqTC8Vfg72rC3Y1Pb
1NXNpDiztqWbcjeEem6k/fvrDWGBCIFoXRE5ngJuMEya5VZfcx9PXnRw6bP7FOPfiUmKMKFi9jMA
EuoIRMoJxuxtfLoso/+rdIo3ALvlyoJTL2vtJd7EvPUzqVYH1fH7sYrvO3I+FD37m5tQAcUKL7Qw
kTDK8dNMJB6gzHsFyAZUhI5ZuXhC1yVcM4P5ZC+cDR9NA3U29rz5vhjt8mQbcgXO+sFNWv9HF9zG
szbzdAzkUj2Em5vAMJAMel/SIV5KHpqz9QAKz78Z7WIKYA6+ZgOQwikSiE9BzDb55irIlW9ss9TQ
Q56j3JxazU+siWCZNpf26hJD2D2Py6Ec5wDHHqSN7ho75LdgOT81l4/zUtdvoBZ5TC095Up6vOp8
3pYWKPAaz6xKfkgpknFtCO1/awbAjGZl8XmHA2nigBBTbU1XZdOf6TBf3gG4Xeqz9RT12M8xbP7e
yZuXRJAB+HxIM5t16ikNx+CMvszxfCZGxMsC9/KeNIMs2S2XA+ph8DV3h2DBG6q9gxc+YsM3Oy6I
a5dDpkrhyHx4U4YJfP4StvUGrORvirF2C7xO5qjeLe3xQsUFUWpV1tNnbVuXJ6rgxLdv1vDaMOKP
9YtED2VFCHS5gD75Y/DA6qSJkTGxL8v7dx3bT8CEyk8LbvF4MQXjocUJBP1vwlo/EQUxpDuUQixp
JuF5d6Iph6F4jbYFmo4iFRyBMC6BODU187xmohLHINe/p+1C/Djpn7XG24JgEQFjsPatMAamaDgH
h/n7uJrZAUoysmm4kodpe56q4Bvn1ZXAmZpuW7vbiwvc8Md14AlEZRbc34MtSdDcfUmBtwyEIlL/
cTJzGlkwpQCkhazVyLg4usfbl3qfYkhBFL7fXfAxY+w/NLOFR8wMylcv+vnfEmuiUuwf8PCLcV0U
OZJ53nt4nr9SW1IIdjG5KlC3HDaHt7hYKR+GS7TV3wSZLjvtpZKgrWOn49bT6AK7kXG12uEi0s5q
oI8tzLbaopm/9B74kIqK7yzjwKlXBd1at8f7PmP9ptvzLzBwSbb33TkUl/uJe+EvrSxQW5PYoqQB
4bcDUkH5MwPMcBgKQ38i4i0uSWV6Svp74D6152XTniRAB5qk4TPQr0LbdSGYuCsmTUzlF0nW4aqj
+Tl6Z4rRzJmDQpR9EJRz1+Xv44Bm60LDbdC2YMH+2NTdixZP0W3MpHqibNdIkKd/HBwQQYoeBx6t
3CcUKSyfTqIA5/Q/wGdyoUjFU3fWxnkLG/jhpZkUsKH9M+AncO+sbabLs+527mPifvLc4RZDKaju
zfJu8SvE9dgDPuwtxV9HAE1qgbUH++TaBJet+5Zhtnf6YO30FqH7urA402hqy1wGW8qD4Tml/8Pi
yWnAwl76NvpXZBZ/ZJVjzLkaJeLpRDVXjpn9AT5mP26j+mVP8sxed5PoZKSdxXGIZv2sWz/ztcnB
ebZt+ajGuWVjewUGDlk0S0uY8Pc0lizvcNhv09QbFduFzKowURR26PS+yxagE2DkNkZkX3AlCOwq
JgrluVfiYpD+enUis2tL6nJwU4TAERAevNcvmtMTr3nnmri61gehY3XgBDi23IUa5qWQStu9Vw5n
32Twhn3NIm/9/SoUnP+DyC1dyiFGpOFiiT7cxQGQkszYttQIUTP2tzA/IlhgonnplO5XuaGyCBgG
oVamEdHlc7EU5hNL+U1xftg5MxPZaaHDRKsNhUxJO2Ck6CUAgruxFZKfpUarS9LfZbDka6TkzQjt
9zDpcXwn74jWbSYgbIYgmuL5YW5haZBK/sGBCTzLgz/1y62YPuHmCF1n9vuy6eokuKyqZ1SRqZmV
XdmEo8lNMVW7UBkV6TReGVLvtLnuMOj14FDyzTidSMuqWN/RJgRgEX+0SDNPaQLVcK+eN/z5BIIj
mvQfEwm5Axso4fR3ysdmBFic2Dgd4LQguQPgOLRWigHeuuqNfocWVFL+i/p/tDThJp4sOloVBwZQ
4AMNr5R8LxcA8Zgz/iOIU6KMNkhSF66YOB3dSVOHUjhFQ5+HCEFENiCYlReKWIQIg7dLc/ROJARq
4v/Y9Yyr/JfV8Y9lePhVcIUIjzHzhlkKbhtcaoQ8MNLrNIe1tr09E2FCn5bqBvXojatrgn2GpEBE
s56BCVceGjugmsO7/RWQr37/9pLqGWxL6tjUZJ6Esa1wAibzjgtK5wD1b3eIAeV+HH+7UtqyZkIe
rYb5HM0de3wTR7+zMryTpxZbG4DJ28AClwajaFh2CofVxClwwuPzsNcQAjlFRkr8P8pBk1j8xHNb
Vp37Pwj7SY+S6Qd0+eg+UZmUSo6mOHFVGF48hZyEelHErDMFrdXo/QEsNuZWC1cxM2jaFeH9XAbN
CxBfBxUlpgl413m5FysfIym4ri2IjtQ47u3Ct7MCVDu4jGZyJuTTkSsFZRVoPkNDHVvpAkU+ZV2S
2GCHbANm24W7R6HbLBKl1ZWBJ+g7N9WBkpLkkJjuoGMKXaD5W9d9T4oYfSBnfYSS2F8BcubvXQpd
bfvXjH3Jdk3Jb0yQh8+ZvPhJwxwEjHR8GIFIkqQcm56Zqqn/bz8pqNke2mVm/xJuru8Fu2yzxp/+
pN4y77ejPa1SS4fRJW7qHM6in9ig3LsX+hk5M2ddc/s1zSwxYx4xEpSt/vp/ySPB0odPdQukJkad
1KpM1JDOQt7JAf8GExTiG1DQ9IbCy+ZiIu3EKyK57M5e5SOMbYBoEpPeuXF4T+dHFWb1Q1+/G3Eu
shi9baBroreDx23ifSf9WM2wEqHhvJVic43b6t6ILpip/gowNjxdIzHxCcrhar9TsDdKUhpRxX9U
1rsSIa2OQpDTDtBFWke0bmCvePWasNWfTgJD5ERgNSMoC3oEiCOjTMt4q0ck1+9depzyrbqf+LQj
8o1EuYWm1Xgmfx9rJi+lAzWqoJJcZQ/6jkenvT5+HGirQaaWk3BmSgbWX9r0nbz9KbjqOU5g3ILI
sav/3Kuj4WAkZtinKtbDsA5c31GNjRmAeDapPZNWRfGzpsvQISXMAlTycZ8EBWHp6DQ7ZTkspIgg
eTyICV9zRRiRWdl/Onrp4DKeFNNWC6Pksdml0FO8+kZeBSsFY80P+Q/r54eOIlVekFHAgn6WsMaA
xBux/LRM732CJESuTjDpa8oeTURrXxFzpTz0i9+oOjYXVFn0XhVtpjuJfqsAwuKHS9sz4+5ePqsC
eS83Dls1sl3jYf6k7Wso+RvQt3Ra2McR2/m9AplqPBmAs14loVkMmOZlqEy2Eh2ceP3NjpoQ28cJ
nyJRV2u0cHQEAo6xg05AsSi7V5Kk2S+INMLghvkQwM35FLgFqZjmKcYPjnJ4d6UwtjIcoVfsZr7x
CYpTeMTBGLB/OrZjkNQM0UsdSFRwOPIMlH7vPwV5ryBzqUeMw+KY85/ReJ/mGEa3PmpNI5og8OZc
D68pBsIvQEhb8OHnwB2i9SpFE7SPONkSJAZhL9HBzGfAK8qd/1Lwlr9dqhr98mMiMdh+bfFzOlqr
ka2GOxEs7OCXLlvjkdGmx0QhmbEHkzdm+FuW/QBInuhVsmGnKF9YIkUcwLniPCkdXsYjm88/qG2N
FKVf/EC4pC9Qr9iCMnBjuBSDT0xQPtagsRaTtqklubZsj+WtamqX1NH6pDjM81rq5HPokLYYj0L8
gKPJKavbRwauNYgcwo72ycWBi0lNuWdWgS2t6UY5DoMNfcqxqn4/2stUqaQv6zumnTO5bXq2ypYm
MMX7AZj2gnfkMb1l8R28alBv8i/ijCH5NYUgaI5DopNRUi9vN+S4V+jnGzGrXJb3PMFj+GDe/qpp
rQvjMU3KdluXczxDF0qviUqMilT1bkT/QuEQyhGk8S4eXV0C64XjoVK2C/usMtHBq4bMqP4mJeei
5SMYVtroTvThJgnw7fG7MC638NSTk5xw8TV9taejOV3kqVCQUkw/5Eol9HwZMHBHHehPIug5FC+s
dT+7FRYEhEbyuijw7raLpYRTMce+sHdmTuBNdNcUj1PsFnKYB+R5nyZnHEdBslB7BXRmbbB9K3j8
cNka0muPU6ceTu9szZ6mAV0q7Tbf8JINpw6q5iSqBJqtb/d3zE3FFSDSMgdSTqFfO75hvnCiGC6S
JBqyJUta4DqD3Gq0TkwuVliFMHFKWZ3Y9IzWlx34F/hFw4dwyggWQ8S2fPbi/Y/uQiQLSXK46mS/
vELYPMxfKJJCVtqJhkTfWYvJhmQKNoGvjU8adRJxoNGc/NWmQxUlDebexhLx6RsTZOE5OttgLDgs
PZLC2zDiplJQsCULGe2mrdCRuaWWMd8LpRQjDvWXzJuFBaDR7RSkB/abDfYsab4W3TsnaBZ/Elof
B6OhTSa9cuYRvxIwapmyKyYgkX11PcLhp2JOBbexcOK32SiGJd5q+oHt1rPE541Tkkj0ZSkpUOYA
7ELFI70rFNUAsaOkPnET1VqKqsLmJlmoF4smaeLjK4Tb5URiscp4vrkQrSUvFgpNqsjbNyycFB6g
JOG0bvpZLm5C2Rnc69W1w2bJQcvxENH3hEIAA2QQ77JzUeVFAKoinkG17SBDnG3EJuohKVQ2cuzh
+CRuzz5lpfJiuTxS7Ju6EtksT5HaBtIn65wsxjFY9QPWe5loynx8XEIWKqk0fvZkVzqoZA5OgH6I
thEzHKvbp0r2cqDqtRbGmSlLDzBJ/BU6dI7o/RuhxRU1t6tcGZdQRDEUN0Kzo9vBmVTOFBkU5zzQ
r06aoUNgIO0npVTWANusYDgRlyMbyKzZg5GA7Fe6qPqnxCB4mgIJzwl/E8UwGnmJvZ/PaF7OCgPb
hSMjKNKU/3exsYnLSEaMAat9rhAgt6LJxLWAfLu5n6c8HGz0wEcVMwqL/bbnoKVBO2HwP+69R8KV
QN3rGUbrXyk6yD/ErmB3UrKYwz+iVTJJ78WhXsZPEGH1+mWjeLKOXaKayA4U0EdaLdCDm6IoWnD0
WFHLSJoR30/0nCCX9HqOr0se3QFCc/Q7hHhK9v+4IlECrdAbbjG5Lvw9wyjhA68GOFkkDV+iWgds
P5v56imL6Cel+sVRV5yLBh8+G1uGocfG4E+4zDjvPpLbIaTNlhKKs50NF2RPyjNFE94GjYXP+U3B
50Y8StKYD5HafP0kYoo+XohcCfyYK6cdWMVSGdym40uc3KO2vaT4YvFnj9U3zzQsGlE07SWJCqRr
a7+lR8y8s4toCRKEf3hA2lpdSjj1RS8uBt3mmjQDoYGEdyxDDGGsxHYNy5pZ2vOi2O89PXEvfLBp
AaxbX2Cr04jYCTM7RbznJ4NFIdPj8yPxweAawQGv7ny9RxUFYwpaKXVirAS+xlhBKqHL4o6Aau6E
CZCo3RqdV4pvJ+BsjhKb0k3Yy+vftqo75mx+DQZmV0blJV3j5RoEqy+LDnJ33t9HjD5331euzQIO
1kQ7aKFW6R7uCxM0DypBOvTNMiqQeuQkU8on53fAfMRIK09y99nT02efBxyZgcS20kTPj+aplbS4
4QcxugUp6PrMNH5bQ9ZHBnoSdikgwTpZgC1NvjCZlSekoxTF9w5t+kWKqAGxgbeTCT1DVWtDe767
nW1D/j+ykstRGKypG91rQZhWLXJ7sT3q0IuZQon3VEsY/RRHTbEsfPkjhJINhKYbgtgeZ0tvtn//
CmDMm6jzQl/Kf8AWp2MRg064e2O0HDSQ0HcHfqHv+wQjxpOdmQoXM7jq5t/8WIj85Pk/tJ7Nxq4F
ze4XGv6kdPSvOYPxsY0IuPB28COaLHfKtzVQzO8fXGOPL/+dZ332g9j2+sW4RiRd1+XI0pLO0hm+
xlZaIiP2TkjA9kA0gOa7delthnPFtuftkEpd708U+hODRuZDzdcx481dgPvl4K91vfRTiOHbqMxQ
Yk2SE5d1bYkSz/FigQ5GYZXmKanH32xJu7VMgI74HGzsHd9SvX2vqhpVdg94SuYpnT4G4MJT2/BP
cQmQd18g6PkKmfYQ0+C/7nwmm5PAk8F0dtd5xZHkcWLTuwVLFPEqTf2IB6pUmOIkGLnSPh+GxLMm
aqJ3VtrFBre2qovi9DUkmi4K0fUtETzvWfyCAplBdpXurJhXKMOT/MSAG127WLcrtUyV2M2u5ELd
uiQdK1EoP2NH/h+bh157Qk6j0QSpzydZ88W8r0JPw5ZvYLRBUm2y6+sWVTHrrNURGHMRDw99yEn9
odsJAq49ZMDRA4S2eXBrxKqqvrckw3MZNOzlQVmf1v/+L5C2yHVlrJnyvC7Z+pjgeanKe0WmX5Fr
tAVwa758ZJZAX+4ns8OGMJP3XPyJW4o0H1zav/CF/k0bXLdu8Fon99w4TMLiETvWZidUksiySGNm
Za8EYCqF5janOJ6hKE9yBVHP2IpwWWXO0gXDt2h4eH5NJzbXR/eJGwrgHkFs5n3y6HZkn6o7LK+n
BpWmfvYqjL7w/RP17EQZKydRK5yFfOtqaLxRm1JmE7LGG0WsJGFbbYSnUuctwM8QREFQ3WTCbiSa
nKNJKGd05sXLoY32Gy+Npav0SEGj6lXdak1ewVKue9wCzo9DkpvcH76rPXxew+h0lo0pzRgNDdyc
FNHu5L3OgckNRvdsrOmKXk/jjEEjV15L0dW/XbEUkvA1RLnDJrGtRqkpVZqySJTmuc9rc/4zdYiD
ZNQXoS/VNEXZ2tp2Dff5tnQXqYnIWFxjM2N/mpwmP4i0BJ9uott03BzTRRdm6vZMmDgK4bnbLoy1
xSwFp3/wz/8TTy/1Z+YOzz4Nhwt9HAZuO3ZsEJ9CkvGIqYq+XHv2oe/Av20gvWPObxsFp2bPpvYL
PXba9NWykwzPQfzHXXpoK+CR84YsZKHZ8ICnMGrfRVQMYOKOkKQl5XWH1bJQMIx8y1ox0lr5j9eT
MnXgL6x11QKa5jZ9dFGS3hecQSVdgwyrMGiD9ZWMmNWjT9Gm7gvs1UBCfG3E1oP7Jlsl+2TC/ke7
bh7pxM5un80gEv0TUdZCFsN5lxBD2e0Rh8x9k1MbTKBKC2B7TAJuEMYq5AfCNxdFkikmOAK+r//k
vCygO+Btbi1Vv0hS1M8zP7fssxh4ZNzLqmckEBy4zhN2YR8k2u5sZnvcffGn6BV+6nPuWrJOeGxK
T+yOsxW+f1vE6QHRzYF2R8pfZyzfR90tWE75E5b3pHqV5CZx9a9yOorvmrkfxraaSyyp6+Ut1OBS
P2Js4Oh7diaarV5d85XBGlHruorFNnOZ3zAVnFjmga4wagg+l6oDhP4MLpVk/8Oiv4GpKkVSuKpA
xrtA0nwWqiGDLHD313f5r6uMF8ez8t+7WvaQ1tq+qButJ1X1YvZlwr3TqULOju0mB12SmJBG8WNt
1asIV0b7we/rpGCQ+12pGmf4ZVpQGIYpUBi0f/6LB5ryxeKXSwLndBI9VztsAzAuSzNBOCJS9mAp
Mllxc8U596i5b5aBE1GBPVUOZywHznvyE6gLEEWj8mGlqK64zMr8RwLk+3ZJGP2BXnQ+/TSu0UIp
dXyRjMa0b4GNfCu8TQhpxswe6J+zs4aiKoMID+rbXmJqiBSJhb1/e1x/LL9EwYyGeRRE1y0N+s1u
c/QK+JuOOXZAY5bPsZQStRklUcPQV3K2zZWFrKLazr31MaoGndwI478kGuCbtK+PFyqw0h+h3yny
+4nUGHva8JI7LjCq81gUhG6TtpYWCy6WOcyZrqQRFNZYo5WWdWFeidW6dznCJHSe/8VZTtcHQVMA
gQVMjy0gFr7nhasEiJEcno6gbWOxXYnvNKoXM7yGCM/k1UXt95WaA6rcUvU4gBjTRM8f8MlnKT3Z
Av8ipaXLgaHDGlGiKHHxIOYLU59LxgdGUQmIyottHg+Y8EwMxZj0F5xmbrST6WGNgKozMlILSmA3
pILWz//luQi4wXDEl8vuhVKCokQCowBXV8TI2IuN311OCvfSxkQnefHwEe9pt8cHRy4V+YzWLkyO
fgIg0e1AvY6cgrIHZ/MuHdkhAZJzebe5NyNIv6Usibn1/w/X4t4hA+CJnjm1zu7L1E/G+WAoOIu8
B1tfXHY5tgFKTNmpkNnNeHIIfDXisOjwBB/srh7bgIQyhXfoUsaHE9tOAQUIV+PGw2Bsv7xCA8oR
NXaK6RXXiv6us9Z9HIlHcMZt81vEf6jXWUgcsqH7YxYVlQuzP2Ht2+mS881X5YdxaSqzVK7fajl2
bZTYqcoEuZkejJ7bnrFGCiD3ytne+XFaxQDeSIqnka9SxoXDXODDylYma7JdIyKYr8sW7oQ4bOd4
Zh8X3EqPYBrgOXeBw47aGDdo2HEczQRBQEO7WgdZniF9h+Xr+AhBdaAfz2KMJtxMJ5PdlEoF8IQB
dmldWMduMBe1VoBZSbMHagnq8UYFy6FdJi74vvjFUiYA3XVRPaVPsc25cacwHgHar+lG/Qsd39E0
RVg4BgPmQW0LTjvGIgP420fj2wK2ssNoLVl7nHeX3bCIxWTXvyAYP7VJcDwrIUk8XVhQV7etslC7
Ex8rlX7Ep5ZnqH6e5gMXVDeLG4GhagdCrIePzKRlv6fdZX3mO0dNsSjoN6zFeBO554RvqM5G0+uB
PJ5ZfSVcZnjPyP9xw5bedaPYMTD50SjrMvmGz6Z+tn6JXOjsW69+1yRJMrhAXWr6dZGI95lb6biI
Ou8o73IL30PtmbrzuDLJPQs3rYhMGtDygpRfuRRw2BjIQulkIyAUfp8/vf1sp/dLxpPiD5ihcDev
Jt7TUwM70iZ+Ca9VXGHC4MBcA0lMt8+f7vfj6Nk+tBQoRKkP0sRxLHVszLqojXJv63+00e53GH+S
MIk0AsnO/XjJ8V61jbb4R2QVO3a+Alzmbm46hMwN17O+Lzh4rO3EAEl17reioQZfInk8s/InXQAn
A74PezlnqoHF1ccxhh1C0wR/xjSahbbj5/ttFbasR2uvCGqo6C5R6imUe0bRCTKHD3KADVJz/AOd
DfwC7MjA2QX4+XAmEa5r5OC6RrwJYFxU8VPDUeSOl6eqoyQRtwRDQJRKNDQnrzwyyMr20s5NhvEU
q6ZPX910JfIDp7Hvl18eyUzP4avyRILuEj/QztuoNwsx/kwYE3y6VZ6gj3yY6h8fljlfr4/AjyrW
YgY0mouubfwiQMeazurcnCov/0dMSLMXDTSxj2VKJG2ocOPaHZIZcisLRZHd8x48xv3ebsT2zP5X
96H44KI+6MJAmOXmljLv/GVadKNs5+ucgxuh/mkfu+17HY4nURmC91hEQOQx69Xq3b20vuuAnsRk
609NYJFhfiyMtInEkd6zVeTyOU0sFwUeTIYt8hesjppvCPO39mXIPHMHqRClGtvXktX3okYoJreQ
mJ89RpA0gyNJ8Ut8f94ItW4zpkVxWEnG+MI2P9GHbRkxYKPWWMJmIJkfJchJZ6Jc5IeHGzMnLn10
9A/5riFuIUmvTFTnEDgmwBn/PUAXwm2VCrmC8Y/6ndM50OvtTFYpA2oO42yo63caVN/pwapdX0cX
F7twr2o2OrYHIxHqQtrkUuKzBwpdmEJ/kVaULwL54T0eJZ53+KtPo5K4tOx6Ru0deErlUlZtzKro
PrHMoyrT1mcIaklavq0iRqmLTjf+2IK+UB3VXSjylCZmrawYCKsCUPYV75V4Xx97B3UsywiXCofK
f1miVLvMSQua76PGh8bj0KpKREgKTQwIovwcNmVIov4Nw4s88MCBYfvdi4Ygl+oW4FV4Inxs/VIt
sG11yZaiamjweKjYmAuqmIY8Yj1xARg4EaM+n0Rk4xwLf8Cu3wyd3zMcqGX+oEYxGsRa42Y4ADzc
q2Hdlmu8gokfW7WMJzEIErdk5L+An5r9Cn3BcUhrzx9803jUvjKJ8ifdzDG3ScDGdBlNHXSHOylI
5RbtA0sTH8RS50tqdsAsNioB2hblhrPc0wK4QURRMSesyge9rck2NfjHdsL2GSQ0TmI9KPHzmcp7
CWKu1wF1wbRyeRKIO39NlSMa1tzKde3TZ7mzQDm8J+bq2DzOpzVCqDtzmVeKa1i/MOa/4SCr3VNF
izZZ6XrqbaND9kFBkhuu6vXobMY8Sm0CjTxIylnb+a5gL2Y74vSUT0pI7rWdmNGP2FrLFFkXzacf
2YGKFWVlj1V5I4dR8U3NsemIFOdxMAJymmbLbuFQbHGZ321g39KHOXBrP3nQRmg601miPn1PwIl/
ZBhn/+PKC2cLvnl/5dXtJUXlOYnZnrSvXgNguhaYE21xx2Og8qgYS82g+FKBDdm33ck6OUw0yCEv
eZPuWare/XRhROJlJgiRK6cVLo2lq/OKxp6cb9DkfOkurB/SaBVcORwQNow3Hcn7T4JDIY0wHIZD
U0ctQ4J9B+G164COHZMopjbL/rcfLufwLU/3e2dmt0JGgZfUAKdQKgXJcfkokRu3mRNX9E7DloU/
401nAw0z8HwLY68Ik8/v3L4AAOL6XTBo1iwVnwRjtpw5Sy21UwsSuKfqwEJDstM/Xd5JMGtruk8+
y8pKIHLZNliQBA7/ixdkT2fgFQb1tZxsFthesITokyXGqjeeAuqtUT2ozadDa5py4BWIRpUWCqAy
olbVDAJafa87FJphmKbeGOe79oEjVEb7syItSS2T3tOONwm6f1KcdEJOdk98DafYwGpLCmt8nh11
NbWNB63m5y4tStdefzcmSm53xLPGieNvcaIdiCZpB1cwSZVdJf0vwDwripwPSA6hOOX9LEPAjNtA
81AfLqzFMONrGdTqd8y08xhFctVNJdP4fg3GiH8pyUDh5wDLwuJccZI4lxZziLCZY7E8Zjk6oiZX
yOL8Q6FbbX6HWMsTx6fd9hRE0fpTfudEfqOTiCyjV8pElGW08OLa2tjqRbBFhbBius00EApCxrOS
TjKr5tBJ/zaMYKZCBq6paRCLSIvrX4ojn1Z2QE8U/yaDgucfI5+dA9HuUAYgWytj6Hd7vPpwF3u6
ex8s+TGLXW7NTc5hqheciFIHuBo51AuWBAwYyp3RkCCOJchheokecMkB72+6fjfQFBOfoivbJ4Kl
Cp+AaAczYecx2b9Mf34ZJdgIQlqRgFctLZLljLFgiDN0iSQs9Yt8w9innfaqWq1G1RXkRJpuD9SE
R8824k39uCM07zem5Foji9uduQ+K+42Bjf+0NAXipUcmMXpsJTZo0q3HSFIXe5inFNdgR25yD19W
+Qqo56dGhrE5o60cqwHIHvXyZYF8kK2dK0yQ+e/w8pHteauz/TSfa/+CSf4bl0ORP1DUiSxvd7/r
si7UrJNYzLhDu7zdJRxt3K/lZ8ALrBRotnh8stPdfh+/tcyiPwry6ohCocVsHZZYoa695W61faBH
qkxqM9NMsC5l0hJ/SlxzXOZywK/nmPkodF8awHAGVjO9zzIyhuyTATeyg02gvH+EH+lALDMWEbve
uVjfAtb9SDeKq90+QSZ7Y8NkYzRdn8M2Ds+Ccg8pl8Rd5kzLSJY4ykcTCAQgx7agSj7olhCUsVaR
fr1i5p8Ebktq8eqSvnuG9MqJKxXc8IYGGCkPxlKLD9DXhIOtpCeKdguRJa3RV9lmKhKJ+jEo9LkL
Ng3rRgU3TKzK9QfeXg2uLpvrUHYN9LTc1RU5uBMD/kQHeKJbH44xiSRTq+rW11ylmHyfg3oqHkkA
tWcnsgo7qFFZKOug0sptKgqE/a+3hL9TPwQkhYpTylmE9qqNER8wgTYYX1ZvLZWm5EoBweCb4tMz
vw+do/YrY4YMQ5i6ipnx2qcEiCq365xKJWlZdo4rkrpvCARUW3DroV3AZ6/TDZk3NmZriSB/yWy/
wZ715KzpWPSTTn6wTQfmZIO3z88a2S2ebCo58puPFkZOXn6v6f7oB8DTMgHjajEZsixFfOyxShFv
DsuzgIzSGGSQDYFqoM1nXfPz+uifvzr6wsbIiEzS3e6+lnGc2MzqkLx1uFYpRQw3GYFNfPo5l1Xv
ZFp7iJgdwf1eBaJ98WGK8i8snbU1NM/wo40nppL2a4dPgtZMVON4Xgh4THGK4cUDVEGRqXSeIH4q
QteSTDZrElzJuPENwIsqsMMn3wUn340uY19ZXHFVty3kvgxMXJ5KVKOc0yrjPO4OVIbQoZDKb8/G
b39e/H8K/36FJOSjHI3f2xJU+epSwtYuiuQq/ppWsO8uaexDki44k6RPR5H1xxyvJeSKqguH3kxG
fzJ1QwXLAJ775Jf9MaN8dm4eRKm1WEIp/KimuT32FkV1WNAJd9kdIZ3GGAaY1TBp0CiCWJdEtNjh
oalfPpMsuLielCeqZ1FU3/8XE+QfmMJxk5QVu69XjXOX2xylNd88YUkGcG2+pvjxr0gfziKRk54q
jLQ9D+73lMSJdGYdz2a+JO7DiUUFwBaQuGLZJvjxW39psDxxzZLvR4vmP3HTP/DzvH/sWJt+GiWg
ut1K7T3zDyTIhrVU/ENxVttpavBJ0/X/K5RkSx2rb4Rkc9YLmNyhOPq7CSWz+jcuMWK28ZI1vqhn
7QiPAeifrLf84z+I5MtpYpRgXjrfggcjeDpmwSHQNHh72ai/1ItKWCmgJT0dEnk98Vg1D+dOab6B
1WMCKziFcoukndLv9WC8nZCy6cZQpS0DH+OHElL0dvd4cZno8a3D/q7l9tRvE1OR8spGKCfjj7uJ
7YFvm/lxQhHqkBCCJTFkeZtFxoKFAQ0ibPb7FMDxQ+PT9Ds2ykUdwnUDzoaPLgT3OdnYSnSTeeTO
AbX23KU1wFRRFNWGOELadzONCRBOJnkNSilVtZePJwOJjcLvlEfAGkEiL5bmZdR5Rh4bXov3Xmy3
o8dD4WG+J6ZbTOsfe7771gwwPUjpMQjNtaXg0Eyk2JtbZ6ZWuzbZdrkATVPW5CuA5vccW8ng4cMo
Pjj4xL9SbTDho8r7ZfgKeUasfLfRPcnAbKURz4z8LP38kjC8rWf2++mVhekXb9doEEtbW96mjeVK
0zTYlgW2R/AqDn57t9EkLLviiaXrf0QlITI3uaB0m4blSgLf2woAkiAQUWBp99AotuJfj5wUeViY
Ont3t2z4HUfNdkeqMvZmwya8QkrQKQ7bOFaupH3ntKXXeb2RRUfOQYi9AqgE7g/ukz7KDzINHnfo
gmuyO6iA4B4WXH1ZQscW7ujyIToWtTBMUAsn2I0Llg8D2epiATEt2gg1Q03liTLWfDwS77RokK58
GvyBN6xMBqKwrdG7SmKZx1H4ealBko/7UWFqI4ckMH0LfR3KIw+WYB7VKq7v5UHbmhr28ruqwL2C
DGLBqDT2Gy8opyHqzadwZUIfCbXzvCjQyqX4cYK1S6ZLIrmzkDh5q5BJerps4rTZwSwq/Dn7TpQw
mHI6lNvvsRTpMvm7+k+FdwlDRDlC9c3v01NSPXgRi8qBsMd+XQBF8XTTU+8SfwZHwAEg5GndADiP
qYbvRoTL88WkpX5RmfdySRm4lK4qs6TjCstLQcJkvmMCe4J+q/WjlV3JkJ1+m+ANxasQV2qDUNvr
ukzVY1lkeaQOQyG7R4IO3yR+0NL06QFbRqnKbOD/E2oa9O7n1o6VE/WQAInZHnUjlgqiDye5oSq5
gcZobQQRKlkluyWF9WO5jfRw2xOTACWVamrBILOxH57dtpwYGJYu2fGKJFVXC8V9BK2OOAx7F3oG
NKPdWtz8qbDk9+U2+xERnzNiSHE8oElE5y9iwW1QfixSFO/SduP9AmE3Oj8zNb39NN0+sgvC2Yaz
Le/zVWBK9knZbjvLJm6vK8IOEuQAbtVzmSDoZdKYa11DiBCVtlsJiQrbf0nJsgJJOgo5RAO915Gm
GjsJv6STZBXdTp+WGKa1Y2R3V/SJZD+Dsql2CeWAwH7fALsNE+6dOfsrycbsTcIhd3CqvbrAmMxW
jLQ1Ln4O9yGZAc+dM1BjD0QbQ5WNUvY3A3NP/FxHKrKNxRc0AR33wmmoAEh+mScguzr5PsOl9Zl4
yIG6VNPzFVb9dOEx53HIN3csBjpzrvVHgg6u2+5cGy2Vce0nuhQqiiikSpF4HHNT1KwzEJSRXERY
+oN4XsbR/4i9XPnb/hbJaSTgL/yYAGX3FpbUG0Cf0HkkIdFQPMGkEc1kFOinRWbosK5xfsLG3g3U
/uFA1w0NMiiEGdCmsiCj87m6Rx7UXawZT+e9MgHKMyQwrFrc3OF6GmYfrCBJav1FV61HjmiPXRJa
1EgIrWwnr2aoH/WlkfuJfNCcONIYMsmNyhLXRnxjP/1oD9PhaEIXAm3BT0bB1PK0KNKs2IIwEFFd
cHlCFJ3WuPt17F7OnDgougqZSGQwn1XWDwUisonmj+LgmE7ps8Divl4u3gIP1hhgG//RAlxPIG8/
c3zgm4KSKBnGww9q4t+PT9gtw2BZ10sokzIyWA1xlZWaqRTIVIlqWjVzcn/+We/K1crfNz0stKYM
7ElMdKukTYSzMcQ5+SrpkiTGqtbrfoDa4yECYFNU18sDF69H0g4e5gdo4ykEWYZQREy60e2VF1N5
USUEkKN/WXivCqCvYOJUYcklmDsxXfyceIyCrPCrnnp2uYXODDOdU9OmRRTdCswsIFCikZHB9ggw
tRw/9rOxhEQiOk8ghvM0lTOFXSUmL7/h4G4cT1nzE1fguS2cbo86ceLRkkku5roIgeM0HKGWfTha
15Kbcui5a4m9PqXyhN2pBrWsA444GsZFzuDn2G5PLeHe0EZi7r/ssq/uzftiWKP3DQOnfiIMkJ/F
Dx8yUFeU78ZB/A8xsJgJq5jj5sKfRw0P8fpv3R7RwkEXsGLdwdg13gSw0nVASK8mG95G5G/GFM4X
3qggEigQDGvTFBkevqB/k0vCQN+ppsh8lgyeCF6rzmnBpLMJBtawmVC8Wp9EIv4s3a9j3V6xewVk
8VnSLEQqvq96IBoDiyY+ecbfuWxIhhktJywcG93xax9tiFu4wasJYHtwnbKBr576jbN2a9M3xSoI
ECrN9uHm9A55jAbC+Thhf9wlftDCXaEYprKE42yX1GwdQWyGRzog0yqXBf4newketmCfin0Lh5fV
NQlSY+Fh6Xo8CFUZ/vdqPv4UWupDbdcL1fYoBMPkkD1jN9dAvwQf1v0+hIcxqwx93BiMMbLvujh9
1fGMh4lTCT7CjUK5PCKFEI4+tclc9oM7Bfp3R0ZVwuEyN7+iUgLmGNUagx2HUYSVL0KMxy2LHYL4
gipDkjxmP8D+TfbRCe149spE2WPk0f7/u9Q0JKDB++34+e/4wSHJ8J1MGqeGaIbvWi6WsB/7ZyfG
5Ty3pt4uU9HWvEcJliZCHSLSinNZlyDXGgyh9EZXivry9euP1lM/4khgrPsyF8MzJNeAKPXIbFfR
Iup54iqtvhwz0XJmEpvQSN/11sy47jLfnUz7rau0AEJIXw7Djj2RRaZrZEWgJoJHj7G1S9El+Xcv
duqK6zVkskEGjUemGoMa/AjsSr8WX/5AKa4+7Tp74+ayrArswunjyZQiEYKMh1TAUol95EEqnu1K
P41KQc5HPoLtUY6jE0vKjMOQROBF0nBa1D2Chx7viOJ1hR+0ZHLqiY7dQMNLI+i95wgjSyaLNnIj
Aq5zurAvH1w9zCucH+ay2GZKSsY12XQFczSyo/fvoLV9phAQiT36hGHBui17098Crx9dDjwFPmIw
lR7qP9EiemkWCCJzEBpKq7CLP/VZbpL9ub6rcwARmIN/utTDCp330xSTEofwKF8rA7mPzLWr2fPN
IgfJaOtSoRZy2Ej0ClX5uaD7Jr6XCuk/uCzAMiXlvPCPO5nJo+QKZfocZhRjVNcq9sKsnWEQJanS
QfehPnndQ0C2cSLFGIULjqK/3wJhMau8isZDA4vIJ/SoaO3TTeYM3EsvVbcQF0RD+kzoYBbBIL5F
UoU52Q7Jlv/9GOgpqt/PGcv0JlmiXElyga4GFv1/59cFmvtNKsyBJr2tSFHIy4AIXh1M0gWZcDaz
bT6JC1ZMX8c1fw891yaB7Wy6dacJyjQTyGsmrKiAGQR5cD5Ox9mVR1hykprKJb2m/F7uHfHnAMTR
iPDmbYJemK71YrFz9rT1TOC4ATVzC7JeP6pfDkfxMGWTnQxw0c/gA8YTcn3R5T+QEmtnJt0Au5EE
w97tBlGKGzQSfLaQZ4nELjh/9I5E55e3SJc9+9EeBLK0s+6CQTbUy+IhnYTB7bVWirKhdMMdkJET
LRWtDdGScpuPeMXgqcDq5zEYETu4xCaVhZiA/Qtv22P+ZW9af7eI2YmhpqMCJWCt+pFg4ut57wX8
izWPhFacnjtqY7pSeqxdUlhGkAlaeU80x1G2G2z816fsHv1Tzb3rvniV4xABcritD7MvAwoRCunW
ins4b/8g2tXMLU2L/EVV8r2fNRjT7Wov6KDLd2KqoeZm5qM1xLKFwXZwxsDaNek8hcgROZyUYSCC
uVF7Z45NjgIrf9egghbgjrthjItBqg4ioYyh3lrLIbjGSSsD155Bop7AJd0eJ9aE7GcSGWy8q+sW
oBeKX7qOi4gJkcUEqVcNlhQbb92zoqzfZomFPoJALfv+yumqLhrafndK9FczYZc22pPrepFowVyF
zitc727E1287O5EtCDcP4tiNR6+m15TW+q4yWNW4WtxNJavxjfTzzs7RYj+0PWhUFpGm2rJZNItb
zoqicghC4MBXVA/P2lqbEiQBIVGhw7oMtKdUls1VPLPPVhLNBRFEwP9pmJ/m8FEIbmQZhk66cVyj
k7C/0HJU1hw7U7OM4+21HcVXVOWDDz6PWTVMAfeDAR2BI7rq2AJSwyAcXDfX6jLIjUpM/2r38qxf
5JGgymZRYMUzC5nng+zqW+e9j0t8qMj4GOOnM2KR9Vkz3hdchiSxY1/xuy3DK/PLaq3eYnYDw2MY
KtSU0zRUaS5Eit1Hb0eJMqvMRUE573syFDPhMQl3cC0tD4O0jVchiIw5YPNwu8P+wAwH+m/81fxK
YRUkfCHgqJXbRNjRBfK26jOrA7B0jRa9RrduKsKUAhmIp1rBZXPGcLYmTfW7jZTlPYEwyw6kCUWr
CBKiD1F4Y3HTQ6fpkPA98HPZCtyEAr5eeRW1FOVKkoCzQtYh0KBRKiZwR2neokKeYJsXYhGmX4C7
pIuq7XfaiIMVoUM4LrvCfhPPJ+xTl5kzcsVh4Zi8b2IvZrt5WaNnRuSvAVb2WBd6Aofs5bJTClcG
EGr09w+ZDK/fg+a3WE/nMSBplUOvcnphe8etaECeVIrsdbVdQBn0EjTUgwLhnfawG2qix327/qb/
dtjaDvosHlOxi+tJ5iLT0lf3Hrx4uyW/0P3dQQAo3L5KoV2b07+vE/ZpICkt/CtZX5xoFtBOAcl1
ZBd3h8Od/UJd3TFF+MOFYCdLEmjtqiONly9TmhmmDTwObGU2mE3r3M08nbFNwoHyTN8bSpLCyxeR
MxksXIPtgemJonVwUm2h9yoDefW4y0i3YwMR5gWMy6eT6lbeqV9pvoE8as+2L1vqfY8vBcG4/YSG
UdG28WKEYwzBVgzZv4tgiu0e8UulAsaUg8BJjnPcfmF+GcQ88qeHxRKnyoKJ1CIqvWDU/epO3KkG
Xu4Ruc4oqle/8/iQVMEaSc6TtLskdJpmQPeZonRZi+KQgQ8PHARXnjD2ji+KCvnzefFSPNaJckh5
6ZmwLVwHxf4s/+cY0dDbHkorbDbKcjHjw5d6uaTznN6/MinJu+efUWxSg6mUiHQl53jYT5dhAToS
Rwol5zQzz+PUzkp4Q6IfxDgFI4eNrgQdi6cVNLm/ALPWuofYmlfZYzgzCX6jAmW0ZWr7vAcw7Lxk
QwZvNHp51mBbW1vAQruR5pwsRNqzN8K//r8VnufnyPtEZ++Pvr+zB1nsND09I4ar1t1ngKTWk449
Gjf3TunNO+gDuQ6NaN1bV1p3huC8X3yfr9SSMtMtKmcVzjEwx9vzgPssbEBJl88IVS+RrF/78Yrk
tvrq7Hk4yStVaI5PcIIqQ4qVIaO15vOVH8vJfrCFJpw0SZ9NXj9uUhx2DJr7Syygh6PwHJpB3i0n
aCMPIhBJBEYrDoqjHpnhphp0zujqJuJ0prA4z+QAdDABim7+DaipOmbXP5N8Tx/f4DUoBm2an+oa
NeamzAj+MN07JHrNrtgtnuNoiaDLdnG83g8LOdawlCJ59DJ+9m1gAvkGov29L0Ucya4xsy+lPZoS
ZjYUIgAEk54ySZo0WXcQBW/b/fcLdvzyUbwR5wLXhZG4kMMCHQDLtz6u+DGEInmq72jlX9C5jrh5
ES0ZfEoONY7bi0KWzhAVWs+tdcNNcqMcrDQUqVaZTSLoXTw/AHTmmgdsu91MZAZU1C2qrFOqZAUj
4i2Iqv+6FT4wk0EESuUni1Hb4BYSuAz/zETjlZeypaQEErpUQDSEZs0OWdNsqYsxsyrs3GxvfeFp
Gu0GrzNuKSTn98EuHcd1cR1qbMDHkxfgiGvW8vIqucVWhfFxWfE4msMDWUP8iU+w1QDMjVjduBrQ
rwGZb3/RbT/WlsLyFEP+Wykgg8QtWliNjaKwERY3/K9AqV8J92Y7qVVL7C9BRWP8RCoMvix9LuUI
TazjfPUUO5dQTaRsyfkec8jM3E0pkFBOBo5mks4HGxtKNM+a+Odt9Qln+x8WUeOlj/aJCVGVJu4X
Hi4pEcuY3vp62yCfvechZ/lTKjgVBFEelbtWMFX2LfFrGDKRozhqNC9FmE6zyvVv3BI5UGouY148
cCg7qJ2sOsn1+84MZZlIjrqXj3Y4x3nGER7kYpoYRn2UwcwQnrFqBl3NDs3Tb7nFPA07GU4L0Bul
mabQHYcW5dYwE8vG0h20oN4vvvOABGk6QZigTyI5hUxn6f7+6LG++4k64ndW65JKK0PbdlJaT1PK
D0+vF/eqRADnKER+CppEtAorPf+oz8yFEs66vxLZmntbapMMsHkE3dHUnR7hcaGfofGi2iJkl2oH
4hCb2RHVQPRvik4qRkXBSXdaf7XqDTrNmdGrhoGOlO9fgbMVgi2c7bKxsiu3mH6kIAvRHhUQPj8K
javdzT8GYk7Ntj3kTtyQqOyDITn1EVRmKNl5GO5KqZDTSbcK8wIqb9REdHJqLMFYRpYb4FaYsUnw
kFsGE+p4PCmqewTbe5OK/JpK+ZzmuA/hAwYN7dmODjt8kco7AZ9QokLWI+XkiespZKbixt8S4hm6
1kySCq1vJKs/sPbVJk92nBGvIAYCs+fB/22CjfBG7dJeW7vKuWbx67i7l4Gt+8LxuLFij7LJUuHp
RSgur5RSi4E05PsupmFQOaji9+9vm3NLOy1IVJqDX7D5oY+MiPvFqeQ+YLHRQr7FdbsAGMjt0y7E
VU3hwPT9Eq5GUJc8i9jPGhz8sJ9WjRUZFCXCI+0u9qvEScohe/QagaNV89RhVRLNLfvtG0FLR5gK
whFs66MSuKHeRnHyXINnUlDM7R1j6CdSfiDw0i4JBDee6/bXWUjIzpsA0py4Wyo63Md/aSvM/XMU
V7Nnj13bzjThVPGuguGBQX1MRbLy1JD9+IWzicLo9+b2AqqWQ13mtH0qPE7BhI3PkTKy7DZ6hw9/
vQzBpg/Fe93SAlbd9LD81I3tB61gqpgU/1gUGsyb8WoproNQ2qAbH1ih3PST+MWVkIABJu3vnFbO
Y3l4hWzPlAv5h4e+SYAAk0bPSchqJ/mQT0lf2doiQbSqOi/cVpiuwYLW+uwS2d0qpOqaJX7ICcGf
Ybz5XBkSNi2tYwM+d4dDsO6FSbWvqy1S0ZTHvRcXfDI6lpYvXhNK3Y59Uy4xkeKQyVgiaFyYeJiN
dzpqy0QeoLSyoyKYoUUVA/fKwxPOr87HDbvjDFTnoZmK6+VHFcLvWc3QU4yEjiu8JHOSeQltL1is
STrBR1wpZu1P2qQMqzIpLbT5MZHNHhKlo5DUap1Ug6+x4sFxq71NCrzj32BWdj52O+vOXg4obF0k
kuxsUMmhfpO/FqgcD9JmTEG7kTIrH1GyovEPBB9z9vFhSg/m6xeVG8qv+tmZqsjJtA4ShYm/ad7C
YN6bqAmOqgntJRJqgEnThU1FnVQp0LrcCMknTzQemzaOwXlCFlBiBSnmvtdu5spjYNwGLd9ALmqj
P5Dpm66pa0zA6n8abq/PUxBx5pmKHE6hwKYnkDPnHCSusTIEuw8SgrMaw6u1UFrC2z31OeRX82ke
rKsQJnFt8ZgvVoXbXwATSLgt76tRbMr2NbCCl8kqclhbhMmNzoe+5xoedDvUnDrcBgytNeW+YgQK
OLm9LYQ1quWEHHg4IoTn3nmjE5L6tLDtoKCslTIB++Y6dH0EvmmePS8LAuBQ0E1w5fjjDCtWi4uq
Utt1KhPV89fnKK+F1TO7NgP5VwUZGwJibyqBsodJD9HOp7VcjoK+0nE9RA3nv/ROu1BF0o1kz/6H
5ev8gizl3+eZteY0TUblcRU1qjMIJVAXKC6UPAQKwKFWrNEqz11nMiHLA5VaPlvE0nDP7L/oeTDB
qF7vnO8xV5KwFIzhwPtLiT5ljoptwjrK1YPXiVL7JnlG68M4NcbVUnQIWqam+xc7jk2FYMQbN3ze
h7S3DDFAJtaZpBQ9ofVwrI7QbNOZoMMdp4YB/qL6pDwtIjG+guE1T9aOMfhuH/Gcm8xf2wlK6i8/
kyTrl/BorM/QRBSaB/rfeD8nu2h3EEq4Lz1f2Ym/MihQilXtJrh80Fpf0+DPtVty/kUTaoVZwhTZ
B1jRNtFo3oHmfvqRaTnb3SSTy0JohThOZMYyp0I/Bm2Use2dtgz12nS3AsgIQn5J+DqRKy3Qm2wQ
aFY5eLwhrG4/jIlhLIAwlDYLzXCM70ansTTfF/cs/xW038l/oN6uRehcfMLptZKfvFqcsWJ4LarV
915S/2x1zFuRcqfawvlvvR0SHu1Q5VI0ATbNGCYQAqPTFP7JQdqgGMSBrtH+Tn19BVX38MHxFQ2f
aSRZdM+dH4j11FrXvBSsHVMFbn1zmHfYPUZ9yXouodP+tmc5BRs/AnIzUbuGNbU/oYknx8/gI3RG
PBw2WskDDrCvA14+jEXiMhb359B4LvVFqVvyJUJRv6M+HfLaP0S76CmcPui8pqAkktpWb2UzMloN
cUqI6u+bHWE6fUh1t7+PATR4wKGY+caYGykoQzSaGqJhoDRLQgehH6jqPhhz31cvpw9cZS+3LRrc
w+rzX/W8nVdL8VNDlPcXQrk3EoOti6NEXw4tRAgVk/MdRREA4j+/KQ9iF/BMqI/wD8E9MgkIsHFG
0ENv0vr0ztW3MszN9DljpMBmAsLWgEEmoAN7pq78g3k/40nscdjviNIe9lZqKJauDxbb/O+FMG5Y
e8/xnID9GbcbqSjaBYu0sh/kmViQUUalv2tZVdm3HsWQnLQ7Rc5Ju3bcWC/AuBTPH5Iil6bAUFul
1l71DmAaerflL1QBi4zzF17CgKCuuqwZtJycSq1Yig4XAlGpC/3AsJPHcQXUEb1KxY2wCdF0Klex
l+/6nJzpCI3TDMklEAUo8uKPWnhJlWqa0VvDSjUcz2AABdESioCiyPC/qu3vf4ecpeCbUM+aLuVv
2tZiZmVrfE5zW/19MrpHpnDqARdUsHTH9/DiU8VdSsG+aa3WufS/KCOqZ570sZ6R0+1ZsvlJM7Py
JA1DJW2JxKfCqv2rmIWMRjnQCfAgKLBznxZv5KM6vfXrCEphoKIGkEFrZ0WvcuxtR7o8dqHl9tkx
paYLGYNzSud4K8Xt3FdxnPSIv3h2ie697eV+UU/i1xxvLcyigyX4zESaRPdDrIazHUYt28v1h71M
nFxiymwY/t8De/zZXflFAFeJ3PB0EUANI2JiUg6sBcYJLk7iSP/kcJCowqT9lH7eCOMzRLMhqtSu
qQ416xmrZpKI+ti71jUyVefx64K06q0TG/WtpA0BR0ZRQ3L1u8oJn2FZzpMvw8s136IRQM6x/hyl
KbjNnRyLiTrpcFeNV+9TbZSDvnQRGHSbQg6YTdv3gEbWeP2X/xYmwelX1U/nkbjrEajHkIiUPcq0
bfqOjDSvS7CTusKsKtHzReFhAjavpU3jObeN8N0zot3x9YCnF6BRG9FshQ/xlQBTITg2UbB2Cytn
2cznP/zamg9TVaEe+Li/cGOCmA9k3MpTGF2yIz+rC9IT9O6yHj9ZzTbzsu7CxRGgbQ9NTmjSeh15
V4rWj/nJpjSkaQNDoNnwch4mYoreEM5IODrS2FCqrYATYiBXaQiXVdupVcIpqKHrl7YQSGge6CHO
k8dccFCN4vAMIAQGu2jzbY+HzPw5qp5sBoJyLAnsWW337I75VWdlKLHO19Z9Ntr9KhUXmA5X1794
80AvXyBqFlbJazy0EKX5cGNrCzXmHCApdNKpgib1sMWH1ufzlJNte+cxZYhNNr5ra6F6ww+RKjDt
ecP5Vy9qGv0Kdqiw3Yp7i/kHklfqONLZkSSrz4KnicaDugrlFhzVw9+ZiUvpNF2SyTTCiEXGXaOf
KmcdRXMyuj+dM725xSxd8xI5QyqM3t28FVCRRLrc6CmRhhhS4j8/IKyyVuuuJcs1SxJnvx3DJuw9
XbPOYiQTyc9CHlMw6oOT8LTRF0WOF8SEmv9/IyQJ1Y6DOAMIQXmLe7nDpHrfs9yjkC7xHbgnokfD
fkkrMi0h4BHfPHywmWhDaWD6neNNEA/4tzpsWKe3i0uOXhs4w0Clg4U3fOgdCmKm89ygs1JGmenW
gHSnc29uKk2T9YylV9FJcFW209N/WAGhGMJrO/mNPg9DaVJ2gkEwWoGma1v3oBYsIHoEEMgTl0vs
Ag3tHJpFbrgg2RwqhpWzf61Cp2IpsFKACFFh60kPTqFhnFp3ibZzJNmSYzFWJbg2aoWzG0SLMitv
/czxrRWi36KektHBnMTUBKvKIRg3O++MGdhZJ4zd5Aokir4SKFyx44MgE/hlFeswZX4/srW5C2MV
jG9W1oajL82vKJbgWgbR2yJS9UgP0wMFk7tfVfB+v+D66/kwCz8Lg5Lbviu/BjIhW9QXqrS3DTT/
D6hJHyvU4XCNzBaIJGfGimbG4uu4RS4jmRlkjn0cPnwZAtDz0DzsEETEeqask0iWPvQUpzmc6Ixi
bT1AtiFQfTwgAeZWptW+wjvstryXSiSExKZyR5eF+bIJqqg8BnpWNF9q1Rf3GyGmJzyeAE2DDXWE
Eg+Y+QRjf5KAbiOH+9U7Vnu8XPAF8BjrVLP8m+BPz+94MLRGra+iD4Qb9soQYYkMWEpHucLHm7dJ
r+TQ1KXBsOH1viq6WaJzVnZxVA2xMQ7XAMN/uH6szn3NMkJ3tYKmEkRRVMKKg+YAauRYYvvNPMGX
Ij7FSQCmWbphLJXNlGikg6Rl4qYp+iqH31OqWzzzazOAN0s6mvDN7WiwQse55TzELR85jJqtZfGI
XgKH7yFZ2aonsUQzR0clQOLVB0UWEXroan8e9zHC4WPTp589UTt9rCfgwFMzRz2D8y7RetO/uuHf
/mhAin7WREfcTSSkLxctZBe5dtcEYVIRf7LIvMqt541X2C4vumOZlK6EwKVftiYv3xZqZLouWcoX
Zri/bshvIsWenc9UUsYP+K9IfbHM3R1CJNn7B59LbL0huyhm0OXOzQ1QYPdHByb6qyJpXwk+FfWt
/yjUW56DS424Hw74Q3jIv1Ki3hFDXYBORUdsvq57vb9C6m7yGif4jTN/iwNNddguevdT9ImCO9w1
unTHKaxuDi6IX1dFWcGRB3WbpQeu1yr+0C6LKWnVICxiVXH8h7vidarxjMgmtnR8Wh1NAjCmiZ8A
CyNIXV13OaWFVb1m4EqHX+j4R77gPz6KDXOSxCz+82QVWb7+Rv04Q491HjjrxbTOnMPHWfc8GKbV
ex3U/rUWFFhyLa+B9w8xhOHLFzke1lUnK58R+Pc8jvKN7JxvrQpkPNLRGiIq0xJKAsCttnQcTWwH
eycxquuE9DOgoEu+OfNOVR5RXFUD+7/ugwty1MHbkgkPYO4dksv1WbXHReE8PGvdEUzRt2i+6/NN
GCDO8Z+z+6SJBQc2wHcfGqhqNLuLSVhFBC1NR3K+nmv9NAZbdlEkrc0xIwk854qdHfa/q/7dLluC
UQZVHVkZpy0kPDQq3HnuRDHPcRhd2GBs58+ee8VN/uSS/IRDjEwT2lIAziToIX5Bu2Q5kjYxvhFD
YcVU0ExRipMHU2Vx8eR5Iwt2m8AkaR+U69zi1kuu/qN1Csl/CuaMo9TfCgscL644/GwAzHN30nMk
YTdfyrDy+V9FI397tslTWBBKk1UW71gKVHxDhA2nQZ82o4GRJ7UvTOW7fNobxC6EtWT/KWgvwdae
EEzB798AJ/IQocTapP4KR/E8PmfZIzrKk11Pr6VnPC9DqoGNjSTlgwstRXF9i5OtT8S8i5FjWjjs
ek4hXVY5BRxe7wNDwmnyx6cvmOJRF78BIELTne+FOaKK0k9EE/16uLFzzAjZ3KY+FBkw5cR2onnE
rKn7smfDb8QzRjYUG6jatwH0RJeIrw8GhWK5zjC3hNqSHotahXxrtOfkMpwjqHOI3oPD05tdZJlY
1vV86gOcWAr8VenlTvN+5vyp1w0+t6mj6W4aObxe9tqG6eNyDtk7Do3fu4bcylSZyTjg9ZxzXHm/
Sy4jdFHviq5CiNxk2GzS7iIxwiDeM0/zMqhQcP6eQW3XbfFrQPZrGJZH2iR3S8cxbin1qOszbeHe
0GaxAg/Eaqt2w23syKzyWcJwoiRro7eLz1UKoYK/PnDtIctYhojuGBccYyLSHx3bfP5Z+ETDt5LG
TBSDWqKTfls9W6VIcxY58TuXC1rZajqldnNfQO2sHw2wavX689Q2X1S7EtVPdvgY8/2cTOtNa2rw
LGk0vM/N+d/ATDKAYD1oKwgu8By5dczvUGxIVwtSZFgFxt+oXhnBe95H5jhBWZJTv4wcw237kWuV
LGevJmMPW9l4x0FgytcSavZA4vYkCzc1XQuVfEjm971/O2Mq9bULkcIpDNFS0jhnSQJGHTWAbM+D
sPh1PxzPqX7pfHfvTV1RKisx+9/opAMAzPuQ8nqu66hCki6m0zc+949DPbIYUFhEMqaO/hNuG6BR
Dk5s2Zpujmq7tLbpSCUogK8BqnPSa1ObxnvdV+Sojr3Z1k1HmbDsT8yIrEszWDbeTI+D1n7dauSL
EafO4l0PX14hm2vYEsh9s/C8iaLMptiO5RCyvEW3RxOJ92qieA/lk1ZDfPcsHumkRbxZyuRdcSmH
qnScRaxmtUml2I5BHmrIMW2iwdW0OsMCZ5J6uuAv9916Gau5UxAunImc2qsKjHbqLz7/lugFiUsy
HBpnIDJrdf008RSf5pL08zMKicU/Zv+ec/W87mfxTV40RxK8S+pg2pB7GCNMK/DcID1Vn5jOzEtp
K2a6SOtpvpN3hTci22YviJY3wIYxn9UC+XralMKaqg8sXgKLvrOBqh++v7J0yCIhOQ/rggXunI9Q
16OhroWlORU/ooT4UDR0i0Q+tWV0a4R6udVMJ6hgpzM2tThtLT4KvKNoVLvR5nSYYS3bOlnJ6H3m
agSGjem4y8BcE89C6YFiSpX6En9RQxKIUSvFOi64bgm3xnmqU9TVDX7g/7sQZhiXQAdtAA2CksYG
m6FXzR+EtwaBu+x0RF6+2hikkawme8hOO9zXQughMcmS/OLLpcZCID3f5X3MTellRrcfrmEDut/S
sL2Uk1iKyY8y7vUC9eFisVLEu9JVlF4IQA2Apb1sEa8Q3Jq7gSiBFfCLpy3CN4bArMFfc6ckuoIV
c6abEvQBQCDsoDrFlnp1hG2BI8RuUqcqtaqz+XSuWTi4HZZH1OVPviDBhnnkZGq0RLX6mM7sc00w
EWIyMfgLDRITjIXEA1f2EBD6rAfRUaAk4jPdP8imSLnpMocVXJvTrnHsxJchqQmcnq7hFiy5xpbL
6UZc2xan8/O4sesustKlQFXeX1glN5ZNH0F7nlwLYodrUcp2Rr4ZOSe81y4XzBtaizK8NZ3qLKMX
L1gRPYbCmdv1GLInB3pt0y5jC3Na1BD7PtOLIJq/UZzvPsnpcgc+KCmrwm6b9IUPknS1lLHEtMSb
Y1D2NzR1iJHCvsCGr/5PSnORN8i1LiRI39duAmYAexTsn1Oy4/5mPDALW2LELIU+1PNl2a83dq9r
ZpWt7l6a9wpbxU214qze1LSVzt72AgVWgwGMkIM1+4/BUUI3YdIj5yGKac5VJlCPvBuQFX90AJos
ySlDnMkQfWpWbMi6Hb9VCUqEXLvaP/qKeuYng1zfoK8e3iQnpW96SRYNeOLH2wXEGcKRBEnbfhEJ
GLtVFxKSkGDxfN6YrVP4BK/17Y8LN4W8aHhBn5LaeQfEv+UvCRuW+uXjgtsjEVWtJypyI36aCaa8
Oi6tD6LjdnYA58Mf+z+X46yK9g0jgVKIi/jkEZ05pvrMxYzbHg/zga987n5wrLiPK3ZIqMsJ7qLD
JoD806FDAaH9iq0nktUxv2XlXuBKALnQQZZmkML2zZ6I4QTnPGV+QTsH8l3zwJZMMl4zJmmxQojg
uwE6cWQ/KpmUtns+4CbsNW4WLNh0gbWiqXoWPVsHQfTB7MANpdpu94pI5vuC2lfv685gKRqk1zo/
SfyH/yzIpm+8uYY3nRZM0TIGisH8es9ZXVZcyzndcfABlnAi8iTw2HO9CYPHl2oHhaIztWeJFSjl
fNxXrMtU8VcxmayISqMiW1XtPTg4g1LSLw5PtwR4uwvRdbiLXGUJAUKpdgs8Vacd1wmzSw90kXgL
+DXrBA6Ki/0lRnWo7vTP5LwLBaLXEtFVsS70zUcQQ/BZVB8yQPVzjSP0Gy2O7/LDkVdif1EcGVj5
eiTKTo/tVj+nM39fHkfBxlad4oGkt4zmz7/ZaVxSndsvWR/JFcS9udFAD7QwBHJLfPTQCPGxh5kv
YQcNAYuAo1UxlC/uyCewS7JtsVscQtEDmvrFoIWbqj6YzhhuqPqUsGF/pda5j4FvysS2rCoiX/JK
fyn7/VJ1nIPZfInC4xYszsC9wFyDf1ajYoGNpBwj33HIxfGK2ridY41xbAj2FVk7+JQVoube1G8k
iXXlzaCWpPKuDm5qjDUxGJbN42UXG+arydJYr/KxJ4ZkpFelsI/cnX6rQwNMvS5gYcX9oVTJj51h
cTPwPnUzJK63WcBGC72OkOowOLMmMaFcLoYiEOMdpowV3eZ50nn7gKXLsdnrhYsotrHhVSdZBthT
9Jp4CU/VQeLKr+DCt/IFoH/zIWv8Yi1PlDsagZggjneFjlmUq5qIefx/atICVI4W7vCKZylnIjNU
0HRPOwoZkAKfbBXMWwWiIJQDnvEYIjod2XyOAfoQrqbEP7K8D/jDo8SwqTEb/g5pi89M1QFva2mB
DUVBcnN3bApkdGjcSmH2r4FkySlGgqnHSjm+RxU+xj9YnT4fju5DNB9pZ8XeYaGfChz5c7sSPoFr
cd5DCGk50lT6dZ4sQjRJK8dPCsmU6cIZC7WwCpWohrQ/R8uMtDk+m+NK/IT1rm3Q8QZvRvncyoAz
07GmIzaeaU06ZRdy41R3gvkI/7OAxKQQllf7CG1TD/obn4a9ct+b0s8HyuHm8+uMNTfJVsopWYhE
c5NkYUCLnWc/9DDGIa+yl7aH5PSlZAm7aT9JqX31R+N++g/60BMZQTozzE9PUcjIaOkE8BszYsfA
mm5uNZ3S4xJ6WsJx02PmPE0ozNtGyEc+8Ae5Cq8ueV4GU9KdgetJoJWbWwxkg49ph2+IBs2yhjwO
4fXYH/xdTwKWcoSJHr6bTTixIoeoKYz0CdcnSzruTVoyB6Qbilpjk54U5SzU51YQv6Y5a5Gi/lQ2
vgY/lVqg9wEW9ktdWvsByMlEIEMtKZLkBl8PUPkcrBNW7MXNcbIuH1sIzCQ+z928JsCInNijEf8U
b53FtwyDhGFvjMJ9Ufj/I59+e4ymyE0OLQurisSgwk86RScCrLT9evmeK1zN6UE4l0wuYuL99YpG
Rzmn0Kd4V7ug62oUUPqoVWQ90xJt/FV0+dVi7ScmRr4qKTkkegXvicrgJaDJ6zayy+2DY5R5g14X
4eFVoyNghYjpvICAZUa1B+Z0cLqBDhuPvUojZgfX2YRITLkUuGg7bawKiKNoegZzsApsr8WfSduY
Qpm1939T3RaQ/LFMWEB12QsmKz1OT8uhub4HvhSFkBzODgCK8a/VGOUn0LDZ03DnC0H2uQBnxIjP
5Q1qh9JqFUlfb7WiZoKS+kO5XhOAfEHEYn7MmpfN7uFXepe1mouWQWqoU1xQY76yRoZW0uWaUE9d
ejq2mdRhdbXZCVgLQKWkAPcMdQlPwZTgAH2IMWVFuS7aG77702ISJk27UwC3LA/7I3LMf5bud1r1
FTQq8yWnRr4nkJOJgVQJCXy3ccYYaOHXZzizvB07yD8nkfV56BTtSmfKBozsE9GB4La+vk7yO0tt
ky5AJt6OI3eHMFLFNOV7yR9NhqcQcVbQVlx3naTN4ji9Og2MBQcQQuS5+I8X2pMsQalOr6hEIw9y
U6I1UUO46Zm2FotydoMS9h0nFW0Tdp74NeAnSPKcnZypkCVbosqIIa6U7niM7G+UjqvskuG5EWY9
lfW82d52Gwq89T/CI7PJsT1RNsByzrveuXaPj1QxOt1/yfv5FZ2fqte3rDCsrgK+wVXjN+YyB/Xm
PUVNKN1WLIP+pgJ2MnqqAYbwkxTm6dloHxfOHYmk8EFnwbsnB/2w0bM3PNhWJOlBXmrMA5MRXVXZ
btEo1TATYBmWNhmJwUPnvyGfwiVUBAKnv7VyyKj9/L5NgrKto1uKZtvwVvtMSjiEIi2ttkj7S4Gx
KyVWM4Q9/3KKOdAMybqvg/yGGZZVyobZhomzIlIrD/7IuAI+9vMXuXaxeEMthD08noHhA0QLjpjC
0CST+pw91V7IvYXHF9s6/oLFvhMYbA13XN2mPphpweyxyQmLR50xPCNqgLZCFsR8+VywOMUA4ecv
eT6LysXqyhLrIhjZN5nwXN2AqLq9Jy71Ph3lfetqlv52DMAo/JxZ163RikPa/XTCZy4lor3G81DA
Iydamn/LVMplIMZ1U3lH/c7BY4uQ3xRFbJYuJ6UAxXGF8p0hirdV2VMPoVseX91cfEAaa3OUL3g9
AWJYmkcAeR+zKcDtZnpIIhjAVJ2Z0T3JKC8LvO5cO0CVILoB5his1nXgLYId1IN9fi0ANrziT7r5
yBbeUUC6pH1cUIL2o3SAkfdFadhuuLJbiRYdzAnuQVWczi/v+QpCv9PZ1YdkQxhPICNEZ7R0LBUS
r++XhpYIzqxpnksf7swt8n/V88dP+2FE6ak0/1uavQqNu6jDtlqB+fvrDN8C0kXb8WoFrmcUfEnI
f3AF7OF9TEZt8Tc7xo/1YhuAH3+sD976dBWmnvYMOyBMbSjFIPl6Bx5za9xUYElzr9PdA+En3LBQ
rnjqiUb5uidzv1ovp8to12KsTBbl+ScgX8hiHiOz3+vM0RhU+HEuj0g3aEZBJsO+OmlKgokMkT/Z
6TUkIcfrBCp39isSH8YsrL1joEHSp2kcrLICl2YObb9iUTBD7BKHwRyoFIe6S4+ESatWoIq5QuOP
02PV2XYq2zKBq58cOZR6BSc2YIG+TAeiGrhkVQ7LFC6lU2Vhp2+rfS4xcHs8IDbkcA9DBx5INTSt
jcB1pRcLXgOWfouIWoIBp+M6A9J2eSJvGB2pYV37ddaEQ/iWpux33Q+zpIygty/6JG0ItBGPNGXy
hDs86+VfGVkVnVwc3gp5zJqIT3rJhn4OUWiduZKvEGqRDL36gGgbuLsEP4bHAg44X05KK1muWT0V
wpHH/f26HEh4HRq3NaOTZGXIExXUFHYzhbvWe/WFr9+eD8TjLFF2HLSTp7C3F6wGGbgKuYRBzuR7
s84OZs/TXQQ5q1fOWN2E9VJlMIADVHlig4lXYmdG1Jb+Wjon1N/7rIv1lUQQr1d1mFVudyeHpjD+
SGgYupyNfCQsqeyecSLeAeflteUDZJ6hjSKw4xGXQBn4f/26wu7cJmd21hc1nVt9NVjN9iIvqVQ7
f+qeCA4jzai4uysaEonixz5W8IvMdgNQsmT4+YawdStDSjaoH+OM0vceg/IO3zIR1yq+SR/j+Ely
fpjohIDzCbhcewVYsC0EIyvHrY2NPeqc+aX+ylhrtBXbM1jhZzSmGr1OhcNlZfoi+FuxHQ5YP4Ly
ncHWEC5tmL3bpYvy9WRr03W0IvXqM39QEkILqLxBN5ZelN4ei8Fsshq2RpT4GF8wZJxHhLYbBmJu
i1gA7LWB+KMDpZ3bhIuURvlQx/8dW5VBc8P98DZvVXHLaKP0yOgY6F3lAquIXiRn7TeUjed7zBjf
6C+qEVgTwjZDFfxHChrlFir4RbRJp3Jgaj5mKuAzBPSdE0k18pc44f+dtiDlNhfCj8eN+qps6PM4
Lt9jbBgLIVrLjElwBUUgzLiyKvSERId8+DuXqmXbJ1JCFGI6yvTBOuFhnNcWWGhcNTdicMEdrPc3
PC06DQUOUQKkWauIBosWIM03OR6vuxsfF5n1fC5hjsZt/F/1l+t/DR3h+2/crMPeyMHTPLf9ant/
x+s+KVPcKvVYF9Gi2DONo42Ha+AWc489L3xiSlmwD5mVBOMUV4NfudS/wQ5ix1BDVt6Gmm+ggFDu
6ql2i+ebIrs0PpPQHL6IZLCtO7Q8m2N8Li3QU35kpVNUwRr8NezuLzS0+Z/qSAD9Fr5y3nY6eTTn
2Rzqs73im30on+1gGRhEnGVt7oIp+N/P1/+NrB2LIpGq5LjHsY84kQCzLWKSm4QO70mvjnMUpZWn
nXBruVgkeHtBEzsJWfXJ0hQtA7JqEZdVuVXQgEyh2mVnTRX5JN1+cJmg7N8AAMxsuHe7pyfDyaUl
mPFDTnEaaf+Zmdn+Qs5gFXX1TCV/vWre+OVSRCVJNysDzDlh8Cv8LUq6u8ijYigmUuEK/c02dzj/
BuON5AgXhgJNeBt6iyKhBL2vou5LkrUF4ZZ8D9h3mOIuoiv8vUFJcALnypVkpvP5xN5ECevNr3Ma
oniegkg0ewULjOLUAz9b0dFadDNPEQSwNw+cE6Do6Y6SO0cJ5z0m0ejBkuesXHmLBBDBzMMfj9OT
LSTGhC+Hn0mtsqPFXdH1g7bWJui7rHM8Lr2gI+bTYn4XmGQmwZre+w2D0PVVi4Oh2ORDDlK1ZXqn
WlMzabCAEqQnv8syLMieAy5UPZO3yML3Yrd4zLJEyMGHBztDys3f3ayHNWhQpld5Wqf+gdPmZCEe
LUeUVgY/wa5/ZvPUVHAoxtdoup0GmtaEYx787Ps/ZNwgk6YHgexzlRMrR7KLPGcyQXgtcNKAS3DM
cbs7U/xc8tAb44KjF8C36HjJ374VHglDNdJC4T9GnfP6FSVXYuyBzSi0eSh8srNbbTygkQXzHvLO
DgfgzWLSQ1bCy0xYLyHmPuvH4ipHhEuz2LHKpaaXD4CtgCJTjZQMf/5WWPuHIbr9AtL+YrdHnVn+
dgGLMo3REkqKOklfhm0ClbmiqToKko/DDZoQ3Ay0WZmoYT3r/PYKi1BkhixLFa+dgpNtF6meh0bU
cDdACHwD7nE1XA+eKEb0Lyp8B4mrU69JU7vAz3t8yLEUcvj93A6R82Fv5RD74JLLZsV8DcTyF5z6
idZ4sRCOdhB2dTiKcQ4dwDdrNazgW0mu3mULGbxQG/+UKxgWQ+HOTY7KLWR7ZOn/U8iFqUFMUflW
f7xGta0TUSHTVypsLRaGh5SEbbw0uFkWb5HoDmzGqoVSEEy3IYHa1wbvB44t7gW1zTArT0jgJJnR
7Qx9E1WMTuG+QMgIOITMVta2EMINU8HJnVdtnc16Q4W8u8KxlKvvyQ6ebWe65WMDsHZX63BG+CLo
zKYbI734bVhHcOIUhGikqCawDSaMiDKOvdz6LYwhiCcmsZHoC/vYHlZ6WCLUtzkvIFmxJn/igrhx
oQrE9O6/WG0YbfiGFta3ebzknkuv+CrmB4K3jAhzRUelXjJleny+771AMDV5U+Hsn6ZrUYizc6An
SimiybhknLTgQSYx0WaDUvIJBc6RC50blJ5Y6qseV446UX7ghQJVWr9eR7EogfdoxZeP4WyDd8mo
mm7cUtaEiRDR2NFJFAP0C4nvwg7nZ51BZtISIY5HZnaHn9P9mJ66ljA0Wzwqf3nNlh6OlwUOGubO
W03XLtiyFDExIzKQ4RmV9CERkkFLRzdi+6YPCJoHc+NeLMuAzzwQftrampq3mPSMaOZwI8ZbkH85
AfMkOl9Hg8OznDPr8tiGXAo9I72W7IYY8s9o10TFjdvlDQfYZOquvvteClNzEDaSR6pKFN4Lmorc
xcuuWBC03ic4M/tKghvd8aB0xv0iR0arrRBGIFK4Dj11Zu1+yuqy5r8JLd+LT+PyH01sWlEI8Q4B
LLD1co8PpNhjmbPy+kfZrZwyCAmWlncGCu5Ufpad5egF9GoqzpceqvsZ0e1CTKkmCldon6ao+mRA
RCQpTubhUHYdHgFwVUOQR5TG8VCNe30mS2qprh/4PziaQvi8s27KmrDSwUf5VzMHrGQQx7qzZbLH
g0FlpLw3gKAOCySX4ukbA3+X6rMf6Ht/nqqAZi6QJH4cc1TYimDAuCBztGNdcZQsZ2p+kJcATVlk
WfLR5KWBqhhLK/c9U9ZMNznh0ioCO0is1VQvkmUoYTMKqzpzrRhWmutZ31RFfmxWk9rWGxbP5rj4
t9wzEHEGbhXxIA1CHkpmPauRCb1n70atJl2Nts42L0tSVP5R7RmTWS9iAH+C3s5mPhjL/8yIBUdm
CkbNt5Ecvj4eqs1i2BOrs9DyQtdtpac8wE30h0ru7Cg7qqasMkf4rUEgP1X+Wjua3Q6cpIZWGHzJ
p15swyZsc1KINAUNX1V5JXG/cgp+8gv4SsdDC5lwGEgZEgNv+LZpbbAGdFW54n43owO0jQHHVK7T
AWqPfD1h1lMNkMqyOO0pLsKDYwZsi+SSc7UCeeXLcZx0rbVJPr/67WXeaJje837Jc61IBfwAalzM
L/eQx+cSLWFolApGYllAaxmzJi/6b1GmSweBTC3y9o8Ubk1Ak8S7vF23ZHGtErnItamzH8gINFOs
GBzdwTbhgk9794OPGa3k2brkLBdF5FeiTyzXcHhiXV038OeWy+4iOFTsGmw5GNLuIqexLEJgavwn
g3kkWdJkiP1a3XQS+gAVkjAGX+4JGzS6fs3u0HPUtfcCvPja5xTvLABursXQ+7Ws0gPxFuvgoQCu
D8PZGPcEFf5ij5nEiUk5z3zUWdgd7faOmCKp2nAwB2DJ/7T40BTwtqJgP4q+mLuHgn02U+zTsSCz
gV41G6oCJMm7Kvdrk43cfaZt5rZnwRHnmpuyyl9FcuK2jDX9/4JL3eBf26LdExjvBtVZsn5XO3mK
Tmf6UwmNwBMi/Fu8t/htaBidNr0lZZgPui+9OFluSKOGyX+nxWnEo2T0dL85VbyUqNDvBvx7VIxU
KwPGmpSxIlJ/TD/EDnVCgIXkNDb3yH97Yq/F54SXAPNUDTRybc1UfCHXjR0br55FdL1AviIALz91
6iHQDQP/1nENDKzqfbOXWRF/e+018XXVlW2wkw+I6NX7p+7GtKcMZDxY9+InJ7Dzxhgp3F5IrZxU
Rn8+nm0DiqpTUKds0MpZ81/ZrSO8HQCZampecW+DOTa3q9J4LWnsRmI8VbiYoYPPCUvEt4E6Zv1F
e4hJ5jaHUbukmS1rgyK8+nLHA8ndTWAhupsxX+EwyYrZFmJp0W7Bs5MuE7mGkcZ+v13NucV7wkc5
K9XYXgVs98D6aPimwft/8E9c/3q468rpa3eyCcswlQysbkthyz7Xr7JpMupfhhKgF2bhLBwczg2H
3PY8JiQ51HZqjUl/9HqP78+bg7d/YZyxh0xUYIhRJFggeXiZs/eMdUsKlzTcLIsHLSw/fA7SilNn
DPQwZtnVBBcLeoi7O/NlspfI4JFTDiW5OogOXm/gTYBVyUCRaXe/EzPrSqCci6fLT4XQLvwA6IEF
6KberLZ+S8i+BpWcmU7stB8/+59zvgRQpeYdHvJf+Rzlxi8E9s0sh84NAe9BLSkGkHXTzRHLeFKP
pGzq7TFBLP5KeQqeA/aoccp/cVwIgpNqMiDS0VOL8rWRLmvgmRhQJ9NMAxEfXz0ReUhJbURtPTil
1ez6sdVpxwqgxsEcXw16aWVV3nKMjQIL5vLksYk+os2pCeV5q2Rswr22m/OqhkCxVB69D8h3SWJH
A3Yl+O4MS+jFE4yWkVAfeeGDZqAYz17hqhr+hHqrFC71S8XvN0Z/whBY4gfvQ9JFja1/eN/9XBZp
UiT31gDzMg7FCnfq15AfeyPoHOwWJTIdFvbEqC9FZi9SPzOQqYpolG3M7fJyATplldjoQA68JJQg
CvxVRcBShomQT6P5346Nz1aekPkCANjoLDQFyWiQF+cSKZGz5HXrFfDC7LWIzgw0LzyyQ+UD2X/k
CZNjlUp/1zVv6qOTOgWGrrC8Q/tpF4cyYe2JVYAlaqmGpwCrAFmZ42ODx0nX9GHlfxB9epHXPow0
8bKD38n3LGm4EqmAdhqj7trJ72ZsJ6Pe7wZX2JpuvBWFXrwjgq/QNhCr1RO237YyXDphdFz85fA+
EGuSOY+/Lyiaa2rCrC08ZOL94yVF7Kz0oDMbSZlLfABNeOxHLtc7VjSja49mGl36xn8Dd76kUJkH
asngw57kgSvGIYkSDgaKu//Skj4TXT4yc49mAncBX7AUqLOqDL3m4VENlsHVTuaxuYP3korPBD6k
fmFzYgs2IzXhvhg+Z5fJwoi4GOPBXjYlelIV2AiO+5jmENXsdSX3sarTmC0Gir4gZBzlA6790hVJ
154UcuZhFZP0gsTCg6dIs1fpOJCC3CPxMpNMnN7S8IKYlJ6h5A6MR3bEgcXMLNgU9KjcJIR8DRAV
IzLUIvquNVzctc3rZck63kHHn31cSAsV3o6UqJq9CAABEI90oWysPQ0awUfrMu20uzAOcfSAy777
lwGC0Cpr5fPoeUtAqAR4oX+Z0SYeyZlcqktk42OcVj+E4jzN3uVgxjjVWwm03vZAh5Vh/Zbr5J2a
Yd2Tde72EAgeKFoMfUHEX/lzLWkuqAbx4rOC1JWgSTt/Tp++IdUaosksfC26g460bztPuM+31FZ5
fG0+HlcdhTypyWTp3HsqlZ08/LjoCxsNvMbXzloF4DZJwYdXBjFSVsjhGi4MXMp72SZjhJVMFEZg
YcBFXr/MHIt13Vc+sjq/9/ee0uZZy+9CRrdLd0tlSA1Ayz8zjGWj/JeQICmJnYoKjwkb6kInqV3s
bcKpfyA68ZhrtVJk3lC7v2TngyHI8YdA/wXIGFOQpwAMV8HnEhhCjjjEb387CPWUc8jSPTPWpMi4
eQGQ+HBI4gSZLZ166rJa9xWMliD9sPjg1F1lw/bAOfhPvCnol2ToFEwEl1JQZMMH23G3xMBfj4As
5ECdzrkKc+g0jVlHJOx1J2l2j2ccyLradRg5r5GbBxEvWJnRymKYq5Sma3pQfHPfHefEmMmxJlYl
rpb4jfPMCuSUJUHsICCkBVH0i+SlzsjEGL/gVCUu7wTuMSE5ebOYoWzIzdcr3xqZ+s7IyLyQlJ1b
mPZdHiGkCJC2sZ3tRinGAQ0GZtzBFcNmglfRflqEjrtgxZtinlBQVyxH2uYFsIvhN4TXiOcIptHM
UgnCRgt+yhS4U7dfxrcEh5gHddp4JbR7xLkIuaLQOfbLr3Q51+anrtu8uMb746YuJupfq3WVM9Qr
aQfyy4jiMAmhdjJmGsv9yKLIK9QQ+vI/iyo4CHlKTYp8jkPkO6kq9ugUGu3K7nRwyKLgQr30C97j
87RLUgXGXrsohtjESmDjEVz1yGJFm2xpTDcnnm2ENjjkkp2C89uXVgDw2sqFaVxIonxq7+SKCMbT
P4UU9HO6Qc/XJ1gDsr+9rCAQi+HtGaacR/KJ1QGr9NnQMw5BzLT+p5fkBDARRNvdzHs69UMp9Bdx
N/ltsejAGdADgrXQU7vx+6Djzo3QLMETFUlbOqfUWJnwxPqGPYfEllFRoPKZPid+oIGUviMDMFYe
Xv2fcFtEuc9tZOdWENlJAWiWAdDqoWUMAf87jWRidY44ESuSUzOHbebMOo5xm57hGO+mTzwhvy7O
TwjtGX0kxUdfA8wbZPezmz+YXW2PsYQUOxw89vzIkc/gnsl2y2Ks74bjzwI4RVxVI4EVsgpRHBWj
ZyUsVj5hSg5M6YOQ6uFro5Nq7vRLlnQ/EoSPLgKQrWYnqw/9ive0AXVEboZjfmHKV1eMAUkmTAgd
mSp8Hk0OizXTKV6E8Ukc7f36H1nKd/MxWHDOWPkg+dovZftlxbW4FX4BGrzhbvwswjCA0NA119Nq
MGGELZLsHk7akQiZoH9OQ9dfcFcwpU8LsiN+kZPZqA/YwS3laKmwyMT4jLc6W5l9OioFpM2eyIom
k8cPHdgoVBet/SMSebiw+Oo/CZXKyrtXQTGpUBnuvGPBukWldiST5n7hxNH1Lzi8/DpYfzfaUEP4
OlHZUCmWfhqFCgR78Drhjq+dreZUMiHIaaHKMyQfAqELnWfa5fGqGx/IBl6obyIPRWOziQRT5bMq
9K9P1Vwy5DntWg8n2k8vFcpIX/Du+bmji3da0+g3UvzIGVj41yg//0C8Qsl5elo59x1ko7ATpavQ
7T1WeAbSewzG9yIc02/lLUC6kdd8w9FsFIt8viLDYjloQRYPdRI1bM9AGfY6ncrOwjjVQJJJpoay
moSiPoVKFK48yEYIkhFpHrbR6fRKJT4hf0ju+SjAvBv4GpobzVBTMW0rB83IT/o1ge8sH4oJsnp0
lX7UtP3Fh+qtcsjZjRHnpze12Ev6kfvetIT7Il40JVx7xdLJcT5cRzFq0bmMtpbZfEa850HcodMu
51XeCotpNB7PvzqVPwDj18OqRTeVmk7qumdgoqzVXj8KOqWIVuDOe627nOLJ8LDTC5FEmSGgHJa4
7xL5e0xd7TQP89pROqXsHyIPLom+P88N3TrBZcfA2UnPvx+I5e8TSsy7aYlz94wd7QON3ikHb7uv
ZbbxiUSq0lRiDqjztX252K45Y8AxDHzz8HZuB6g4QfufGCofYQ0f+8bCk9HWxtkzKoWh0NCRk8XI
S96+xW9JxJL8M+3w2IQJIE/9X3Wo9fEeBPjvockIje5w9a4w7QhPh0lzJkzFckYr/jPZmsVVxQQV
mvLTKT7SnA3X5RHoZxGj0zFPcSwDbxvh26oXn573NI+Nk2SCegRHcseh13eTqeWNKt0ire2nMEeJ
sqC2vgN9HXhKA/9rOTtUM8zip++jhXqD8JMoLDecLIvle2TY1qz9dRC5afjGH2TO04+6/6O9+vUj
UPc1utS+c61HYp39jda++IYuhdaMG9BCOoxTUT/SmHcBAji54cE9pNsuBR5fAriIR7NN+zucfdyl
FURMAXLL0GHP42p24DM4TON7hZ/Q+UACYFmFPJ5yTftVeTCJqX49QKC8/QovNeeAYR8X2+s3YiX0
zAdOrHHpp5LUgqC6H1E9niX8XTFPo89zbyn2mV26aoEpgG11wSp15Y66epO9HGA9lbodLaH2PgMG
++rxqORdF9F4C+KKZpwubST0f/HWJaHmMXEH1Slr11ED4DVeMkjywScB34onGRMzg/Mh4fW3g/ph
1KKf/Su8Dk+VacL8INspJulhDfZQceyBYsEQW2XQAHQSqv0GGrTnjDN3GN/FEL3geOyh5M7xC5X7
eWj7zvdm+mQ92P4QCAjaLTyGCeXUz9B3wTaMNqmepT0gSCvh9ofThBEit+raxZ8aHmY8UAEhTi98
FjrBtfyQpy2IzDmsiDJ4rmcunxqeT56zZ4jyYKHg1UoCXohbYlgqhv4pZORlOTmXAXaL2TCXZlrO
VejVMKxG0f6eZxULaA+opfYMvEF8NPESKxOxst3pu7+suHHc2eMrXmuqnNErLXSId8pCjHh4IHlt
b3PlZVJthypzLRQTrAKXsefZKekHfUCksKz5fOl++8G1FWGZwyTbc6802iWEAoyBW1FXXcxn7cZe
VnQh4W3Fj9jkGOLjp2jCqf4ZiCen91toNGLdKMCW7WBWZLHqwLT8iWIJQzRDRcooOdpv5W9qnX0V
UoI8Gt44Hvh7b9bXEoVQOGZWS2zHFIt8/YrvTu9wBuE3ExVvxdgSHKm2tiEzkJ6/844nhS/U+vgF
19rrorl4i/2vUVod/nZnt9Dci+T0ghI7vwyJ80czso+A/BBxDGRLZyQV9FoRU1hFGDPCS2MgLhjX
yLXdJ6zSg5F9Wb8urGCgenPj8cd+0R6Hn3OirX/JHtZISHNeZkT3v0kFmDATF82ujU0pMZffaHB1
5eXaMYKxaquM8uIq5ojvlim6eoQktcbp1f5lFAfSK46yTOLZYFkkpD+oJ14qaitEFpy3cu3kDaHq
o8suP1OrXa7MQSXgsJzAFP8XlCjFy46rD7vMA6KAeAsazz6fc91xbo/oA6bcTCEVTfBUqS2bX/Mz
NXwZ00ImQJ47OtOODzT39NNgz2bwdkr8NDsj1496tDzxIWmojErYMLPmwuUxVkXoQZbSbP5NwwJ7
3WikKrulMY/Iztwr3pfD8u+e7jPYVJ385FQPPSZm49QqCqEY8yF+z+ADJgcbHNeVbO7zmjThApcV
T0BMqVjZQWZyuXCHVwCSJyugAeIaLpdxHoZi852yn4mFdmJr/Z9k+B3bfzlOVdVQXb8pYYC5Fe6U
YNBGeiguhdDDL3svSf/hPmOOyVnzn+XIlqmQ+TjXjeSM1sZcKczjQHKOuw7kikkLFk37l12RsIiT
R7JPyNJaHGNOAc4Mj1OPsqy0h8/Z07DkPwEu0MxHR/oz2r+jHd5LexjndV10Mi5LqhvsFAbO06az
ipgvkw3wxoP/2jfehOWti/Bo08rP0ObkKK5NiZx3KoqrkOfIfcBdZbpsgBkPA12kxZ/l6QLEimsC
zuMQdC7g4+j+57rOEqYZfm6fYK2W1yEFh8a1yhbh2qLQ14ezSBD+uRROY0Kd9yZ/39mJa8ZVWaXq
ObPDvlGFKldhtkHxtt+73bcs0/9BADfDxdedu/TcD+J0JvtVspQ2eT7QtLxYUUDIRDOHMa5qvFLN
8t1LNbucqoYXHAoNhX12eZxA/tvTFBkrOAi7tEABgXxAV89VyjGJwQHuknZ9ZW1/67jHcwTeo0Ot
96DRTNa9mk4BmKek+B/NUeRtR1VgzF3Tu3dxkHOAcOD46rUR4Z0LXTK/JrgtljLg3dMQVCre2ig4
9RTNFPYLmntMGhgW4AMwclL4QdbL3xL+EdWQYvirET+WRid9gIIuxD/9u0su2rSX3DcLNYA2nWM5
y9c582Ly18EBq0qVYMg1kPpa9joW3tUkkOh/pD4cSpVGhUrv5ATZbioy6Hf0uwGyRQ+wg78Y6phW
IXD/fuNT1zL01Fv62zWG9QaIaO0wuTfsv1jHGuGlPPoRVP7IAMGt0vSSWEhntIBIcHnkkTeWOlos
I0rNbLHT6nEjSHqq6IHtQSieREHAh8GDNVkNPXpttTcpb36zEwrfqcGjxb7xMifv0LII0Zhur8pH
cdzg5ZQ1Il10141kTfZPv03Qgmz6DxTyQVK65Th+cYaSAHp05OvdgYjYH3Go2Kx0lm6uAYNOlm/K
Io74eXzwEAQBiCLy7IMwWMMWplEBeIGfn9j8yeVY1bWy+sZ7988UuyMD6q/0FRMIQIJOx17nxVur
zQa7qhUNX+Vx4IKlMr6SnVINxxPClFQ/JZ4FeCq0vzhCMIxoxE+/yeCB3hXnjwB0X+ckDZTIB2iY
MXMAzilMmFmUgiH876K8bw6/f2PDFVe+Ulb7Q+pVDeLEfxW3Mi2OAH2ps4fscjMPrRNn04Rk+teP
lU5oybT9eXUYQPxSvk6Epc6U/5Ap1Tb03pnna3iaQKP7svTwrWYbsBWhJEwd7s/86gpye3VrojlA
QCRxtXagwQ6gTvxrd+YVDeQafh0bjG/L5MMSOmBg7DoSa/Yqu1Op7IXMcgDcVX5z47wX/7sJGMzZ
jR26uqoEafYdIhPFp1oklQvTCbtGA/KElCSkrSn+wQOaYAHFmGV92aYSFuAlADjYdyV67A1z1yNE
r8HvfDhke1jL7U3mwIs2VFfWcUlWZR9MiVBFG4tN+o4T1y39QwvUMgV7uKUtdXZz8QUDdPSpbL97
voTh/d0kPiFYOPIh9fQkwejg8Hr2wY+DxJ92qczKIP7gQxQRvpWGAjHSh9X2PGukUxOCyk2nm8sm
bxQRRlQ9p7skr0otE0vZ9b1KJdmqJaPSO42Vp023FO10z58uuzOqApLjq/X3hozA0IDzsedFNGOv
NAojyg/U+wS6uGdfR/xbaQJhd7DtK0p1gRX39YCmn5P023WDYNJrBcyidcPA86QdpT+uWBiRoZlE
X+xxOrxM+aaPgzIs7l7qP+8kfIMxnYYF9QZ4l0DoUr90/r4cID7YpNS90vL12VmVO5VdJ0eeZ0mu
LiULfqb+odX3eYv5CBVEobVijR5NNpbqXS6Ma3HB+kGG06ekUonHYAEEMHHkDJkBo7T7PTGfB5b/
4CCFNo7O/SVTQnXAYOaQe0TmKDIa8/SMSwIFznkeueBQEybkeNFDN0wjPVFHoGfYd7EPRpAZ9VNI
+EqPPV4TuVy1zWeOtA35Gb0Zr44Z01hFAm2AGm5qLpmI+m9LAnAN6xCkPgaf/PMl4/LgBjkFv1jv
bDFJWoSaaLUIIh3Hl83ZjTS5H6oT2qpDhfAVgZb+BEbRSJdzsP9li8yb1iOt4b6G9UJnMbj41S+z
8yz8hNNs60YJz7thBmZdWzNAdDOw8lnwPttyJlDEt0WpUyQk4Z6FrqFRplxJWMnZUpL0sN8pc2XW
kkbFZPeQSq0tMEBcxz+YH7oi/xOmpdYcVmHeoBbMQy5oFI0F5+QZqU9AtZ8s+2db2q+MeqRbKcv7
EEjMfdx1XBjlmTlxqzGLQ8aQPOwO0NOeY5hwb1/JsdLH3ObTXpeL2Vn/5Sl3hZgt96yBzoa7T4As
1XAhiyWyfLCQyyT0BrfZykF8zqvuRra/mlfVZwB++QmUoYXePkyX68cWpUZnma/YzJ/upFZALYea
taIU9VT1N7tNr7KXC9wRHyuwEJwICMBNSuMwElBBk6zIgiIiTXnFi/MyeTwV7T71KpUZZo5+1s7Y
+NUOvvBIKxzTl4L2g9b3dPKWIEYGTMU49qmJ5SPenEc9VrpyJL/XpAjgZSTEL6AX/ZGNJGTeUaSd
XFJ98b3VGFim8bFjWuFFqhoy/Yjd1WAABjtBmPJRIJoPODJzVChqOznWCyWIl5LN7H5Z8e8RloSY
c2CwB5lzDPZsILbeUIWQeDaf2dpx/qBESCNzefkfjT+mj3VZDTtufV7g1s4xMTUs5b4EVBlHDWKO
0/SZ7S83Iq+PSJdak5y5Hj0GGi4ZNRkUuobJjKgAM18mc/ptkNFk52uiQPLDQTLzeyCzYzUXvge0
IeDnWB26LzZD5gLuxu5b3Jh1bbZ0PyGCsDre3tz7Cf3MWF0EPAYwNwfoEl/54hqSp4F8qqTQggFt
cVKXvCqgNAgdj6EtKF2ZBUILzbMY2x+sEVNq+Z3fA4Oj7TBz7yx3Cbv52dyD9d1bno4efHE70eeO
RHAOkWWo+SQCqyzQvkY+0iY1ZktCsOO205fhJjG8UmEx6NXwPCExWsQoAIW754tlXfrR91BXWbkd
ceT1xdd6oDthNBcrsY639wz9vPqVHD4Ito+Z9R+sfb1fJJqPelsGiL298M+592g1f4JXPhMecpH0
ansQ4yBPg8mYyxFcSuOdvmt5HmT1EAdD6C67abdt6RXLcMEOU2x7rdlX3l35mFWiAepxaO4uSmDA
aVP+Ct+x+SwQvVr975AnGJZTFcC/gdaaHKMczhsM5GnrLPR1r/hoWZnlICkennx5Fkt8yRA5i/ky
NN/HBDPUxoYEML5ZZQ5bJtYsrUCWIz0eErJdvpe2KyTv0mD3WqMF5uOVHGbyBvHGJT/+XVgU7+4J
148FMJXDWv8imQ2sKNUmA6QYZ3vIqOGETfUzOUgrjfRnQd6c0KYXGUnDdZ6hdWgLyBv9wy0tvGOw
VDO+9S3Ss0bqCh9HRri1LH+i8TgPiZ+l5430nyJfq5cM4Sxt1Xiv+YuynwZhiDIatPUBYwJxHXgH
mUU3GQe10m84m2Ys1qu3KZoM/305V1cxqtzD3CeqKPrrnlTiOR7ElzoRG71BLKUfAWSp4E2mLH3x
Y8QIr+J9hH0NyhkOegw+DzPebTvMLvRoXDu+16HRP/UwCtpJ4gKS6CgSAtSxykQenyhRRaSHw36m
MuQDDf59NcQLDk3oAn+//BoauHbyBKpmuOvjtnVonN7ea9PbimsGO9SuUMLH11gvbDyjd+0pYZRU
Z4e4ZIxuWXwAS2XAkHuauyHeHheuueLAlzAv8oD2MgHyj7wDBsoDtLTXnItWlv4ojadbQ64GWPp6
iDNRiZfFepyb3hoahaHqstcgoKveZJiEpKnZGWcFWSMJo8uyahw6M2uYAfyZ4Da4VFmrXYOWpnAO
mUhVukDtRbvu59LaPu063gI1KXaB8n0VGGXQM+oJSkyIvvSU5GizujkOf6lWmakM4ONqMbyWflIO
j8TRFVNng8ktGrzc55VvOaoQPaqpHEyc9JDDtJRPFsgWEooX648DgjWtux2N6am35kzPvlrap8cF
QbGIiwQ5oF8X06R7IRhi5hPdwA+6oaZC2PX1lOnZ/LzK0HYGWcJK341v7csZUCiR1fqQCI9bchP8
GSRqt+WHg88EW9f3ISr/zpC/IArPEfH+Wd0kTJMpWpynj2uqslxk0hbr1xD7KFT0ur6ixGkxRrVL
r4j+LJB3lbFGG+X5Xjximw7msigLL9y2sKQYpS4GhEt0lVp9eTOjjvoJmMxKFdgcttcCsILzJtcj
PpIygQFnAdzFWMFHy1+zMYvSbx9b4pCVE7QGwNWrarGyPqIHC4+/0StRPlUwrCyUv/Y9GZjGYenB
LgD4p2ZMVoVpqoMZdte+p86y8TXysHvbY0DBoPtkfl/0z13rhMjhIoNkXQZS/SsR8XUXVA8DNgVc
NwwRV2meTtmvy34Pkg7OT+H5NZw8ZrY21y9L0rtNNgOHg2XwGZ2fn+rTgWhbEBbqO69k+iqPe9rW
Q6HD1n5zFajSyWEmdTlGizPEzFoiUnhDDl6cBq9/Z73KBCB+5R/Y5JhK+qHPFUrnmjyJmUw8/RUm
BAJUaxbRjm0uWG6BurEZhhgr8MNHyD0PEq7R+Ya3qxVtAXvNcL5x7iBxq3nUrIIcKOfJa4oJI717
F7Zy9EpJt2FPwbO6HRx/Bn1BXD3wUx/VqVPMa8XUdRnwCADCm17dEkT8JYqSy9OtxrVrcP1cjxZE
J83M/OOtzdYvQATA89bMweZXuPfzvrNCyCswSeQW/mav6fUR8PF4e8IA5sFD174/CwL5VrI/Ro2H
ZSO4hdxqHWBakaguOWMVbPi3UzOw6KCS+QSDdLJhzojEtDeUpik71SfxFMMpjXlnvSaBTxJRSYjx
lar+t+XJgymEcnJms0jndSyU9KV6AvlzSEuoY8Rn7OIgs0psF6oUlECPmDAezkkQ/yw3hyYcH3ga
ah9sMo37uVJP6LruC8gaukNBiNEf0JBG5C07rgpkoRPk6kOwOHPk2KFjV/VXvxqOzwNBlTX2yaa5
lYPXlu7VfuO5kX7xD/EHDBcY0qdKFWWzRDyAAdcJ3hASoTtmeUXYi3z3PBIQvWQV0Ms2JUdD0+iE
5j0xHtlDDMUwnk45c4v5oJIg1YrqY1smfHaRlgU7CrZZkQRRpuc3pCW+jPr5tPK6KZUoAVFxR7ao
F4NzoTRPVj80e+N1AW/+W25c4en97xV8HJXBw62xClfeO/HCr8LuzxoXV7BUnbG1l2DYda4qtiL8
WrxFFyucznPGULNOgn7/3r6WF9NIGl8S8gWBm5DgUPcT2+hcZw7CF+H2tkB+vyuo7WS4JGkpHPSg
XtfgtkbdCsMnViburzeG+XiQ7u8opPL3y380u9VYNRS3XcY3rRynQ/fEY4Y3UfgLrbnMdD96dgp8
LhcmGvnv2ldRABhkq+H8wdlJQmDO77N2XQLOG/88qQBpxQp7LBB32v18mEEyZVLIrf/MVKTIK5+R
b0vleueUMTPoCmMlUgIF46eH9idEiywDdPzWAUx+/W3XXFierU0uQOoeg5T2gE+H6J5K/z9J337w
ymOdzl+cxPxR0cUzoU647YTHQjk3UJWAWY0vgX7FqbQcHJ48Oc3HOmZuzwCJionYLSsn2ENZlWMW
bmlE5BOBBB1EYONhrHtI6SWwdNwDbUkHWw9OvxbdttVTQDt5VtPebBNln0u65Zo3btAW4Y0VwPXq
L34KIiBmHLnhWr8vX4wnXQo0mxC/2E2eaIpC7hl8pp7nwQpR5p35eA5HPHWNeYiH8k8XSNmu+D/8
aYvUPDYklGx/7H6T9CwkHbxG4NbY2a+fEdZ8vYtFCHPa8cC59iuEIhSgnsC51pRWAlxls8qLjYNe
23f4rQqEyIGoqkRRs3gsiRJ3cdWMGQiRMyUhmULwGbWTiXk1FaW14TPNbrBBLGHltsFDNS3an1mp
LeCAYhN1OB7SJ2+KmYwZ9hx/h2INoPLAEQWTkgE8uF0Ra+lJ8myPBa3SmD7bKkYAXtItOeFBj1bU
BhnwyLtJadgMxJTr0XXhUTVgNu17VGb6R3vY0oLRIH1RroLmk3SAn2WcXG/pL7SJIKb0gMiH+DHS
WezAg6mKyY9Cyd8dE3PvoTrlUT7vFe6/FCV91nLXDzbov+uP5qgZ/C/XKseyk4xbpeBP7D2MGZbb
vaQ07IDon+Ytk4k+SkbsQQHyo8ssULXQnxn/FEwiJz/VGYkJdCmI3nIn1e5VMmWZkSa0TEBPsDoq
QW6QPJyXcuenATCuuED9popLsTCOtbVqeQ+9E5/M70X+XHLz2f1ctVXBYVUxeelsl/xzLImWZv1s
6kzYOhYYz9sN5mLdqx/cAP+Z/NDxsprf0rU7AJntV4tutrIyhaQeMJxHVgYV7Z3kWZxzWqMcDoVf
kFv4cIg7TPhN09HIzEfHW/ZzrhRA1OB7MzdJZcVH5Jh9FyJGBxxM+PtL2BA7WRP0QHoOA/cO66DF
4LyYZVy1R+MTu3BNjRvcNfkyOuI+ohV9x9/NtGxWQZmsRDMjreOdDo10GwfsBRWnQRifkKIyQHuY
4MHF8GGSbc5R4tw9d3K+ogUZ8A5EcroZhXhsE+EVTB7souFjuRjrBQkst0gBQQVm+zji1Gxdxp5W
EHjgl488p37qvDH5dvNF/0KykB3QcDgfPJd/ctlFJlqo8qvrqjxPedax7Kvoa5LCQvQXhlh734bn
EfeDU1TgSYvB9D7DgrQkQA27B//Mwmzbb6JKtKmgwwLJq1gsHk1mXqHAHnK6QtxUWSa8oRq01MY7
30Dv7CVD5+cgWB9XHZvmmn3pblDtGiAZqXXEO8q0IkBUgmAwO9s/7mvKS5F8jnAklmI3tfMTnEG+
kf9OO5aSsznF1efDyK8r7zpqdYSzEl2NL/L+p1v3zuRxuKpjA/o69+g826hRFuLw10zn/ou9B3Mi
63ha0ZP3k5YG4j06BcH5Y9phhal4/iGG6KiWworcEeMiaZb6YaXgIOEQ/XoR+wzSPstOyh3I8cFZ
JjCqZ6UYCuRaO+igQaQYjMj/ZkwQcNnHhPs0nJtbdkW8ZbUNFBET+MWfzb6K53MwZTNeWLVDStZW
BnTvxWoAhwLAJ03xzaQggU3C4uLtWK/8nikEsfmaXJYpAofDXyk0SipekDMNGBEN206F/S63ccg+
Vnj+a7NYllUDwevrTh93dTsCDPagjjdY+GHCjQ88VwMzGOQTTXNcl/1mSvJagOd1Izj9FM46pUV2
sjTIlXAXPWgjDQxmXG7P9GKiMoeuYGFJiKGvw/e9OGzuLKzxVgoJWOyeWmJQ8mDHjMHPsTwZz51Q
aZhEk/LJbwclS535G9Y6pXrSB5gH9IEes7tb2TJ32sf4oLl2mZ1618pNHl/PVSUrghiUQ1tHw0W0
M39BXvlpRB0XfMVCq6BB60NPeXeK1IxqIBgHJIUmTci3W6L9y435h20L8Stx77J8oRtgQN2ZnP80
pCrXg0HyGCkd15ZeJkrCipl2OULBiU0jU46fgzAXJKR438yCgBlTie1RsWsC4/OIL7MzKLoYjDnE
/fSS7W84eKdKaJFzb5TdTAyUZt/G0589daa9TLp1e9q7WKhPF8nJw1eSYluEpc51qWjTQ2XR6X36
ENvEtdJkR2RfwTg/sPkNlrHHae8jvRdp8wzbg1erc5mTo6RgRs6S6BwhqsgiZL9XiezolinMYmN+
75qm0nqO7K7atNCqCa1d1vR1pav5eIDD45H592+2rHutL9MCdb8WfuxhMhRxTA+aq255wRDrcVs+
4AWcGdIJncVgEsKG2YeLwPH7Kj3aKL8L5XyS95quEdjKllIMWQ1k4T0JMuMbJ2/K6qsVVx0WBKBP
YRZtBf6TnWtS6gCG5DFlIp+bwoipt24ueX9HsFCgQiK50bp9Tr2gbrE0Brxo7RuyS2v20gAKjscz
Qm4ro7z/JFqqEDmZR8cPCNxqStzA7GvCO/6UxOV8zcwBH2iNtxIRgLCLiVHjj4aA3sksQq3R2Pry
8t4muhQLo++5fnW35z3DahemUt6O3ox0okEypK7ZPAPK8HvAlFlu7hnJUCRKOPDYhpiFDko9rgtr
NsTD/HU1du3bpTFRpUxvx0ZzbEo7EgvCcNCFZZK+VqWTEpVLC8jcNjrXow34DkrfcDtIBKrjG/K7
g7+R3xGE6L2xG823H7A3OvNOFNxpXuEao3d+XvWtG/GM6zkkuT2rgs5rGIQTjt9N0UZTdZMDyhZf
Li8p40oHlfIYsNkPe3Kuf4YjM1PdYoOl8phwxihEd279hy7AOXup9luo3EPx6KlADc3ofYiJXcui
IUI0V8MISK6BRfjIlkuj9jsVz8D8I7cp21jsZ/ba04KcczRMDeL+VU+IXZyzhzCaGQBThlWhh+0h
O1hfweYlWnb/7qeIjKDgvGzLxvSq/h+ZqjO6N7TBUclLcPCT6IHSwqNn9pPNMXf7Dmvx+xl8+VDz
TVoQIZ3WBG5gjILS4dJ1mFBANzgOqxInQWbPHHnJaBvd1b9PpEpsiCZ5JlUO3vByPCzB4I9EpUWs
brjliUT5L3b5EBXz+HdcSmwbUWOe2f19e1uT3xYt8OjINdxVJvFB6X1x/6/er3AtLbXhQFxC4zxY
4WiRxquC+/KB5kA9bYLObh8fo5A8KyRlyqRk1lhm95hh9yv0j7a7apawiEBUqIOST2NrhZ/ONrRB
SNJls5STgKoPDuALRvqaUeBCGLUnRxOmnDb3QMhsOoeDakyH0RfF95f6ywnZ+wflKBctWsJ4mLlz
J1OnGUSZj9x/apDoMGsfFHcjnrs4mxEJa0HQiNcM3mmp8nWn2Irz2khGCjM6XujhOWP1Nd60M8XR
IyRMlzoxjIAy/Npxsdb5hRNpp/XHTYpkrrjsgD5gcNZJDkV6AS/2QfGVdy8uHowO22KdKIJrccou
hyfdwr3gO2tfwxX4lpOJPhl94sThcTZwXIvEJQJXBiW2IBOto+Px2aFPo3fR9jD/REFmnGVL3RY0
WbHs6ewawHwq5tarEQ8ryAH2c8xz6h5EC0zgxMMEeV3wKMLcAcOIyHqdcAwGC9GR6WmRLj+nAVfP
PN/OIwy1+XpqEGMmg3bypGcNEdeFRBus4lGF1UgHh16OJJYI3ymCBkNN04GLaaC6pmqvO8pAjF+V
EWrWRSpYVp2YVnjfRQl2UNTJXt3ba20Gcg/UmmsUj2efJXRY+BucuZWL599xP2BKbaYkThPNmuuW
WcP1C4NmBx9zR2bA/8YAVJXKRmpAYFdOJIfKXWXp2oJwLWa35ljutFkvHnsH/c7dA7II6uVe5tgT
NOyIJPxfoNcQno2XGBGEwQdB89G7f4oGzxGV+8jsLkhzsst7MUvO2mkR/LMxNuhO0eIDPazYFX9T
X1KqOIxgi3dTdYYESlx1k93M7z9QYyUqT3HgXcM3HtiPCgvVNQL3H9GeMkBpp83oBadIlkKe6Jr5
g2HoYbxaq5dqpJqLZYqrdhhh8Bc0WrR1+UjBTDOxS4QaMcTxI7P9qtxVdlGTWGu5RpHVTUsvHSAX
JpamyisMBcoQSf+n+fy+jL+fQvoiKszDxDF5IrYhWy1UCrrbmTyUYZnf06wlPPC5KNN39RvIwmHT
yndc1Jh5po3aR8ZQv10tqLs+u+dxiR2DyAH/awtoFI9xJ6AJQeaZ05MfNDyIzzRmWqep0N6iX4T2
KpJMAUa1KuQkDcaRXRKymO4ViTcMs+9OQvDYnQSCphnPya775QwlJfq56QX1eOBoAcalz8q4RvLt
H8kys+Obfvzz4U4oI0MzsEyPmWEh8Lp1m/8xfmtpQje49mmEnyaFtnhK5HplLpHROtKSqJ9nFST/
uueFiHhs5zpDKF4Wf0eH3dHf2KQM0FFfvOf7syGEC7DwdabggSQPS8HXzMfnZDO/Sn20J8cnl/G2
FeBTePUjOMz5MvjhYMv09xry6v5HDPYNErL+kc+Ec1bpecn31fUlG2/9C49uGkJ+0KT13tdwkB82
+ryVPOjbEAZocjt8tjPvKyojIndPAKKLHzLc2iUkVBg7OkGKekPfOerBaCRYX8wjqBkHEkX4jXlZ
yx9yB6qPknBpn5n9NHR/+iPGM2H3hv6P/LMWJH5CsI/2l2lFQHwsh/knXe+RdkH6OQBVP0WLX0XD
QONIBkYd8pn5tfucLTq19DW2X+w59ifL5B0VIiUARzg/1yYIe/ug0hoqfzyOM04dJqZVYMRTLCfZ
3xgKqOc6+zwkWhcaZIZqzm+cJiUBObmnl/71B7XUOqYxS9vj0nCd0M03BMbe3sVezYZ8SfaWEGXa
5i7IruINScamNj46qV9P9wGLY2QDtY+mLP87ZVZgan6HNzFRZ0pMnxko1WPXFjPUwS8gS7ltOptX
bL5qIJCsXTs/Ft1CMHvBO5EIXN8g0jLyZxIndx92aSGorGbUC0INtC/nlltcDqWU0rVuxqT/48/L
DuQ6DRgqR2WoAJ99TJbeYdMpd5BpA6C3dgE6HVEOcUmpIclAjWw6RyBUcM6LHjpbRt9tdCKgl+Kk
LolanA/Yjw30LgQABzVFnFRZtEE1/sHx//0oBepWMUf6BD4lzMeW1eA/RjdV4q4xG4nuh/nqXv/6
FDJaIn1tnsu7BFp6TJBkYilLQ7UYQ093sYtZH4zQDiffHOazFvIrqExN9axNsz7pKBrPxWZJP+Bt
Rj0o83MrX3iKztbGdU0awzIcFZ73OHtd9dXD/OPSJA7AWYoz+yoQwdRxGxjivw7/5QI2W/qffgVU
zpq2A+/DXiG884J3O+HxLiwX3Gm2ycewe3WeNEwRHuvcZdC5hiDJ9nmQkV8rr+O+JAnUVpPAQI0V
qG2Y5f59asXAQTPpgyhwUkGf1W90o9oXdCOeKtyY9sqKqM7+O0VzWgrwgVuJBq/+yTEWj1Eom7jB
sH8JX8jKZtitkEPmtjMawp18tWl88C8vtsAaZGxJ6vDhb/zuMSoH/V9iG+ZwgOoDvkfUKrngkiIa
7lWWIBnX3wylntjrCoPv3bx8qV0fEjW9U4ABnRbgREG1vAJ57HOe3Syj/2caQc+pmnBlgR/jFVJQ
rPn9pr1EhwLwZt8qxZ0v2RuQhD45DSfK4Q8ptR0CikEZTSEhMlSXQckEKLoHn5DjbVSHwFwMqWhx
qy5hpaRaidfAOLh0O4PWLOpxXs43CkWH3ykLChQ7fFlo9aFf3vzr386utn0Q5IYLpCWEerWMBHp0
VCg8MvZTgyrZHJ7WFhwKbUAIFz/FgbSHMAwyRA5yScuz2L8S9u0ud94coBRmGIUvpwXpihPjOLDE
z3YErk1huqVkszPCEg3c04HKL9XR90rkBu2U/+l8NEt3tzQOwz+x6JYxlC4GMDpEEWbyU0Csukqb
V2YFM3Tm/0ICOqT7AIOabBAhBw/PTUc46Kv+xW+C//3zB9nVGjxxbp0VIj+avffdmt9EdP6mTmSS
VwIVl3+HoiQlxcOb4aYwiY3HbwxVDuQT8GY5GTxgGriiZscUWUVXRIZWZosM8ORG8NwI5TaFIQ48
T4NXRpTDq6OVo7G75D2kMlqYK7PQSDF1XLGyppmx95uWANxqjaD7ciKn215CSCWvvnmsC42Ze8z5
dcg5DkZBVZARbcHewhSXabqqqhFdrUO02n96W4CeJ5DOjDRHhlMy3ZVBDG5s1Fe5N/pnS3PHBgF3
oFTtrQk8Gh4g/8wkWtf6Zp/u1C4+B8XY2w2X9CthxEWurG/X3wSj7txea72Sn5g5OLXf+XgRtxC3
HTnlNXs+xZeUSMaKqZmnYOWcME+zJiHuq+vl82Rl0eo3kBaco3Iz/oYWrARFhfsNdzZWzYqQ9BiI
pRIN1cyy2RhD+boKgcBrfycrQdXnHAalVUCES+Rcz1S1MUJBLGG6z/z4ODOCNoEkqI+qbzfd6J95
0ObLPfbpqIrPbisIK+JQYX9YCsvMC7nuxEKev2WPA/y9bNHVnfXT8rlZkrdH2NHeeaL2VDNQEfDf
+Hn/K9VBzGK2Q2b5NILNjpMDc83rrrU9aeel6CHjntO+LtvzuD9jeH4Y1aOv2ECvEPwAOA44dXn+
BlaFxsRV+9R4zjoFOs54z7tjtFTYsvDvvkRq4NBxib/NezANS0qm7WV/ogkoPYRuGCCSPeRQPxpc
9M0ADUZuIaVkLt8CZgu2AvgSypgT64gjTeT9HTrA3BNuIiG5PjYAHZUQ6ECQu7/823XJY3x2CVm6
gtbIqkxj0gAagoEH8E90Zg0WR+3XKWKFAiEUqnp34X6ZkBITUbLKfPkdyjQA30IgbTbI7pFN/5Qp
8Zm3aBCcdB91LsVTvFXPMP8Ni5zMr7iCQ+LZgUbZGzMFymunsBGKiiBOL5GAFjAD9D2Uk8g72aR8
plTK3SGvbdT1r38/beY8dODgiB5rL/zz56eYENtJe0cErEvFWlfShM9Ku0Uq+SVyhl1tz/5h4o/y
g9oFlBv/6GQh4BfQQ21zOW/GzgTP4ncYO+DIOqH877piYieTFYPlu8MoNHvzZQB69slbHRGeSffO
nMHJWZYEvHwElEPBL7MwFuXfGmOr9Kp6KL82p5IO2Z7bRQR50GDoha8kGM43SCqMH9IvY/UXcAdM
QdVBotEYLlhZumb85RSBsCJoA97uGEtXPsvddT4w7IR55CiKQVZc5vps0wQDzVM7E/kZBmrdiJYl
xrK+Mz7CcFLWv8gDj345Uh/mTbpyisquMPhkT3/xrRp7SNgnB49XprB82OZGNH/KEsufYOVs4f+W
4/MsPBix93KKxrJ+Oev4u01hS7GGwoCN6NE8d4rmQ2uj+NOWYFO5mva8gEZOEazl/q+Ji8crMy66
Y5OGp0mnOMY8bhpUhIvT5uxtB932/RyZDDrZAjmbE7ci4EWuUVjCa3af5aqQ6fyTK2xYbwCbnJoG
VvHwW79/3Q/grQ0pW0cLheBFpHCq1O0Hg5/C8xqhWdzfFAlAIkVK4ttuZj1BoiCwIsGV9awoMKaS
k76a5+0fZOqwHqU3Ney13p+WdDxapc7Vks4yeoqS6qTlRuA2JTICKSBQYGfCRPkURzdUQngPyrDb
Wq64Mqj3W1SR0aqvUDQb0KN/z+Dny6xV+lUT+KQlwea7BGzPKM6LB4j0Vc7nBuLg2P714EdIH1kF
gSHIlX51LFPEyf3i/oD0nL+n8ydqOfb2M6lfNo6ze1K6mliiUHSRN4/Hm1X6M9j4U3BoMswOib91
spiXSwOntyZSiqqFsKEaMbQ7Jyg7yj8g3BMcynbKcjhNqao7gRZ9hFxE2jMwMQqp+Fh53/Jh4dL5
bJipbfCHqgltlXCySKXYvhqIYHKqMJRvKKefC9dVNUe3XenFW6DwTXVcafIQedkEEpJ+fII7ChK1
AONmPQq4H5Nn3p8DiG2qxmfVgmO8dSNLFm8+/c2uIL6bfhjgiRjvQlMLlMl8dyAdScxr7SQVP6bF
5rU6YPUN4KadcXpWNEF4RzM6gNCeNEiLfY8TwUAwmgHN/l1k6i8LEpejFEU/tgIMqvfRCs7Hb7jJ
iNJ8I7wIg4jD245hPULUwtDTwx1hqoSJovlf82yYenwP4AQ0RYdmEPyqnXB7Db1iG1J/sAjSOtlH
kD1k9OqW0FUvvMPfFt9/RvBvs2XwA5P7Tf7Zjw8rxgxATMhPqAJ8+1Z4aKceFE0txADmQ760e/f2
8oDl+hdHz1MrQgODMuRbm97N+9oEaaOClSyH5oFKaOINpq7cd6jp2aVpfDD5icPYjWsUnfyiCagz
sxde3lLnOLDffryxlizYKA6gH2H8vkJ1ENLqBR5pRer3BYgdY4mhIb2Yv7yv5QfNUN0b+nwPXV5U
TB4a9H5vbdf3qC8ZWzD1i30v99D+2tOIRouG8a4eVlW4tCSL+5d324Vc9ytFvIYkxB/RfduLjPoq
KFWsGlamKpkViit/hPRT7SGB+paxKWxMhUyookfShJqVqapT1IrdxjBtzZ9jjmlCN3DMC0sBXomG
c04LmMqDd9O5bzyHqp88FJFsG13LuSP5kF+CLOsWhZ2gAkSlaGIaI8ZnSxoUhvtFI66UqASDp2kJ
BW2eOm/dFTsykiFXA9f/yZKJdEN6YDaOE9EgSC3J7SAIp9u7xvLM6t+m50mw1fZXeR7OTAx51a/O
xki+O1F6HVR8FyqGBc1PpxDw5AcFd9+XYnivxtJu/Eo89QhcoGC8J9f2VloybHcNgWn0Vw8CTSmw
bPn0XITW/ywGEjhv+xmYUsTq/sgtgpGFnsBKMQN/o37LD3gJj4QoD54ZpkmXtohr4WFpMCco8yAr
QIW8qLjStsEilazNsTbBYqhfBoHgzeKkO47IQ8O0DZfv5zdduVUfeEmDN67mOmEYw5Z5sMshFHZf
PaZz8zeQIdMOQ7XJYjKeykTZJEfhTZNdrSAA9PXhovgKhs4qe1r9GeaTopN2M527MLKgE0qjpsXr
Cs8wCq21N/I05eX5ZMQs598GVUqF3Rarg90dGM7Q95SLr8EqODbUiaCqSJ6KV19We6QNHI6IvNOO
Bu3sDMcWO4yirlZigqIlJ2dv1mI7OxF3i0R+Yq/48D44ANxWeEYyX4Rinf0c1ke7nv5Tafv6OnQm
afSqN30sbPAXNmYurvt0WH0Vu0gNOBK9jC4p2FY840Sd0sIQErtX4UEnH1Ggg/Z5kaEnhwp3x9Us
Lut7SQvA/yamiRs22+/rohO7HvBk+D85EFW+pupqHVLHdXPpB0JwKU01kPRSjq0Vszbp2iD51Jq0
EFFI7bAFgGNTFsAx6TdFTsTgmDrCCx7FAuPUAqKp9h7HvilpBYLBZdd/9WYmQPX1H7g54qCl0ac/
LR3F4SG9HMGQmSKzyC5NWqYborPX/Ew25J12TceIkBVIgViSz8GB4OesG9d0CL+Y+MN11LQtfU9J
5aP2kr52/Fg5RD+rSkCXpp6YXs9Qa8QHNHKFROsQ4OcIjgXPaatGnQnV1770r2X737Bp2RgDbysG
RQvwC7dpFboeGD3ujMeuNetRgLGyDALEcNhlAC1cDCdfvhohXD6QYXHe56/xL7BXRPVMY0I8lUhk
Um4MyvQj7dOeqPMdAD/iDce3eD0CN8WJZMZrdDBr3QOXfiyfWNG/7UFIIplYsoFO9eYOQvs53SOa
sHR2BOvpmdjaFLIjXK3aLkkuEcPNMCZ0k+2sJ6nKtYvRcrFMFNWWKd4c8AKtAIRlHkPJBDxp1i0Q
5fwXDZe1aPxbxlJgVGRbAiDKgWtnfZqilIsEy5OKzBqxrEvjwzcVpTSDlP08FtW2QG83Sh19KpCx
5B6zEA76qq5CdcKGWH/9UxV2LottGw1a2Ymx8XGoFvhvXC6riRSbZwPPnVOFIlNfnXl0iTXO+VJY
og2n9UTRLvKRYv+nY4YZWHn/Nv+RCS1z2lboT0zyxj8kvOtteo8zHS6bXk9Hlis8V4aRsDCbciw5
T3vIz1gzYyLV6X79BJwsErwdJoRswmZ6UfX8HhAum0SMGaSBnFcFnOX6eIxdr1J8om46U+ylJwRu
EATrga79J3yilnIobsTo246MQhg9uSOwMS2hw2RPUelpz4vgPdCj99HtU734cwuqFNZYCtxIQeSk
EDsXhunmqup/zHA81dHedwFDCPkGhEa/QU609v7aWpVzg/7mZlDXExI5Kuw2m9CJ7DXuCULp+03R
2tU9a86Dm/SO3whizAexLZ6cK4k6VaZecz10mqg6mZSQ8jYRZ3gFtgpEBs45mvro58xN5/hJO8gc
+WZJ/aiZn0tBDBAsK1chiqIo8JOJK4CBS098Y4qo2hU1KiNezd/GrY+1o0fbkM3a4W6uj0UtYK3G
U0BXyLLkSvK27VOc4xY95XWC+2fxWqqKIrqDB+TSJtV1V5AuEIsL0yE+zwleDPMsVYHMbCXe3sbG
PhXhxu/ssJd/I3M9eE1qC4XqxAsHJiDUDLQPqbULhLeGNArAQt7JpnSTl9P/SnK9D7qz4Xi7vQpc
EJndx8/jnbNUibaBXUkDisASpuquYpe16jgRUUy+EOXzLAoD1boJikvmtR7GApmizcBmpYMooJZy
yFVkdRrAa77VM6I99P1dbZVSCfmE7Efz1iLV+4//7Bwypq053I07OHmiUJfqO+3qhIsrGkze7d1Z
B51KtjoiJSklE/SoOzVkMtEI3t27MLL9JuCqlWvE13xEikDHdeL0kK19LxO1KhLeppdvcBJNjw4S
qh6KVcfAGsjGPpiEIJ+sFDg8Jls6uAHN1yBnaHx82fAeNf9SjYRWqK3Jk1NTQoClvlH7mZJB99aF
vIftG2tLZyGVdulpVYSqiWuj7D/POXFi+HvdZ+/HSlQEHHZ9Gr0I6lFaL5gPpkGFTIsk3On+Y/KP
QFmL/YiLV8gV6lJmRS2m+YReI2EpLehfUuJKcPg9BTv91XKuRRdJQ7rB8J2Ne8HSqiQ0OMTRauT9
T7ho2/ahryiwlgaA1bOR5/jaNrFudYFX8tbLaGtfvFP6hpCXv7mjUMJlN2qXqbTvBVmtrEHvhFiX
FZzBMjWxySSlYOTHCu5WCJtwcMRxy4mQR8pRgHfD8PTVnwhmXP0NPiAdyIjwLVD1iHoRzRVlQ4/e
rBqjBjjIAwU4vB2xj9jQRUUag2yh4Pd1K1ncaB62sR7OCLDajIHDLjC8gm0dEXF/DnoIenkIQBZ8
ISMMMkyTIpjnb1oPQtGsB0OLSyO9n20f/sJy2twkHdB82W9w6n8deMK6TIk4uCH0914j+T85t2QT
0pT+faWDc0NO5Qz574zO22UQDMnie01gERnRIBIMAjyrKZIK7vvOSRWSPanNMfeTmSwt/udrpfUq
WboneVj+HVCMPwQvnNbRDivGe7+DmhUpgM2iRX8dJSXQgp2Lk9rSn5kD9XoFYREAs7O5dpywcAvA
nZKS8yjlNmUhu5BJidyh4G1N6O6aRtdU7sRdri0/6CuT4+EALvsBsreEyq5hBmsSqtBtHtMHGLoq
hhQ3lRiuxZ1Y9hCtPig5YhA46kzIz2SlJuDktMpOOzn4aEoYoRvibl1Fm05f4lyilPK9cMBvK9F3
8Uas1HjeT9yk1dA5XvGChj73xYCH+NCmaafzV1KO8ekeH9PmEeoujh5R7FM9us4SVxIUAA39lG9H
BKoZ5uG3vjoUqfipGj9SqEDxcQH7OLlj4BHG891xN58MX529d1EcauiYIQDdXiDM3viwlnj30hi2
1QG45EOoD4L3uex4S8NNA0gbueywo3VDGGu/BndZ5A6L9kS9f55YVaPRV8S+X+gs0BwoY+QQeA/s
eg3eD/wRW1icUQCK9y1jAlFkBuCaaFaucoQd4Z7p8zsj9Rd/veLpFWMni/STjsaMN+SQLAntpGHy
1bVEZyRtNciJ2iv5K/rM6BkRzzEujXCdBZx3cKpXIRuq73xLs5lUqg+b8LOBdb4rYV8ZdLMfu1Wt
/yAN5X7YMx64yyzOa+0t+wtJKNeoFhJqjKm5c1Oh574TDsmJf6Adf7QzL8oFAr2xCq1LZJgc+Jnz
mS6VRGhHZkKUYG/olzA6KdN1VKsKDXvZY5GzYmDzDomouDtjYSLnUREWat6LWloI2bGUq4I2SF11
r13UhG9uHxg/aJWzxXrvGnae6f73xU/9sozgA13ou7qbUta3tc/9tGcwq5D3lAy21euKGQWJg7Oo
uWJ6OGVSDpRQEeLUWZ1QOok9HkSlOh7w2akqvaljWjCT16j4fizp+B0wAaSSUbVh+7ySx+tEOvdq
rmnfHYsDzbAFAf0ZYbV+d4QCx6vGAXg0A0h/4aE+MXG/8JhUvVt1WQp+Vd0b3O68g00TyNN/H9G0
yOuXz4PcKiwl+6HuC4zPUgA+iy2rZDzO7TsW7njOt0bIavc1RTMGTVFvMoCE6a+ztEV2ZK2NOvt6
suholiUMT3+TZiLlTn4zX6h9h6HTUvYMPpYfmrxjoaPm9THj+uLBZuUJstaXjXGdCtQoV13zZ4+e
1u4ZzurBeFKApCvoalmQnqauDoEtrrE6EhaR8SaO+JtHgrGBd1AsOqAMLltGIWANmj2EpPQ8kZT1
Sv/xET/45C9P47ci05d7UnOaQmiY48IBnrvDDG2JdcNF23LDCWf0+fE/FQce88nAdVws+8rvweCd
JYwcePGgSeUityTa2pt/2WuUpiaWZL8ZbDk9w0BEtvCXCEZoAIqdg4PULoA8/tZnpTfBI2bVqUN1
nmJqYjC5UGH6/IkdlEz2iTlZD6kOUGVGWoOKAHMqO4KlWMNNjzkcYGIVBCu290KaY7xarYdhWDyn
s5+s/laOZYp3tpm3V4huCtt+y+YlISCceXb41p484F4zFzqSkK7oWcuLqMtCHZnO9YCRO4sMhyc6
hA5UDoMXs1UKJLAs7UNZEhBFctRmWkpNXfAhghVELrgXNzVl6bMoK5vFRo1RdYB1nrENl6+3+q27
GiwpiO7jkfOvM7xVREo0t17y2A2C6DMg8R9B3IJPkYlUcR3iOaff8SceZrfRcJ9tVFGQ5irOyGSf
OTMP7qt44g5E+GsfsksofCeNRzZ9wuhwlqrp4Lphn18DrFmMAm7pFwdXz5mXv5B7BuI3xOdU3a7G
3gVjTqH/Oz35BD4zedR5v2qvEMs84yRC0YVjUZWCdQ588lDXIeGZzOuAGOq8EVuSuxs0AlQzLGhn
iSqlW+RIMa/4SRzwZfLAQJJ/dgP9tDt7Y88pIZtbBulfnx3nW7t7xZ/ryLbToGc+EKNlR6BqQ7n/
j+6Zbt8eguTtLY3MtMs+qSMobDmbtDgxqz/I1dn559lfXegfizPJj7Y5PneAYoBp8Wzk6KfVqsJl
Q1wn6p1dbTz2mkP+fVAuJmU00RoXHymH+OrsSG0YxdFWCQvXD7FLg9XUfzyqF0sGnGsIq3lkgahQ
zV8W7TQsWVFVcqZkFdy2Hs61kVIp/EZ4VVInM6K6aVIMP4CR02wuKZVyvvohG/CkwwzZ2dD1AvJp
jZww6a4l+fGNmP9WzBBvzkr0hFly+0ns3gdyXk0ABEOfboFFVCr4KT4QsIOlph4prwKjitl5ntYF
UKlnVHEXLcD/zwR6mH630UI0XNruZC4Sky7XXxERoOgrCKKq2kTMSVnVa0xmSAPS8QmcoNaii5Zp
qdk6X2Lv6FFAKledBmGlEx3F9NAZap1SjLcvZZm/2QG8VX9zXjHncMZ4dnw8zAZ3uLbyypfBcOsb
3r4N5l79h+UE5qryaFNh0RFXJHJO/M9ZMoa+uNpC6SR1WSHtY0d5GTAgIWF6QtsgzgqKIu7AswrN
HBUzsqQ98v8lKdm6Nl80y9osbgRGCmsg0cg6Hw4H/Ghniv6OoiI+AoHd7k8bVv8UHPorlRjvOaWW
s5Vh3lPoDKTfsQMm5XrqIZAQtXNsjM+rReA82meUJJffOpdi1smFQCR1+eYWQvZh6VVYtrUuViyU
4ftDXqaFvHAZ8My3zZE196JPoGG6q/1sdGTe08bUeWhYo6qZnwoPilaIKYmwrgt5WuUto8NL9vBz
qOXj7thynA0u/xCwdMFjWu9WxoEJ/YuxcPlv0ghjZuoMyGcPEx4d+XdPBohXq2VkBNOX+OCXuOYJ
btt9qgo/HbuNWG5SajktgzdGa+1TktgZ47qbAcxRRNiyWz05vGq4FPU6zaRoP1chB7+LmB8iOOM1
1cxVVmYBsDcMsqOJJk/Kjfr0Fep1vH0o90PY7zukn3SqflkzNjyxgmu8HdO8rrOTmnzdhqglcDMo
tUrB6LTsphKhd3fAjpflOkMtLxBlhpKUvPCpl3y0Y3DzWjV47x+Gn28kZHuETBqRhdNr174qnGqU
PAyiTlTigISXeP6q2zNII7EMBAwq9RLguflRnJvFAuap9+VBQM6Az8+ilyQ3T0z2uUSlTxzMZhey
AlVKH7NaUE2hd9dF2i/mqB8nBnSucoBNGcZUHFvXni9xCmKWpRTdGW7QatFV3W4a+pawZWiVNQBf
bBeZpbBwq969OwzyYflrDTAlZY9D6i89Fdh8d1eROTOdGSLU/SO7ObIespCpT7mqnZs47eTY1pmn
YYFR7/ExYQ9Gv1tz1fapuVr8o3JTAL6t0/pSzcRz3lOJf9iJeakLUmjUxqbU2rXaS9R1rc/FSipJ
3tUXqcYWVsWv5zePUZWzinZcV+xPh+q17kiAz+H5VDO6GM/fFH18hxPcz/010eOYoiioPoTO6FTB
3WjLVf6BHkLfk4Ld9egUWmlShLhYPBTy5MtkkRbjdiXZvaoYgPuranu2nxUNoEi4JA5ijosAL9Z9
6oq0B0YX+JshiO5uHArNRhP69gyBHA+MxqfN2hZHxQJkP7av/HIKgrDkJpt/e52UoTif4RV1bYFm
Wu9b4VWgZN80ZMtyPAb7evxR5I9y0GkQfWnSRfljOmyJ6aR8emDu06v16mymS0BHXVZ7wtdZuJeu
u9zaxFbDehYuJekmX5HMKi3qD7ahu2zJ2qDL7Pj9xXy4W4yyDN0DZMrTdUu4tbM1tsG2osJxZrL4
CxlJL3N16XT6ZYVKcxnyzf4mC1IDAghhG8aMLzJCdWoylv7UXuJ0Pd5rKliDyDCCpNS/9IgOkYK+
T9w1TzJ62xmQalGMZ2ULhvbDWRXlBbiECxPPk3dASAmB4DBUaJuzvxXRP9H38NtWLX0j3PirjMMC
vV3mUvoO2qQQQJfJCA8zsy8EdcjoVxT76vSex9AbIzyroxkP6OoCmttBcAmzlSC2+doYnTYF1taJ
xfQA0aNJyjiEme+Dhnk1IjXPYmvyf8gUnpXnemCLlMip5v6Banc0+rVJM0p8BaO1ttK2TuD5iqHq
81xbvJeA1IJY5++lQIzEdm13mNS5q1jsFaz9bS2dH4JSNinEFJUf5D8pPPDpNOMaLurwr0S6IgTu
VW9fvh+uU8ptzYD4EVpbsfGvdshDuemR1QCMROfgdo8+TJxFWp2Vb2hZWOF6zHIyx/zwzZCeTg1W
t7JKOn05h6tHRj87TpfAq9QJurX2Irzti1btQ7bN/0YYkS7MCv0hPzvZwPGjHoaS4J98GyCGekXi
zmyE7eD4tw+oef0xnlsxRFbwRLT47/FwReLwON2oJME7vlPq+9eEiI4MU5e4sBOEdLsHO8CHErwS
9XBN0fXyTRguyxG262aFba1rtcQ+HV0T5yF/8fjFwlOdHiQd5AKNoK4MWpGTUlh+UIg/IkGund9E
z+jCP/qYUYib+InN5QUpxVWrWgdQS5+PBBsFxEc3PPRSm/cXVCDspHe/YpPxWWofbYjS9bbOuXjq
GqJWVXrhUATKyWHdn7ERIj4WjNkj7uk90fETObdxpjP/nZSSl1VY0nnx5+A+VjZ8Z2o7ek7BsaXQ
q13xpm6zB7f/Qvew/BOAaq1+yknuRqBKjKbaOMReofF+q6HvSVccCqKCKNDjEWle6mXw9R0AcoEI
e0UThEWJtVRSdDhnZpCmGf76pYzSLMLY/bkDBRQLDeH7ngoXcMqQV/UIPH68ImAlsh8hCxdjcwh3
FpArmWuth/4DTNP/ipSFAeLv5H9Rx5IAdh2kzJatlc3n5P2zJ6IWXkAeroxzDHxrC1Gc9cucd/hd
aV4DsTEqU8N99syOUgjNe+abJEcmOzk/+faMUCZtn9b17Gz3Xd8rAjRbP2h4ic4VDjQNrYQjptP7
8YyzgZ9mE4PxcIPMcW2gllmE6OU4589NcOJZQxEqddIlqbgkK5PV47MnRTOfG7LABQtYJilFr5bA
63ymiGcir47epMbpZbIEaUEVT3iTVdPEnsnPbEBCX5CMrOfNH5zNzQ0KUaJ128WHGVHIGuNjipYd
CD/zFg+FaW72Lx6oyZkCI7k1i1Uvqlpulgyfri1ay6UWubvCHGu+JIzITw1p3VNkwQbIaxlBXoVY
d3to1JTroFR6ecjIi0ostv3b86cWXs3PKunYG9A6pC9gdzM+dSeg8JrRO7n5XgdzRV06DD+l5EIr
1AyaqkfzROaRwq+toq8e5ZreedtVBUzFPzr+vbzqtsUubgSKSgk3igN2E+g98mVJoCoVciyOEMAx
IoNk/++A71PIfjG0aPIazn/TNYheADZHd3i0pDFSx5R1O9HfAWrQmd/YAzo7uW8WIkJAUywDFY1K
x9qmkP2ZqHpYlIEdImBApw2WiEGwVfg7+UomSVfmrJK73Y27ya6YC4bHAEF2giL+1LaBl0jxmoSm
ZKrdGKfAyqDN/MFaU0RU1TZdfROSqrEcfirM3QdrHx9HMmUZAw9WxZQMLS82IeNPmaRAjbbaT9+V
F9xzPgFJfsFXg6wf1AM3TLwh8B5Qb53BuEKHetSPIJc8ObRGVb1wBEIn7eJRQJ9oZyc9l2oaEYD9
mFToRMkfRHASGirVwtZglR58kuN1jwuY6cQp45jDfcbrl5wxahGbtlPho469wTbIa6wn59OQqTbX
3JxkQ90ZdXRYjVC9kl71EjGayXKZj7XfuzgaW6jrjZoV2YLEqibpHdzyV7vlAvFLKRVFPkhGJ9G5
/ca2nGbtXW7bC6dugrDWyXSWKWDBjsLygy+nOsIaTsyab3ygX1DAwLltfX/rQPYzdxpEypkxmPyq
NuQtDmZgWKZ0cvtYzohNN+dkvLiYuF6cfFxTFc9x+ndfgp6Ti3WxcLL+8JN61TMavI7IkWiexGIM
sLSAzxQPOzIaVA4+p8q0GgcLwJ83FDevtz5ii8NZocTbJ6402PbdaWJ34i/uQBPIrPdJ08r0s2bS
poY91iqRkuzvRwKc6fcE5hh4EGSU+HwsvFcdMWdAotpo74zAlAET/v8y33xSt+gvKKXZdQeeQE+t
IxSKcuQIx/3Z0y7MqH283sm3aYIr5z9KKS1Wesatj61P9pKf4JdwatXQsjJSBzA68232LXGfEUFZ
heXmz9ez8EJeSKvUykvYcQamfNC2j+bkJ/5aGoQicbt9UAaPPvU2gfXTxY6ICwo6tfTJPdLdujDr
hDkwMt4joYdqz0oKacfvdjUfg+T6z1mIM0TVwCFb3BgK3nMDwA9d3dpWgYuwpH08b6wQ4qF+mcfM
js+6Acdmf3VRpx8LAI7fw/ycPQjd+UO09T44iAxFMgFNJhUryh8d7Fo0H0GWAP8aMRxuV3kCLSjQ
hxdC6fhrMUg4P0X4CxXUcEzuhyQM2mPM3ciqXYSvXqmKLmD6syG9Agwn5hMlvFELL73ZY0LSub4+
bDITvmpmtADAJun3th6CnmrEUs20rPLLb63Uea/LJDwijNvHTYyhd67M2j2+HkzPZSnC/z7W0O10
MQHdStLe99o/MLHYmgCKACQIi0gxsrpJrZmVyGaxZCp+G2U1xSpMLV8yFE9X+xP/jzTPutXa9grc
FNFKEEoNTwQNNWVkvVRsfjd3epopwrQ1pKeGLqxrm9SGqQ9VDDxkDjymhBFJKNlI+E60W51eBGJk
0rFC8YNoAWdinDradh+YPxlG7cD70vhiZAoVNdhPIvnRLSbt2Z05hy4D/Kr+c03TwDuBVr+b5egp
rXvibUZW5fL/i5qTV2MhaSqoNo4qYqvhhKyUg69uK+qOmvY61BEMeZV8TZDT+WCxEKJ699LzO+Rv
j/ueYEZUNYllFc1XG6ZlXUNtkev177xmzDl7lcQpZVSsL4mBAEE/b1zV/yQKwD3Aanu2i3IOKDjM
TJkppqa8VLgrocUFvnkGTff/4yivxnGIB31peHyD4nm63FGortsSK98e++9nmEql1idK/yNQfmp1
jfidEz3cRafV/3boDNoFkmzfgj9DkErWlrA7TElQRoFILUD0R5/x75NjdwV+KHLbosnk1No/e4V7
xQk9lhY7FpEQQe6QvmPWXiT7xLGVMng5Hrn6P0+JcDOSV092vkaA3wSDU+OIkfqXLRwxUOIppd1q
PMYXTNRvsnapv7jfgt7huFcQzvCPY2zms3DidtdJBFuXA3Blzkb6R0jmUtulttUGQ2RIHirGzT9p
34bsrT/hEoSRVxKq+V27yAwEIzG/BvQ8VhL205EqpnGaerhpFFBQUXScgGQ240HeAUJcn6mUw9io
lso8RR79t2fh7TOt1eHOFeg064V3uwAQQSRSxS6QpUxuWG+2DM8/sN5b/GOAovehIfgUFXIpnNjH
ChKrS1DE4hWBRXZNidCZ2azBfE9jRxvmqkiKRIl02R/+VdwV1ciV/YnAwHmWce3IvY0mT32ckpWp
6C0t/J4sUtpmylyX9vPWxaNxo85B/9Ud4SXkbB3g8UZD4COHPwwCmWy8X+FTOW25/Co8B9dsvnhr
NKEFwv4RywHU+OzzQdy6Pgb30hTjYS3jw5JkwgU1UpuRTdOrp2GYSC2CCpOrGAzxi2o/mrqHV/r9
gIoqswMMth52XfRdhkCshwkvk3QDDBJFkXhsIPUcrexNhE5dK/H1H9VwhZaLpBaRQLJtxUPROz0y
6dl4yGFwh0fe0U3SpefPI64I3xKga2DjOQsAdK1w39R7oJfMbgMayWU5Jb363LLcta1VBjXXEYan
+cPjjwkcDXYdkiJXcx20mf7ltuu03DgY21jdO4eQAxzvhhcvCkgzbMvvVDTirH0sQerQXaxrVw1Z
+pSlpJxdal3FMMf4R8CGMOH3WyAWoDIboQ1hGrpUDGsD9ly5tgpjZJ654RFlz5DC3L68tvGSYZ64
kJTfsEjjOcfK5oCsTNnnVgpf0X9EZ2JXmvbSxap4gPS8i/kwlmGB4e5gfhGWQ12oPB/WYRWSZ13Z
o+pOreUTUdaYQCTsEv7+5I4pT5mH3WsPykVuSgBG3DJOUy3URTpAmZ7CVYAIXgD/kHwVxHTRSz8n
RzRimwfnVZvT+sTn58CpIOj0gqy+dCNqIt+C0Mag514mCtl6bY7So/B2vpriHrTJHE2t6r9YiUQ+
HZG2/7E6TDp4pJTreP+i+d7iYBoYMhTvqYmiydzg0DD4sCuK5L2wM+FSgL7kilq8PupFQ0yoc/6I
yF7YmE7Wt38Ylx/G1EoNzvTjfoVOSa2qYMRUJ6ed2CgjkXKKmOcCAvjqnjDsN4/kjQsnva4u/Ilq
35P0bZQ/19O6oU0IPVyle7VgfRuc9mBnIx3U3DAkfjZQJ4Nnc24tz16B2fH5lVU0sl0C6fAL3wNY
HJ7ByjI/G+SRRLHz1Qkgs80xUNn/tdlrS12E9NVUUbg1DH4FNFzaVr/zGdKiWvBrcPcJIgsp8rXe
oA6uFV24JGbwHvfbbNzz+Hm4ZxxD2CzmYpRuZN7DLio1XFwt8K4VcSMDJ9E5V2lIqix0B+qVL6MA
SU0awE/wp3PO5/oRWgVOjbs4lD2kF4o6V2vHLPYbQ/SUaSose/beSZPZIUhSxlxndwt9vErd3NJ+
gsc/U+ptgM3HrrRMUK1S7oHnhZ0+Ru2XdRCTEtb/i3Y83Jca5MW6nT5iXc11RimiZIwfoURBD3ou
rjHVEUpKN/1Za5mVue1olZDnUW6FQBCGwCKHe17GA1C0hokycHao9it4l14I0TGVatMHqVEI/Yjh
k0ZM/OgUCAw/mpTOIiO1eCCt8fZOtndXadD4SbIOki76Ory1dpwy8yD1C2tmqgLHYrERGn0+QoVY
rNoA4efocZlV1JhYlg+w4AIquvTaVpCmId+WzHwzBUIPVfmJFMfeeXPtgqjNxtrBxxxMuTE78UDi
vyM4VXcq3asOL/VlaCl1JEiU5zKyw8l2kA6bqPhdI8XOKaHOT4OrJJTEtYvt6K/qzl4uzOxG1J+W
yUir2VjnGyPMraQWZZ4hWfnhobCMoIl6HEap7JXGZEmVdYE62eaX3txxPpB2a9u77Vk4UqRFiQkM
L/z64TB4/RcsBpLxqJpkACjtxCOGPPx5m0puWtWlCpbQ5YMYxCr8RJIuFfZc32ZFNdl6dTrT+/a6
WoXrl980rbrXtR82TWTbvTL99lTFVfEzJwq3Gr4+6YUzj+cMmWps2T+WYpl3Kd7HjEP2Sw2Lwgu2
ZcqyxJgT2Kjgt3cdUO3zOv6RgwlLMAuRSVy0Tx1uQGqnNSr1eVbJI3MJqR6AAZ/arvuyBCxVvm3Z
2/0pnsNWXA10lcMhezvNeReTG7Fz9kdORPgA7PEGr0wQofFb/Rdj+nKrhK111ccmqFwgCY7Vq4vz
VLNg8UkHypbMXEgjz4Rbe14w5QSDZ0TcXkq2h/vRJ81DbGVsNE793UAuJ/XbKS5Tnu9n5aXtGtH6
mqn07Io4A9j4RmpZPRv/+eOh7UHBK+8BIff4nkn5yBeDG/kzD1I0AOQUaPqRD3OYVrZ0mJs6JKK+
BA7D6BI7zLrSfhOchG2zncoHFkHbZGyjLpjCovwRc8i2DXaSDppr2BSvMhMCb1NvQ48spXoWbZJl
SCVhIV/FrE0DZTU+azGiCEnhDngZbjJ8Zs6rbGiqTBHH5y42cOMghykS4vxrrWa786Poao4nFj3r
vKvY9+BilngS2V0KfKjrNRHx+X7EFGBtDnc8OkNbL2h0IAGVLvcZVe+bXmtbpXINqLNB3B+s8Lcr
CLl3PrqhY8D93S59ZGeir31F8yGXg7M9aloGwyPF8j3CJ5kRP2FpFSu63FP8zoYhXxV0M3kbbK6G
xmszFkK2qpaXa9Y4iX97G+d9eP6Nsw5SDHJZ21xJgzfsRqQ3BQ1Eu011Z8tlu0KsfkqarwVLEMJi
UBuzcLjy2bpONadRqGkZ+eCSxpt1XSKp7dultPDSmxNkQxJDjeaar9WYLbBiJypQtTeLWkzGonxE
xWL8ACZRU8QOrmScIRClAB7bYdoOZylIJEPdpXLeaTM5237ZJ4SWaBGvWExnuG5q7Xmpii41XesZ
4JPAFoRuAINifozW9XySb6bepjDZ28knPU9Ay808URp22AVVHWcuaB88OJNY9gnLqCW3mxWdJb4j
eCElboy7J3YDVuV894XFyGxYEM1aHnUzP5MF+szr6kqrFPPB8CTRh2skGH37KjHhRBJYhzRZoENR
Q8+dBtAmjYfHc2to9Ij81OzQb1pnTZd6mI/4Pw0Pb98Pb7Wz+eBwY+tJrWFxIY4Ghj1RsXbdEr0d
GwAGivk2emuPky4bmrA0YvjsgIb3BjfR+fHAVYx21nqMDFz6xHLA2lF6uuo9tCUxZqAVX+xcAkNi
0ngxGHMQQqn1l4k18N2d5/2w1Agi+hrZUuNjCd1FdZG/7S1suz/hLtDIxpbBd6lPBK+2NRXAht4n
pkn+24cAXjI/tvk6HgVj4j+Z+BeR5rVkP9B0G7tfxDTrBey+cXqgw+GX52dGtTmMH4+y0bPyjcdv
mT2KBF6R2Tys6q/1I+sEtUycdi6jQwAJQBtDlHLN0IBBCiliKpKwnqvVv0wKKanCGHYnR1o2cjc1
gHm7gFy+FbfDcS0z6UhykcjEyWZo16dHOVHT3q/PXqDwBrpzlR7petPIxqmwfbAPzYuuV9jcO9hG
rGxgzNxx6KtMrgcuvc/zXT+qww5O2/refCYg3C4cstbwlpZLovWnSCbTi/OsN22hNxNk7gT0XSl1
DpEF2f5O9aBFO5uC1e8JqQiKmhCsImTfULtMgSM3o0maOwrKrjBDdSSarfKyalUWOYduxwBzh8Ar
ekyjBmU1AEwC8BkHtLBrZ53oabWVxdge47gKy2aExDsaQPvE+gSfH8gTDJaPN7B9axqqh7k8sQWg
QVF4zX7cSThuEaQqiJd39iMAjpNtAoNgm9+S4wsKaULsCnp4OkfmQ/nI9Ux+RDuESGG/Ib4TnBLs
mM4aUpBCbXwXr/K0+3b3U30dU1Rvxn/lUG8TkoLSP8Sp94LwtrLFZAl7NT8Mv6aDT8+vT98TNbiz
V1qkivPhwXljArIS4eP/AKydqX6rjc9kfWzGoLjGDy0Vl0HmMG3cmL9jW9VM/IuWlr/j6N4oOc/Y
PDMzxOGDzjk/e847Q58CDaWh5Fr1Qs/DJ0dk0ONvl9VuHC02tYgbwugT5KTsx9aSiDouB03iluWV
b2q3x/4mwAByqJaxIF4WrtU54v+Nv5nMmhkAKUgQB/Y3ulP2rWhLxZ+2W+wTbR0fIpZ4OUDSXQjC
IpL8SnN0fMj+XWHoy6lL9Kpm5WKAFplwVLakCFn++Gsa0ljqWM7fzWtfj24rkTqLFD7zf+N8S2vS
2/v43YGV86RzG4RfODy5Ionn4G6t0ISfvRMBNz/R9T+06vKKE721Jpmm+D+gvLp7yGvWqgO0dYy5
4MmFihDQwYpHfPIMfm0ktroRrX+z5C9cmSAbesa96VrlPGzJKu05rW3RPYBM72H/08ZZci0XhrTH
IVPOg25QuiMXtWaMtgdcPgVQeelhNS9gNxrP19cV2GRECLAHQ9fqMrUjrqC40oMde9CUOLcwnHHE
hIpzZNYTUHK0keNrL4c5Y3fHsoKXYSOnZcjnm1Sb7HwAr8q7E8y2RPhouOvgd/FIbW/dfse8hmuJ
+vfuDSSoiMgkEzwiCAx1k8gSzr6Y457ooYod2AToiZcdebUp9JLkagPeJtsFPeRY6ldItaUQqSUG
K8ljtAAuwbD+Gaa1Qnn5XqXqqmeSK8QFTazzI1I+HjQTLH+Z9HkGYrqVnIeU0lGCiy91Uffo4BYZ
9t1/6gUcJCgb9qDvrgSrJRj6gPKvCNXxvOLpkrB4x3R/LeXbxDuUw1jTXuqzJ0tOCMsZvWvchVAP
K0ut8Eg6JI7Z8mbVxkI2mXf/nmSoRjWUc7g/i7mByNaDVsN7xcARkYNvWMcQ3KRL4CtLIbjVLY0B
EQNMdldQhNGjdUunzks0GQ+hCZZH2PTtd9d2aeoyEOzehS3pxEOonNsYlQD7qrU8TSfTpJWkDKDV
sqm8YHo/l4jxGNf+GthYpz91ca1kADrxj2mvGwjXwQTZdUXhUiZzonYDYqy3EWW3dxhM51qa0Eay
mxZ6fUn+YBRjRdpPCBvUbR07X0Ka8K7xEDpSWqpAc/d7Ebc9Q+z89VE7JYPE3138hwh4mcw+Y/k7
D+8FV8KGgx7Oc46mpb/fs+VKx2tIamQavLtMltjyDBzTDCNShUlfULXBp+I4qG/22kfG1U8eEHLA
XK9fsya8tzclODiPZLBFXDYfLoOmgN80i3DROWixJW4t+QzBL+smEqL1lcdKVfmL/YhkYffOikB4
y/iwuxQ7jaIMpOphPfn+SH39FX6AGPxwH5NUBTQ6S2NrcHFAJDTT37eLK8t6vXr6xtYHguTohzXk
sTzYp+bcL59B+1xlRRtut/K7LFE+8kydA9ies+cwQnflk7L4K9FDOSTZ/tzEpEdO62r8KxJFByoe
/Skob2URpLxOE0eTJpgBWgKTRoOu3zEXKGMi48zTHivp3CpitoXjkAWmYoU4HCxQV/Raz/F2QAQp
fraVjXYTE4axqqaWPGXIg66SyiHcYMnoWkd8+HGRFP1Tok26FNSvUAVxzRIpBFnY/vogPOYytxN+
hMLUszJ+vL1hDpt8DVaH+3vRkEGdOV1lv4MMwf3G12T6xtBarMYH22LH6bcAerm/dZWakNBnuWal
NDpaVJZ9p7n1XH5JljfP3J5z5STtIThD4WgcftlDGivUanVQxoYPttq6Ud6iQOVT3MMm6IzPJKH0
Khueew4EuSESQ9f874yxFWKyvEQWj7MtJU50PfGPy1LXeNyyj7+XbdOvSjGz4Yq2BsbUuyyEgIoF
Ih5uaSkh5ct9PFYrh2YgmoqgL8Ko25mvFtNJgaIHZYyndaNzxoGVVUb19M1L8rzdWzoYjPXn8X+U
zqmkAa/ZFqSNPh0EQLzFifGfk9tI0Sc8KFNC8lXdpn6tMlHBR76Z3a6DH++H+D+FL85IqgPjccMV
kS60G/gNUFapYPcJQWDEWa8usWyVnP4auEuy+BjHPO2OdDl/uUCVuQjNzizB23K1puLe93Kn8/6a
GqYnS1QGLMepreh/Omtfp9FFL2GWTFt3ptzM/HU98UQDLv4qYpKIhMkfyGBHtjAGWbngtCb1bLZG
AnxNki4wzrhsJUPn+LyvPbCqZtAe0nIRcZSQcObIh1PhxHrhVmybHom1wP68RtyM2vwzwZeIivDM
srbHFPR3/Q0ic3ZaShNvA+dKGWMmkOcbfLnvt1KHinZ04TJ9nO0z4FmGt3n22x96OIMQp2zca+0I
XnemsKeU8mz5sMBGTP2HjgdQZVYdoRI6T9XWZKDWlw05rrV6aL0u6NLupG7jS5XP1bLW6NIwTq9O
dfUjdPauT6LXGuYR7O1p3bN0KLLLKor/j+k7Qz1a1AEEUuEiGw8ZKekqPlNqMMkuCGott7EqwqDK
7lLBLCBZNNuBJkwW0//8WU/bhsiJh/iFIGllTlKZFy1dEmdZmW8bjy0nNcc6VtwMzCSd7x2loVaC
lf3Z5vpg+41IXZOS5Z9LbyKUaEBmGubHaNoZ0NWzxfzipxKF9zDWXlihHBtdUebqbyu1hOHd4341
8FrE25zS4Vf8lxhI/YNJkOuGn4xZLhzbwvbrAOKK+83AeD4ZsaGmefNXoBNvQUkhZenO/Wxt0NPO
H8/ZoFQruxn3r2o3D/QVIRqciGvz5R6DeN8g/j2koypBbBaXlAQRlg+GUKpnw7ZpPksYKDsHXwPf
ZooF9tDCq9YUYt7dp+1Ueue5m30hi/BWRABdt5Dx3QFp0Rvw7Xcj/ZRExvcytQwJGDA45z7v5qtz
dnAiu1IRc1SihOHEc9IBIBezE6NOHtNbD6gQ50hVUd1yQ0F4EWghyUVp4imAYqRgofeEGjCfd3hI
Wqr33vpUcQVGLfaPpIMiyefcjr3zAcGJWg9mamJnRI1y4jN8mS0dxRNu0hke5RHNgwrp1pwMUjMk
VplRurXHwq0dm7qO3pTNWKCBpXFKpcQmgjICvtPftueLL6NycAxXcCyPupSt8fAD30areDFagOZi
CKAwVvoSApIHLzfizi4NxeeYrOKs4CUE0fG1FLr88EgYBD5mPK414vTcPyqirao7f+dFaEk1AEH9
qi+O66exB4+0JL8+yUdBk4Xp0K08MVUoe4lqJXB5pLYg8CTpjpLatbLyXH+tUgh0Q0StjOZlSoz0
ZkZTaqdtPcK3Z4MKpMpLmrbhzpfwQp+0QO6shJfIvmgh9Us67dTTPENQAWRRt8Qo0m/UyDEp2W7P
2thTPxkFvuwg4nBYSeLDbZ6qSSK/+xl3fhwXmsEkVfaPQjrVZfNcRNKcGO69HLIJM+01/FFiedzN
//VsqktGMswQo3Xi5QrTTkK6IzDgKz73+2cAqi3i7s7Rb93JKfg7Gy93mvrQeEo5hYZRN+raTyfD
FDzwz7cUSTf7qo8C5GWDKsRYxjoeSAbIaEJ4rFU5BhIHATJdlDGzIfloTEwz6NECe3FtMYGksXxh
lU1v5IgkkW6ghzN5PmgdDvfNqgofD535mTosQ0dH+E8075PIfEzxuzePUziAGDyOoYHzcBLiTQEd
5EUMh8IYawNFMVKEzLFAf0G+ahY79533/UKXeqf7jhycyP1yAWGb+/qMnJtyOCOycH8WwvMCOLTA
WQovCmFgAN4a7YzElysSImIyqaPzwwNtfwnY6x4LxORzN54I836TO/8DKb+fFldm38BhVRiDFK6U
4I7T5/yNQigTpLWK/wgkO/E1SqbrxH8J1tSPEQgjCqc6lTdC5odC9q9k5JgaLCvhxg9Cp55tj111
04USwZ8cpVhX/Da5mDm2JMWNG2KV5a4qj1V8d46m9o4/m3EGKaiBXxHzxb3//jkJJWY8NKDGAkKp
hpYZI0YoncxBW715uK0g83gHKXvEdF6gIt3iMoEAQrM2dYLY5n984UFLI5Q5lq9iJjD47UtRl9Pt
5N5Ja8qGIszCX/v9UdvKtHpbXePVDC0HzuPlECI2ChMy30Woh4FDmEVm9Ha1kVEgrY05kZHF1Yor
c1M7IBo5Ha+2q4SQYg1s632APuJkfvuzmTMAAkKnIWwyvmqv/CX5XnAHrS8KhwNoAbC/xIFTGt9L
q68+7607Oe+GNZA24iu0PQzhZEr47m5biOSeE8VFATSMHAR2T8VO0I6jBJmhSe+D9WrE4zTIVLmS
8oVHgrONSfX+C5LkyJuO40JB+DjKiEMKR1xjnLktHDOAsYRuABDHyd8PI1BlBFuSsby9q8kP3rzN
KQx9Y/7dRXGR6PEp+q/0R5cIa0TaoChArWEzt+ldqGGMXyGkPz43VZW3SAfPjPoWQA6ikvAC8LYm
EntudiBaB8d8NZhjHDB+qxrLSatPjI1C1d3CaWBvwdZ/f4NDstvL1gffJ56Pq063TmfqGmbnwvCA
9Esg+2RLZ2gYuNUfXJlLUa/L7t3KiInEGh3KZcLlGuldh3ylRbA8oM0nwdJVNGIohBfNBNNUpu6j
iuaz08/3RqpT9SpIRrXn7I4TKOf+5rrcSwUr0kwSpNxCjo0VdS9GVV8ICvVQTonBGDHSXca4XVYD
4Kk7zf44R74dzL4Fu4ixLj/L5eBalrSucSXYVXxlv091bHz/e7D2NNhcZG2kZd/6JtyCLtT9OgFF
11AtmZsxZDk+13DgVjAZqbc1AcKc31mnCpfYalTpphfUgTxS6sNKqco2Km5Kk+sMs6OHgWmrJWGA
LINvPau/vjSOhrNNaPdLurGXgOsSF5E7LraTsFxsoqa9/2jVQk7B7v6ccHz86gMU2G+AiLm+GuKQ
jx74nOwRFvF77TZDKwUIapMd0CnPcfkV8RUEpIPDncIhevX9BJBKzjjQVYdFaZmV/+9ev3wUDSJC
LiyujWnBXTApyNcAvrLwXYYhU1owsL1MYtlroJW2pV3YVo0sDlG1ZCTQQO/E8IPlAGsO+K3q0q9j
ZKTHIiuzsaGPbvOJ3YL9gevWs2PbztXEBgtXhXVIMFNgIQEzcKJItUjjexSLGNhyyyWaEEuI6iet
kQI3X12jN0xoWr0QzOTL5hsICaEmSv251SE5MSz5K1t68vP3b4tYtB4TlTytBuY6Ncrlom4bnnnN
8L8vmd/oVL8likM7blxbaXx++bUzhZmcPx6IpwtxI5Tc3+rAK5fnMhWp3L5FgEasHu4alonrfkYm
tNvFJ0hacta0upTOCRKKuZ+HLvucMV/Dh/z/V3mjXr0OF3U5rEVAb/wVMWXORWaP9CkjBbxjzQUD
8iI0x67FWeDizLrFBlVUEO3ZgOpQLfk31yHwe56AHqY38pC2Jydkf9mOZ64hVjyyPnd1Zf3CTbmo
HcbJaSWHe8ntDgZaSbW00NVbWGlh5qUmx6u9IJb1DXHx8/LrMsJj9WlIO2/SlPfDQ/wPKbT/bDqR
6FeRsCpLGgbhl/yHdn4Mo8tID1s+LZltMJgRlT4py2s235sL+I2h/1by/Xy79TIYINJoHxZ3uNxD
9f0WtAmpMe034ojniHH5w0SoOMVMCoDsa1b6HD5dLRTMPJSZeb07ftRrEZKFIJ0X0lssa3DIxsDP
/wqAZQsQMXKRXLXMfX2BVHa07IC0jizhEZiWTBQ27BGDsZaT5CBSi/LaKsCQlB01i6iuA+a1GEYK
2AeNpv0VXQUA9XOlr3s1hG5Qxue5ktnStAgnGQRY8ZFzm7AIdHcRDuOiWSY0ifJJ9ar+DYoS5fLf
d6sC1ojWiLr31aLJEdEE36q5sjHO5X2UF0JSa8NdSExFU74p5ttHDQuwGSUbdF6JqxvQXQSeOeB2
tElCB3MdZ7py0tThOHDm6QMk+09LKfQ4IzhxM/IOT7lpeMFdxtpxHIvAa+nXvVoM3q8uTHm/Akmq
8snh/QJOXnEFF/hQLG7DWR6f2+qmYnvELaIOxiWw5D9dKBvzFVAAIRjxVl17eDuhEfBWh66xHZkT
1jrRvdnEAhA2PYpdaunwCOlKDo0r6uhxKdQCZ8gff5l+fhXJBE3s90lz6N5cwXSuR8CmJKYl9Wp0
vtW4i2uufJU8h+GiVARxbr2PRkIggmnJDP1K9mcAVj5ulTMblwYpUe1erL1h7cKqLL26cJd1FN/L
9cQlG2he/S8oJIHVi3mJ5nNmRr/EzLQ5mzvmK/Yc0I2YymELNCkHOeyvLXgcf8+v+XKRPWGHQzga
b9WBI9kkt6y0Z7EAkDHVOrP5A+cBd6+Swl+ENFTFNhe3llv988lbpidJkbDYSimhUHwKjt0QIZp7
Clba5iC+nlhnLOaqxbNU79imCHjkOlFeP5opVmUjdXGeTs/TV3UMIrD2jdYC23YdPvpvs3UhLJnn
3D4nqYFn8h/dPK317xr5rKOVgINN5gxgSBrXwb8iSse8zIrDD80A0+3SWoZM1eb0wBNZjAl6euC0
uz1daQ9TBEEWAmGivI0OwaxvFELQF2k+23rIYnpX5sFucNJ2KdSFLu4LkUIiq4Rg6+Mab9lUdKSJ
RqejKsb9EXmfW2S7Jml34QJnSLzbwPsgNcIrglUZ9e2LoTK7u6sHty2u3PkiXpzjAQvZjf7R5Ul1
zq+AN1ktpHLSpTbvvFIiqAhPfoQyDmPdfUfFbqCXze23W2RHVAJKW+DOgV91U7nlzd2quraVamjC
Q/bK1pyH0GwQtfU437LlZ3ro+RKUIS+joA8bY/Z9lLCGYIqZgFIbBjBqhdEUxNHlGgqCTfZWdGWe
C/qK3FbcOpcWlUOlX1jCKDEQGeCLMhmBXCKFPR4mlbfddosMKLJ96pQFvkk6jG1sPbLncILSrBRK
atjgT7bYQrSEzDM1EMME2x2J6rv4xUhq8WvwPs8IsKVE4I9FHE1BGpQMO0AztZ+Z1oiUw8QVOIhL
C6aIdxdQKuMDJwRaVm6qm3MAiCxTw9rKvdM5OyMrKR7Ua9UBV3z8cBcAGj92neXVaZE23CZhuVT5
qOpeN7usXDzRcBvMT7osbish5QU3cTlodVRJqeV5ODR+Ncfu+w03yLiO4Q/8HT9BtayyTB+MUDAY
fbjGUzww2vVfyXYMdR/b/Y9ZP5jSFpWRIFbifUur78PLckRl0qqBcVqa3kcZtegGqZkzDAv5whaD
STlnaVJ0puRopVDQsojR3uWK1XcXokD+hRN7M7IBMdtQFhoqJMhhseASMFbw3W8dPgPePLvGB8G3
bfhU8YqLZSqk99yqYrBtlckJiSeVy5F7fAPOQ1WVqsljaQrWRD3bwzPe/W5wdVWDjoTnLdYC5Wt9
YBXINKs6eMM3jOW3Jz+bddE5iQWEnd8OpLwzQrvS+rHSYNP4IOcZrXOy8CcaA3zsDYYpYgLyTfJv
YnqP56HTsrGptThHPxzSdS2AQMs0h/kTjv+/2Ago9ZCn3xutbH8R6eERjrMy8+pU3dKd8xzH7uR/
huhJUe5rptdyJcUL6JxvmB887dKaOkS2qSv5EQTE0WG3jTiI5zYEmjPGDK+Lcc+IBsd6Wv54TaIo
bdozlY13PDnLKj7Nmik1nbwT9QQt3DP07TqxCcHBLHfkmEo27HlNVr3RSQ0IKE/KX7+irJtI2iZz
n6DXbxzi1BAKGxcPvasTZkRP6zxA8ZwUdVqjnQwIQp0ckH4rRDbps5/GkdVVdMOeOmqidFeQTfob
5XltE19vtnQzkyd+BtI+WgecN36HCSD9LAFfwGddlgkgjdxjBO1KWwxm1A1xGnW9H6etjp1DVoNV
QTdnZLOFpSBDeKleo+l96P6i1dvdkFHVwEAoPgdnMzFff+U8ctZKJlMqu8Jy5ZQzr6PcNSPqJrzX
jUEkm7LQr+20GfJT69RjVSZpd+R4ZGKxv5abmz2A+d2IPs8nMzu7D54t/LOO5lEmz5jzp5+q1n8J
i5CR5I//tcGWb634U4pmMgOHIMPeqa4GnPkRZA+Ruf6TuxCJSMi/D7nbCnb7C6zJBY6HX+bLGOBq
byx6uKuE5aIvRMmhpHH7kUa8EPojhpreYvteFR8cH7ygp6kQ9FJu3cCo7IphZgdlVHbASeFrUKKi
YBG6C22ERN8lm+/YooHUuAM2af4pSp0C2gUvXP/FyS/Fgx/lcmoMGxVRFjVinCdEgtJuwETCc/Bn
pJ+ryeR6195tO/6BojVbDsyyAiXQx7tzoms4LPg4nVZv6HcBsgv9rvkkhHGGYHKvM0JO78+iP2DB
9vPO5KwgNZF4hfp2EWgZkSgFTQpIfnZDDRVhkMNefAsZBXzppFKt4ZjJGjVtpB9qg3JuGLkMX3Ed
StG3YlRxgJQYM3v4u8D4nn6OL0oirS7FfQQpt7mGqsx3CfWbd+c0QiGNNf6kAKVrYLoc7/mQJNns
M19xBEBKrWsHR+etq/+wRftF+hTYt0WuZHf7mM2FvcPZVNw/sA9cd+sfhKj/U7995lMzMsVeodCr
RZ5i2eHY3rSnm9XtxiuqbaWMITyTmTNAK1Y5oj/VlojPqYYpPZZS+bO1xM4nDcLC6VLL0Qqyh7FR
NGF/jl72iieMobjJiVeeo5rNfkALUL6vbm3W4oz7fTKJhFvYvSb9v2OEwMZ9Ck04Ne3VdMlVgQH/
7RfzEg1DY+D+KvFBPxAWHZmYX+jlfnfa3FztL3TJOgRhwAzyNXDPmsBicFZ6O4fgCFrY/41XJpn/
tNE2KTND5ihvbEcakHzU8km4OG7iPGfVXV66c0dHTI3Bo6lJBmplM1g/MB5xAHfDg4WFNrHuRIg9
ww/4a6iUSvYELSEA+6xeWMKZb8PVeFcPHa24FxXr8eatPCm0A5qpXnmP/Wchv4FKlAoMKmpV4+v8
y9YQ24DH6WZT9YbIfNSN6O4SVizRlc41BdU44kdIFHmE1Xj+6/HUTsJdk78lRL3NdmGN96CwtTJc
sYqlzkcIyzmttVVUWpu07NuQu9je3Iwrohb7U69fIETDujmRDiuHhOw7zlzwP96fiUfkxLxa6X+e
UkXXs2FVJkMTMr7Lb7OMUFSj67mgDIa83UPD0km1WxGlsesyZ+nrrHEckr2dXqd2NTzvbb6GBvTs
Cr3zkHMKs3JHlnmkoz+pH/TVExYV/aTLm+USwPRoXHiDdprcQsTjGSnPTyeZRJTnO7ut0y+uyK9i
lPKOa4dP27KsVtPwWZvtUcndr5b/ihRixZfg9SIbITkRq+gne1gVCp3FhXqDBdo7TLsqPBdW6NHc
6jqKklfQ0eEGaGqJG97+vVEoCzIbkgoedkHPaMgouB4EkifsaeRMjZyJV/pj0Y43Y1au8ENdHjjJ
yYrwz/gGm51x7Kd2v4hl0Jg/uFbhmKHUAKQ4cyuh8m7KPhBUjYeUNdHpZZniqM84R2KU1FEn6ep2
1L6Fbn9yr1Z3fGDNovtAtEsiVrxF4GlygjRnfTNvDf3PEJt/y9sTKeOFyT0qmvl/GCsZmKJYJK9H
6HXOOBocqtThjzOKLnZd6ZXIZFZ9U4K/G1TGQcEyCsoV4bU34Hm2jdZAYGwOChKki7zkJ0PikxiS
QdSQNWLSsAhYvd6BC8pgYo/RLzOMlbbynJjXvcFhViqbOhkpJrwI50iLuGGfZtm04x8DDNOppLuv
J5hiH5Z/u6QxhHOnPspyIiVRv4RI1e/AXp5c14toB0ftRALyTlpHZCoFa3IqHKIxCUgUpKkAZ0uX
6OthnWXTEwT2d5qEghzUtwqEduS/MPeRL7Lem4AYHE2SigzNq2sINCjNQZVv3+zuJozcsYj9zjpz
VS21ot15LH7uH228eE1gwlYRi6tlYIcPuoYM2t/IuQxk5ZwDNofeMOq8ttCfJJvAGp28FgZstJ2y
wwXov43MNUNK6gJSDDAxTq+7MKOKoZaNJ32yMTi3zt3sWLs+H+2/mSBvBOoKMO6x/l+/LO+0JsQZ
icMvKbDqdKGKLTkkk9bglOyoSnJ0sSLQbbp80PRwaLhM63hacOIjGBTmXXiM9OXeizl0wZ5kdTLv
hTlNR/lqlycHgSSneHH1aaCssvvjTHMuPLw3FsLf77B/lpkOVKHvE3Eq6CRZf66Kp7bOpDDIK/1b
oVKoPuPG16XJHUO2b38KviHN+RaM5Gl0F/29sgprBGbwzDRhQn1ibQF9Cq6Z9oSrV0fdxe0pPSQX
ZIIHWigFuGWHmHkucXE9OiMNreClad6cfrkNBEWM0lSlefgQPxrY3zIk+qv3WrOQKrb89fS20dRl
xxb74wO72o/XACjxiynCMXq//pDOAv548/TgRkcpDWoPIeNad7eDsDaup8G56oN4RIlVoqxfLyYz
ug4hXT0HPtQXe/dst2PoSEORqh5YMDodeUbmvsQ/KHERtvo7bRo5MXoDa4dr5fUm6+tO9qGRVU+K
LXzDo8nXPgyPzIyuoCp6EQP1oL5T6yy+MSgTX0/N8gjqm96zKKLr16NhuX99EmBz9Jrra9voXG20
/fRO7z/cmAnLiQ2ISiKTq1PUs54RC6YE+L78g9B9oDC3sal+E+VentcpMwiXoZ5GW1VaFxlUoU2x
HjADDoJEGTxxiEshQxZZm5/ISTRx+l3s5MAi/1jwxHV3l/JKyAQ4S8fGzju1fFMB6Y2GjqbgSdmR
ctyT5t12ZVYzceG89dSOJ+cQYaJZT3mPyalVQ9tspVZBJAcyRmpIX3ADl8VFfK4aFNXbObyk3+M6
0AZwmtl6eyJ5Ei6ikDIqYPjw+E0dsO+xYyJNUv+NEZKD8SwkfGM9M/Zh+rpd/QEMd0TjGgkI8tXW
cOeVfeG4Uxj7fsM/H9zPJjXBZf3SilCtOrIti/VR7Ag7NgdLwdXHStiT7IkJ/bQYPW9eITqbzTU+
OqldcJVuTRTuhDpzdksVQOsc6dEPlEPkLinBmtyRbqQ2asVisgvsmdj6ifoqYGRRPHqlmQpAEinl
ipnLtctOVLFdB+f0PGZW+c6DLLIXLwZ+Bfh9SFTAL32nqSCYpSmtRRwpUn2axjw6yNwMY5i+xWOw
v5Taa/6dEHe3DjqGre1oH5Jg22naslGMGhT09XQmLlVoq3QEUaqph0g4vT2FHhwuPf20ff4pX5n5
emYkQuzvlB3J1AxCRSMpgn4XX0obaKGntMI6gJcMIn1oQEvIkRHHadkuxrPQrNyhozPqAS84yfX4
5GdafnIoQjbs1hic5ItAbcjEttGSoFi2M1aCESK76KMXAmUJxdyeeCGUgkxspuo8ARs61ENBlxe+
6jP337t9lfF4NzB6No9FH/62S3t4qRvkqF2JN3w0tWhduSb+MHehatXeRJJpDkoh0a5MFLVDC1F9
iCkiIjrCT0x6PLbKOD5A0Q3yvU0RyAW5ECMdmwsx8jdhUdfSzr5+RSV5UynFH3UXpQLURIGxAnlR
Ep/Bhw5L/KScL4arMF1miwdCage1XBuKO98kLzJCm+tjibeLl1cR9A+gIQ4Dt2ksYGCBxFN3Ti+/
Y7R9sbTgS6vlVHk5xiop3lrC5rRnbS6bfdjCM9qt3TNWGLdsmyaII877Imm/NLuTPDhU4C/qlwW8
GbyrDR1IrXLnC8WOelCd0OAgSxksEOP6GvvIbR2Dfogo0QTTYVYZOhfGuEGznf2QBLBK/0twaUbd
8z/KNJCJYg3dguSMDjd5kAGdQUDfjvgA4ZAP9XQVu27P2NO51eP0S6H8Ar+uHcBeRfGdcrJ0cq94
WCUSGBxfFojxZnRMN7jq6+Mx6rXoEK0+jP3A3EOy1R3YB3TDCjBVK90Ij16aTJnXBg+2RDYCTl15
u/dyiVdXjD74cFDOWdp3RFT8JfwYD0PLI/KckkCjjgAZSP6QUbxKHLwVTfCx+AL3gCCmEpNpL1RD
mmlcLsL2r9lGRW0rSiNz2plSbJuoGB3fCREK77+AY/RsODy147NU9tZvNVGEltM38LUESu/GwBmZ
fgUk/ZcNNaF1QsPdESgAbU8bO6qga5Ed9a3ZNwxVHmfXZas3W68sRfuexezbafQRU7unzR2qpzxV
ZU8fdB0OJYgONYYIU05LZnVdd8KkjMI1QPXyRjlVm47DOlksLm83cOWS3tPs13iWdmxrxalPGEwz
nAI9NGygdomTeqRPlaOd1lFUR+3WYdMqaUbhFzze8X5ToqwF6z7ETUW0K6TRVrzftmI8VbEaWziT
7H1yafDp17z30E/eFe+fDg/ZR4Sd7zexq7J+tKMEbSHdFcyxISaEE/+GnsuEMOzTkMUNlYu2n51H
OlaJFGeoH07mTxSXnSZuSICfZr+3bwNJW5qlIYleCp3XHq5L/FYv4jyr06C7lcqo/yp6RdGHnNmu
dy2T+QR/b695r3p0ij8qjKwVB7PeV9VmpiyYJBuDvhPB/WUDaf+a4g/8fbVIMq+eQ58Mp5yrihBK
L9DF2RbVzzsjsZ15ZpjIy3KFyk4CR53vUgbXegwAj+FlvXz0Pg3PenuEQwYuFRyU3M8N3qEa7QXc
kTEKZWhI8s5v9Ss5WysQQ0DcSnFT2Wwz3kXeb3oysfzKrTu6667PSDq2+h8rBNzhDiiG99jTO2LF
VOtv+aQG/odNT62XjKVyVVsXcMZKCuw3+dQgtvFM8HCwq6XnloTa8HacRE+WknZDizdR6eSAL214
I2hBcFta8Ke5cqxnHqXgiqWn2jrHj9v38y/uGuRGHv0dHSES96yk2pW8indtKPiPeZ3uN5onfKkV
G1i9UYRhQmPakL3QB+TFVaVdflWsHwIh0lhHLzSa28QdzTqbR2dnYyW/LaxnU0l6HxravFYGNeeR
ZdQCLLbkadN6Wdag47P9GbtraASNFpSwpblko4csQ9ueLc/CgFwiAgpainbVfOjGCQ8mPvHtsG7+
+DW0D/LOO5UHayFiJ44VP3TPeVrA9glokS4+FleeBKtREVR+DE2xhsza2l61v9awT9igSPOsnEeZ
6zxJ+impv7sjFOp5TLP8oke7nyUS3kZFz6uDVc0IVv0tqavOWKJVk4ZgxSZ6vLWJbAYEg4RUB/Mm
2UyeFtMFvwITdv47xLkeQkQKTXtDuZrTV2gBhYUIEOLFsqkPdSnwIiWP2dSlkdBAEzceuXLdJTic
Cbq7fqjlr8xFYVLaeIwwwTW7ZBzkdUBbatfezz/PXY9/AY6feyUsTvDALY/ljjhu82nF63wNphNi
J2NE943lPAzbUkc4KVKof+QsMPSzO8/R7O5l6ET+4B3cvF6cCYa1y+0+ctMTtfE5mFmHyX/O2xCO
4dEdxhwqN/arAtLSI1WXRjeRRqebcxmCe5HL8IX7FhGQay2RbTn2meGh7HekogOGnTQnhKyUi62h
kCb0eDPpTAzYnDpvfiuZm/H+voSuJn6R82byBhTYFPDcUpxizisM4er8g150oxWHsUsFGfdMz2oD
C8JGTAz13Zv5D0mjlbhqjCcRyoOluthgpTXeofIajjy4pnN5V/HGdI5cXK4bYCtCgkqBfX44aaBr
PTOtxk+3xL5lhDhn683TXRDxAcGfBBQ2ubqubPwU5e3dQGeqDzMEIptAmqhZvVD24CIH6W3SIFzD
mGj8Caqdt9iCmPF1O5V/dQPCJgu0GquOre5QaZ9hwBucYLZ8B/JvkJbP832SRApFFHxCMSIq/h52
9TbFWmywxBPJte8TMi7+W6bqRWE2UBh+RWN+vI3tQ6mwDuaX/xsWCa+ChmjIfhwBOpEbd7WsGt3l
kloqglH+nyG8JTpScS+SL0C07m0was9EpSpKOgvF29/OHTL5eHsOz8ttJ59zEkrKMbPlOuaVFoX4
TuEgtBQzBmrYhDOqx85VL6Ir+XKo73uYK0/eQIhYqMe9dluCQLUuAc5zQhBrwlO7qqfxiP84WwtF
13moGQYNCE1LbYsTi5po1g//QKHb9SlS/+dRWBuB9mOQGmYRwq1NiQOPxoXETl1bc/GNw6bpD7bb
8E2UBtjiAHo6gXraJKqdSF4iUjODtolYbMlchPaEBGvKpoxzH7DYdpmtsYaW64ctT+sHGIgk6HD3
ZDMP4BPs99Dq3GehZZ7t4xZ/p0DVdAEpFhsiMLj5IHh789qnHtyeqRrw6GEaAtP93372yarURIS0
T+ebMtzLJP8Tq9vI/O0OQ0RbaK17LTszAYHaHdJUNVMHABjISVhCp+khD/QwCpZIDVF8gIihIkol
uAdHLFRFqfDAeD1ESnRr6DqsNue45W7AAcaSfrZgsay61pR3lhOZk45zOXOcOVrXDQayqUcKkqS6
OztkbjMLAAEAT7/p8fwjKxI283sSYltDqwhGquUvv4sBbbsmFPGnMJfxBmOU0cjXbo2lQKrc7bUX
/NBXVqmGyXbdbUwrXcR3asFN9eee/N4HG7HHaiNCslt49soXgKPfX9paZBCsCgZMYZfFQBNnv9wQ
/BFHXZeo9HNODiNHjybAWkEZivqnX8cIe8d10/9GL4vnheBw3aOoKl+icbimPcrSnRwSiwkhcpB0
uKmn+61k15P0MWCjLcZ/rs1viG6yRGhcQmKRqw6inEOpeopvlQUnE9Ii1kuortRqMrL+fZsH7r+n
1kZIVG8em9RJx7VYkiFPsZAf5T5i1LlfG/SPsQ7U0x71jaF20Wgm20CqT/AJ9CXa9Z4EoCAE6DMb
nvPHDiyjNas2Pvnf80/SKbfp2xzdIF7H1xZOwAfKvUR6y+dgB5L3AA1Q1JAPy4Gpi+faTAfpish/
rksnqsxl4IONTyHyyGdmdKPpMwPQjfVxzr8IzKstg/3KT9fqzDly6j1xru4khG+SBCRtu/odqyS5
5hS45aFekdNz4nrmzhrXYB4DBojOXsWGnQr+RMGiN9IQJLQzNxnxH9x8oVi44oBywOJAjMldBDn1
qLy+rVqNvpzd762tGS4+ibJn9YO9phLlyomV5fs9JHcuwegs61rC5F/Sxv98gZaNl8Ep8h91JNkf
fK6oMqn7z14DCTxztzONUfq1oVFoWSPc6m+sZjUa/gzH5xCUXkQrxyscaHNNIYnTRwGFf/8TXMCi
ODTs+hzHzpkElZ1Mros/P8uIRj7USWQcOWbcFEU0/rMqnCkeRRZmhEoOE1kSoEvUEJz6US9Ejp0J
GiGvrNuSZXZYgU7EmOapnqh21aXzoklkDFoYDlaRiI1xEYWlIRFfSydeEL68tGfTX+g2hq3CX1oQ
UqHuWCV71mdyVV/KTPjmDpJrL/cqN3P/UDsj6Apu2vbYDDgG6ZleTSvI5zsJAGnnPtjumIDkrCFH
/7LPOFXVp4ZSVVW+mkDhk7qgz/WgYLCQ6fG+Db4vYQnAYK64mBdhPhQ6HxDOJEJ0pe5MgTWxwY2s
HWQ+yOb5dcpc7l7BXJDEM09HVeM2S+KQPrLTVpV3Ikp3jGE0e8ziFln59sTTKLOH7ArbTUD4cFng
KWFNVWn/jB3TbwJnyuD0YV1zaTk28dBVQ8df6fnekkRtvLjHM1UDRDkg8k8fBCa67hnm9Kre/Iyk
FtXIdhw7pDL+tJ9fVtsh5hIOHOo3uAP3Rsxg/zHpLNRR4J+SKJ1YpfI2xq/iSzLew80Qfmy9Dhya
zeWdwAE0boTJIZaul69y1PRSBQdIx5NFUfY+V1lB18SZ0F5N9aMhkWYFVtO2+TJmzaHnZpgCfPOr
cKFSl3Bh6IxIzMOB5zS5zftw0q+RCJjPofwODUILesMSMl7nKZnamW9SbHmrly4TcIkP4KePHrES
9DgyWjlbWaquTLqgzxRwWmZXS6l8GImH3Bo54r3L7qUSnUCGdOsa25Jk+JG3jr+V8VzJcsfHOJ9P
YHI7SUI2QCeTpZyofWrEALww0b3fwvga88i8UDgJG2phz4I1XHsWwAdwuMhfSVSjLXDnQpLQpfsI
WmbzReviuFXmpXrDKbOsxE0ApIoM5niT7rVCdjPrs2VOWUcarMvlWdD/IJ10PbeC4X+oIpchJulE
wBYm6QFeNKJAxxjFbJRQwUXFH1RGAXBtTj+8dXaiDuFZfwyJ2GbSo4FLbdOoAFeHrkdRauNXRlSn
00YXncDS42jP3TXD9/PxtVNu/pi0gZB89S+zq1IIzZ/SY3sVFTPD4mTi9Od+HW+NPy/voJmmF69f
cK4O/LfbKRfvv+XIAuoz8NulFlW+GdWkhFKOi+C4XlOMNFOHwbghY+F0NjKdJM18irhq2IaP/Ngt
4UmdSJHp+peqhuErSipW72GGiy/kKIefAYDOS0yfY29kAu3mzMnRdQc8w4zUg1O5ObKM+8jSvRbh
Ffq1DddvwzMxlrx70jaaUD4BnLn4A0Sb4jVK9YJetkVkyCju8cwQ16vqLSL/9DKMSzOEfIwRjafw
2jnJBfk11TazUGmoULhuQtdbe3+QDxMZId1oavmUNElRocOZjHNfpQ31b+QBf17tnEW5mgOZf7yw
V/wc6VvHePJGlylG6j2cQWha2EFE3s9gMkr0mZprDCQ7D+DDqvFFGN6TfD6drhJuWdnuyeqe+W+h
rTwjUKgoc3qlJIRAOwqxSC+WG1c0fk2NYrtt5IKNrBbGYfofgM4UaZMvgaLKXp63e4YEJ5Ayiax/
fr/CMI1ImbiSNzSZLq5MjIQsS5u/MIUd7mbuyz6xWs7GusCIAQr9PhI/MMopKnw+RUCaHuPu14gg
gwLBQ/Q7VQK9TbbGs5Sa15TalibYKoGiqewC1wFVrE1pQ3CWLt4DpIUNfqBCkZU/6HTCorLRU5Ht
9b/Qzd52V33t8gRdIRJWBdk3SeAieZO2eqh4nydgWtf2/OWEMIwqcw8YvH12LO0yKa2dKmtNM8Xa
8fgdoMMk4ohXBCu632kI9RqqOeAUnCpDHGB9fSgRYCApxnJQJPY0Ulz/xTWnuX3r7+QTdVGq1rId
UV3GXNR/fLQ91/SO93yw+aHWkC66fgC2ROuV3TYXWPx4pneOZHD91edzU0Dzt+XSWK3ZdjMJxe5m
KzcLhcOO+HTpabJ2q9QdA+djp0mgNtM2xnGwxUjdQIUWbPzv2III6nW0sQUsT5eeZyjz+b9RDVce
VjtiOC3zoo5WTCA894DKMDj+n89nx1Bv/k0fWq2TXDnJcs+lo3eSYp2+gB1ZRCJKuUc7ODWD7hjq
aH2WkIqrs7b+qlFxBQYTFGrJOwTD2CVri+hwXhsdzdLeqXwF1p/HqMZLg4cxBPyth7JkUrU0OYyz
N+14iB96TSOdF59ScZ5rQKCgTSCm1ZflW7aA8R5dEA65GAPbWQU/5j/mgMRjuY8cIuXsLsllgr5W
QbZ3sRrjFjeywD9kaYGSFe58K7QtYgtBZ/9zLaEV1xniX6B2DlC/THnkVyTQ9LCYJSrCicK0rmau
sRp9jOk5Onw6cAr+vkD5smBmK1KtS4LriCwh1SWIhm7qazUMNQ6de49/b3KUEo+q63Hchuw6JUS3
GssxclHti+5hpi57Zkh7f7K22fNKjRjFDAHhdr8ZkMKFztgiPLFcDIXNujFbcWVWEHR8+n2JSgXH
y1N7h/Oc70Zsudv09hXaonuJrkp2w+9y7I+FKduoxt/7Gzdg0jgyDMPZVeogFi0ZtYUPQq1xBhMl
+RiJK9N/dDtN8rxiWZ5iriPQ/FGTUKLWu2fR3fz0gJNzTdfrWRGXG9VOc+lPpQC3GhipU1du50bR
9EhbpXlQ6Wa68sqvfOuOt4sNjr2kbc1dk0zgwIiL9+eciXX55/YmkbsLOjKaNjve1ppg5BuTk4JL
XrAr88ZXAzDrZos4rVgwURnv1sq5glBcz91bRO0lQEclIUK474+ZCBRPRz3ZYUGxAL8EXMk31vbo
s2P37R7qo+BHW3UyHooB+XMH8zF0FrKSxyR1lQlbzFXiwWzzN/4ZB/9fMUs/8U64uwZRrpzPD/9P
ZuOJIl/NiyAFQb/iRlHdr6zVm/q2ED4WL5h/5WgQ5DMqwKrQB/o7PSwyGd/y2ULgd+JxADell/yW
+XhLLYwuaTsK97rWcUKYl/kAPmNdUM1CZTbKbBwngoJqaKyISTTClMQeSAj9HrDiSJ/bXpkt6rZo
GCcaktR2JsEaBlAB83lcBkyIKh5WUVOyITXrBgGg41fIDm3OrHwVyMgDQ9EgomNFomsaSJHEnLK7
YZ3IbfVQitR9oMuvesPeDzhx/F8Wb+QDKtGwVVa9dPpH48UuNKiYdgQxjVodfKuaSgPRlKl7cTyf
8PUXvZpufBw5F2Vq8GrpFwIKHWd/o49Vt0um5Qal/UaIVhAg78Uc2x0Ii9inL26LcRHVszjK0t6U
ZLb+3/z9HzlNRBg0El2XRwKAtulHIV1SiT+D5sIgC9XnQBFgQDgOe6VqQmXrrvFC4YOjsOeXZPJO
2e6lkWVgiZy5TVL5iOMKgVViWLS99F7HSPGryZZuxb3wwedmefGBI8vKA+1EcDbK/DXMplEBGrQl
SHvVki7JJwSw+jNeDcIt7UNBAGU+XWH3ZfjqS5JzxMu0AipXibXJPDjYLEZzd6Y4s29GBDJbBpgR
uFq/ySxew4dZSHPSbHW5250TZaP0sABoqSLD6O2l6z5MzqlwxBpIHmaAyZj6ax6oKA+M1nxyTfVd
V0uqH2Ufe/qONVEddlSp42Wwcd8Ll81YKJpJG67lnXn8qot2uqmRHW07faCzZZ+iO2PiDSf+7HNU
cJFH8P0PEnid/IknuzycD5+9x3/K4xE/UT/chbfVrg4oKPeCLbUMxMaYudfOtA5qJwJJw1yq2kEy
Ex655CGpYiZWDqMfo5zHGCsLxndhsKlvYyqGN5f2E3e9q5S2GyovdFGeJXldctFafaBE2F+1/m+7
Ko3aWAdwGnrf0FTHCrJ9wTlHkQBYaxMFwFCoZaT7OXK9B4UOjcsbTfvPjZzyqFGRlgVn94M4Jm6b
HJL19aHidS2aY/N64k3uFqzfsloPwqUlPa9GgOEpIWvj7UxXIsH9FimMIkypoFXJsBic59E47wlC
u3bpochkn6d5mlYCJGQENBmOn4UY4at7ekvirdqn4GKQPWDl6XRUkozahFm9TwU+hE7yuxede1+/
zQEvE6fL1W6TXW+czKFqHS0XvN3CyZFjBTT8xlB/L/altKPW1I7dGa4QRaYkel6r0xYOgAMylah1
qFegScxUfSd9tQVRhyQOhflF9Ivhb9gMj17NJYlTFTHW1g9sZuT3OjtiBMu65/o2OKCH9uJFv6pL
1WfzZwiZaZ1mkOaWo9qzE6TVWlIMzKAWAyGWlJuKHM0qrtUSdT4E6PJcve32E3uPieJ4Sq+tFnM/
PprVy0ce96PWbFlMgPUMJUmYOPWjh2+RdmwSB6NtqTPPACjwpHe1c7+uCvexVjlVCscqoStiT2+D
5IFmqpOzGMzSh/UU4tnffyKBRdUReAHL5C8cn4BnCaU6DR+Ns2O/siGFxhfcYkKY+XDCj7Lr4xgm
pLxsVqQo0W6bbHWlupeofwsVhC6ShpPR8xAHV/jltEfYADfdP+kMbw4LFxohoAuNwRIQnY7lnG+7
Co+yu2iT+Hc5n8bpoCyZeuf0ADSmlZdiWZUhwxgAwPT+FWpLXaCdVWP/xiRgC8YVtgFo3TH9T9/g
a29j35zbL6LBedXsH1wRg5/k4OsBhxPrOlgG2Dr2PTJ3e5kUw9SPf+6RO4S8ZPRH/wlHT9a0x91U
R2vaaaVuhieSDlJAaFyxA6sojny49woe7OgJ+o/y3g2sE/LoHicWBiiPeRofsv9UHSYEX4J2oZLh
77T11hIi4EgwyBMFGvzkyXUWO7boRyZXU7YLjPqWk1+iSXe6jo3vld5HHKqv/WKYQOaD2/cB1v5k
o5kMNKF0UJ08ydDFNsJJmDx2PvaNEkrPd214PiY7pZeo0G9ELM6bxyXwRSQfCBp9poiqTfEF1WTe
R4KWK5cF3SKNCtLcnpmK/HWZUr2FoKaKBugd+OItWyOJ6SQRmbpkKx78gbVRTLp15oYDFSzuIwql
iaQrR24MJWSIJcnZ942mRBczzGNWcr0Y2uSd4+QHWOCyIZNUKGdkMnGM7aeB+jalRtC147j2DNjV
hZ2V/MI8LdeoZR28ULYpvTp9qbKgo7NOowfS78QotUH4uNhNw8zTvPw17qdsWrClx29j/TzLtjkn
5apJj7eH6vxV3YLozqRfB6rlolJQ5fmMItVmsByj+xWa0b0XT9QQb6qENvNW1WZ9kl/R0A2xeZaK
teA5JQb2+a/6D02/PCBGqYlNjPDmK3hWsmJlQyItiKjXbW7glkfNZj5sa+oQZ4ICfhqdjzGwWtl1
alw70R8AoniiMXF6GkVigHd6rdabftN0r9NClkdebgDD0WKIC69OadQHmevWEOuaCQ2GFE2H+LR8
GYX2LH9Tc5TjA5aRjSQOZJqX3QZcUDsZ8T8MzojByNEa5xM/fmMEADDFhHN0lgB5edUkqqozN8Bc
Xw5QV71NYf+eGLKhujTAkrQB8AmS/a7nlX88KMo0ALDIDkVo8dm8Q/uTao+5kFXY4tJZ0NQNa9p1
qe5wUBet598crVgeG64uGtfgcuY17uOqD+WfEKbzhrxtnuodL7kZpKwo4iaGMzu5sxOeZPysMYgA
/giY0JOi0/PhaJQK55QsnDNZGt4U8f1N2XyGlat8wCtuQ/s9lzqqVX4NPA9fKMlzc6vMLc1c/zMi
t85VtLeE6JIZwEK3njLbdplSOB2O1Mg5X8bFfBxKkca/WTlv1gffFWBix0LGQS6wbnF15Oo5NgjP
bbDdFUtIpkCXMWMYWMe1goFMcT4ySu7vYMAOtab6WugrSPYDhyNzneGS8y+9oNl2ZnW5l7pkIyC1
dMp9S90czA7XZX0kq/G7gyN0AC6LqMmvCdeXiTzfNKqmPSiBSWZS17T2HqGixo0xz9c9YX84JYyy
7FqaKMiep1pkQUNzBlygaOB0LAtPvBj2WxnssFrwZgW34tgo49oS0qA5XqiSxDyaPpN+4joTxOML
w+Ib56ymvBO8Xj5R6k68l/mACiMULkYPlSifxLahe5G8oTfggxz4LelmjvYZqLsrxUQ/Ti4jP8LO
qGGO2ss/OeQoQYIoFQ2Jy7LP7NhZZC8r7lTdg5A1lkYXzrpxCVk6lQslMva7vDdvYa7gq+Ui6vsR
POGdD2PsvWCP3qc4IUIRgfcm2KsTWW/RMR1khpmffg8mdhlhLZOAIPv/YjEpra6ElQRKNNtbeqf7
bacMdcuOLer1LD0mKuMBjIN+u1TzGGg2sPWw2zLtOg9X9MWS1nG3ITlj/wYT56JTvlOwNXKvW6eM
MvsRDvNnuTW/in3kOrdnF+MKREWElh7E2FISRn8H6kY55cyB1Vq7YUB4xyyiqeQQ2ZZMMe/WccGA
tcQgEm0L8XGwm9kCJ8BRZ5FbnkdOJLx0dw1x9OXWKJBLakOeHjVHmqm26b2xqVjZ9fA9KBfIQzUq
nWUrm9uXnU4EKPIjY+4UaZyFZXtXdoR/sR7bSFSbz9WVM9o4Y3hUzFJRbc+lK50ZFmNBQmlqee8U
mHA7hXHD+1Lsod673d6y4ND8gooANcoMLbvjRrLNJGjuHlPD58BUs7ToXBjyRc8lbSSFrrFuauKu
zA7BWIpEku0hbhBQjftmsxeUz13KP62ExUEnbAmUIc0jJx2Qkmd3yeGzAeHjrns7FPGuvGiw3iWx
9t3jqagB70SOywr6wc1FyXPsX0tPzCYzQ6/dV4KJi1fTgpnTtWLaisZxjB3ieXfGnTkgD/KHxa1w
WzQoEqrzWin842Wq1pEVA/glQSsSUEiX5/vfRHitjTJII0MNCy5iQGamB9QUBi2cYjb1f5eCpB+a
BObCuUPfxIqD/eh2K9G+q3wdAcZFR4mv3nm0Y253C9NY9OOU07ZaWSD7jc+cIX91W0ph05g/Ya9g
Uv58FGUei2GIJFJD4GsZQdCta+xjitBQawj/44uORK6r0rxWiclqRzq+62VXVRGFid/CmpFitgIg
73V/qiF03P6TtbDoXX7ulrTXho24MzezGrlXPuQkYBC9nHwClaM3nSSUxaiEHN1ogQvpgAMNDEv4
sJcDPo9y4L2yvukgNIPs2G40Ks0zogfVzB3CEUBRNFKsqVtcrRHYI4vVUED0o/gKQ1AuYjEoKKIg
6AMHdIJafcVrn2JlgVssgk4Z9ib+xHVvKO+S5a3VvjEzh2Bv3lQ0RDSIXzqhEF34xRlnJiqTEOH5
bVw1cnZOP/+VDVZkImkyxqnXkL7IByK2YPrwCR0PnzQejT3hJmlopNZgh/pN9QpT8OlJVAcRCiBQ
aVIsZNkN38mDl5njYxvxcqe2B330OBkxnYuAUcuHA5Dr8fsXCfekG0SsqPr0pLnU8grTGkWhNtA6
VqhEtTskwkr0g1eudX9jQMusLqIUcZmdccZzjqGgwNdSsMJX3IYg+shob+iTCVy+rKX8svl0WMfi
7h9M9CICQOsgnAYdKgCFU0VdbES7X3nF1qOdvrnAY0rHZ0HSQt07yF8duCI4K3/ChLObpWKGFmju
BGrBYUpDZomCLoLZiDO8Whix06qfSCJJNb8x6ecAJLv1EiBQwrKYYC4xKBV6lF5ngfiW2/76i/6B
phDHGm7BH/FUdeOS5C7TH7+HQ/SdroS2jJ24CkRciIEKCodi82k/HIRePhlkEJxWoX1Z/ek0xR3W
fvldNvTQ/FyUBqLmUQVoio9K6zRKF+YKqpbHkYf4dDoqmYx4i4SqlEOciVZN7USXhHEF/h1+gFyT
P1bAJMzLccgHBsqr1Moh3NRzqgWfDu+sdxizGlYQNKbrpaZuJRp8/009HbCVlqWqcjNZjrT88+5R
L8rQSIn0+UBgFQ6y7SkbyPQBwptF2Phml0ho63T/xWcDGdisALiIq16p453ncGikRmGkW8eCA6cY
RxtUXh1xjx06uLOMYFMaTfMe0OfrSTubjvmcHyG1JSqL7vVGkisq9IbqXvAuomPCJl/3cIcoH+BI
WBgg/zBOYaOcKGLUVNnf/sJa2kv1zI09JAwN7vbAALdPsnw4pNDw9kgJvu5c1br8srUsnUtywo/Z
dPARNtZOKfV/6XWCyXdIvwjR2nfs0fjhd2/BMQ1qqENSa0sQA5iFU6FSnkmNfveQZc+mQVDmI7PK
u0qsjTjgPzcb40W6Zih5sc2aMu/2O/yA6yaFqQS9HCUE1gqv90Dvbx2OY3ksEoYq5S7tUFQflkqf
JkiHlJJwh3ywG7twNKsY9hcvRvzELk5ZQEzUgK+dOeptUfE1z8/9Angsd+dv+XYkBaB9vxh7Zrxi
IM/sLFzJ7UO6+s+Gjtg0CBcQ6bqLp16vWwyxGuWgeaDhIsUrrLJqw3J75qNRQ19kYgWQWXW9f69l
I7hbOfFxtFUz8jFicBgM4v8iErgwdlBsHBpxjdAJCcZ/4QhSWBD52jzy72J23cOQd14msW/jkGTG
mTLfe1ZIhucngUta82P5Y+IKzPqmXYBdxDEC9+EAOtwhfAdZw4IlKP2TwL7HbjMBv9S7C/Oy7ikA
oIFtmyBvNV6h396kWDPIE7jAy07B+SGWC0M/nuxHKXb8xvLbE710WN6iEoleRKDXRG/kTQ24R3tO
JUawP2ciQUx4zMGB9QSgWxw7OEKYd2fMdT2FQ5GwwD6QRXba8yBgr4k0Vo/N/YFJqTeYtC/yFdXc
KQT7TxZi7BOsud9za9CpTJ6KVQIldEt1ukQbHZknV3+qZIWL6j3vMx1lGJ9X62SWlR0nR/eNEHKD
Dx/ymuHE52oZwnSkMOfbnA/z5fxyCqjbkN8kiyPg525xlE4rwbD/aNbRDYAIPGYimEvU4NtFDIVp
IVpQ+PuZBdv+9WFLluC0UVYZpVmVthAGqayPLMA1uwjTUeH8D3bN49wofhXycE9Js9jSMY6P+YkS
055H7+xbGMl9j99cURfe4qAFcyJAZkZHzGNK+hP4qe30Z/qXddzlDc3oX12fkeLLnhBAqNlQxSwo
HGZjPM4PYPe5CJor3GY/sdgTwXcygkWA/+9gC/0thBOjLLLP0Vpd7R0cr19lVkjHW9BxlmPOa9s1
RAIlYOdTxgVWvc2eL84KuzzMKylTWk+fW+gWHulvbVuI+Ogy7vrX1nePPdl4baOPH02qTk+miATc
s6Jf2nUkfHDwS1WuMfS8iCoJFLUS+3pbY6x+UeHXKzF57RaBB8u0sQNZDSWf8ymfgrtVfGUcZGbg
0wx54FA2xb3grK9DSDbz0eW9TDkXMt9k1m6PpExA9NOj5zxhO4IBmaEMcH3J3bBoTrG3R69QQ4Ek
G+GA6ss4Y9g0AqXDGNNsJhZGoDCdMfWrNxxiF8Kydfg4rVhZ9+dXs/wdD3sXQcWTuM204x1Ix3tO
T9erVrgUncLLtqxEuwLSD6tXrRdim2H+8FB2uS5L27FzL6OATLGxewLwDSQOmueVT/WFOXUA0OPF
pMTMCuTuhywvD0ZVJt2vdQop8oV3112pEOuuJUMJWprCZ+T/s70Dl31jyGg8oE/f354syds6Trk8
pyDP2/2nvkK+kTTngPrDfyCDSkm5r2v3eRSkZJRySJorP2y6AsQ5vaqi3u82MKjaw2MjtRzuc0kj
jRd83uw4bLCkJFZWbLLUjwBPI6S50UH2c01QxKpewaBxngcGQFGIkmJOidm6PR29ToWj5LglWU9p
Empf0yYDa6JXrSLndbej4cUFYc+ATLNoJ6ddcHymrnZNr1jfxoC34+q6W05oAkydpS7fic+YQ7qD
KmYwMYS2mqL6d9hFcRckXnHl56QPgz3rqcgup+lsoBo3MrH88NbtycKUmEjRMoyTcCes1UQRN2bm
PZoc1x+ZBKUr0NQLuR78qyNDqa1BDcfHUszMhDhixqGsOhbaZZi7sSoamgyZ5osU0WFvbmhD4PAB
NXHGWWsvH6ZxMgTG3sLJ3TbiRv6WDQ/qlWv0Vr9hycEv6L88KMhWx4YFFgj5BPaGJKzVTn7Yd2Qa
kuT47k4NfuEGPETk/yUu1igMcf8i4xCTAdQW48nTOyHmkCe+y+PDJ55T1anH6UWYOQImVDTYjLAA
I237ph9KzZF8Ql9aFEZb38cyLTmC81Y6NbUnqb3ToErmRS00EpTOK58P6wOGNUMcw7iRQV2Z/Z87
aXQ0ACg77JfqSrq9vtHwLTmSvjWU+qozrb6E68WpapFaN089QaFAuhT8PbTJV40UVX8Ow9KD4qQa
bCxKH38MYZQOF5iL/ACg4TRTHETEV+2XCtNhJ3oaIhUpg092N16apKdb//h0SUxvw9ZQ+CF8q61j
6/ApTSMgNAZ5bS1ZHcIvr9xdf3R/Y6LptCKjBdfoeMZ5Frn2b+/105M1XJ4F/GUzwLCkQ5ka5Wsx
qBgdGNA0KmR1UHtO79ROlyJEI5m5E3UWPR0ZomOErBJ5vb/u+Z79a1dMRx9h1I8quDRCCNAvJiue
+uezau9fHLkCKbh8e67YTjLQJevshEbSL57iARls7wu3ymmN5hxyqzj5uvlxHUUpzESFK5KUSR82
q1Rtk7t9R/NYlPuiwfyceSej/jyVGSmp/xciz+VrBQRUFf32tZi/ks504xmlde2bp8LT0Ms0dwV4
ZgBWpRq8APpML11cW6u+I1GF4kpuP+SS0VgjqvUZpRO8hgHtH2jmkRoRw/N3MhCtflZPtp1wIqut
rFRHsgE5ERGrNe4i+AhBOygpexde4nM0QCgKha0M4l1HP2mEhMNzhKfQgE1P4cO2gVLqg/xCzIZR
YzNcPO8e1E9vwLBPbXK4Rysht1fkCJHK3aLR/RpOw9npTNr0tziAqmdXA/Wx77YS+361MSIGHMkY
AJAyg9/8NSOZNTcn7OESkDErA1RThcAJmbzc9O7GxIiB4q/6SBidEvOIp4VMCcxSJOPnLTAR211J
bX5u7R8Fzibp6yTJHYSNRKc2i/x6e7Qhu8OyE6z4o9KCe5RA+xrnQHi6xHPXWdVJXloQZicMGoAH
NIAURWA5iaSRtEhT/gJfjHqIIpK/zk9MmPCP/I/8Kcf9LH/vLuR2CE+/QWc/EBT+yod6SE+ntw30
o5AqtQpTE1Nu4LJW7zYaqwFTI0J8kEuRuN1jJ+eEVlq2uZDelLYBFd6bxv+76VlesFR1HWWoeVqT
euxF8VM3VlLw7ftZ+vI9aKtCMSKMQ3NwkxBthBH2CFqJgjnaecUqpALsozgjq60C2/nJ3iSyKv7/
KyIaSDKUJbcd7sguon2afGL0I3SoG+AO0XM8f60/ixOkfy8h9tOxOGEFsc4lqN/dhufHevUV2bXL
cxdfTGwzcJre8jahgfSo+UJ0l1SUC3VX8bz93ZaAzfslO65GB/BRhShhC0lhX9vvRobmQUwjV7tp
EKd7Rm49psTHKsRUGTlNLpylI57hp15q8NaV0dMpaqnYpltGKltgYMl/kIVERUU/dOFC0KGr5p5u
ASOLiL9BUNMQXYjnl4ucLQ7sC4BJU3Wo2QiaCtJ1iwabBtWj07lfTG82vKz1FW2ZPq7GB59HoQn5
iyso+iW+qb6glERjCPe+YQFjvMbz77/3DDyHDNKxzoljGIJp/IiW/wJjvwwzAIzFjs6uu8HMzJsw
jCRzn9crDvj53CWy1pGPAih4pZdzlM5KimI95M8kjxb3SKmefZfkJaAKqT9lqPDgJEhsnxQJYDY5
DuqxsAfwzcrvcdnjmeulemzARfsaq/iCQfVhWEXvQNDzXxoakHRdw/b/Attfj8srYbwvClZWZoG8
W/Rj6cDmbndo+TCOcdojxaVTIqDlFYvUynSjOl3FN8+4xkyrPS1AYJ3Mx9xD4FPtNkhi0DNB9ivX
EPhRnBHO9cVR9W+z66Bf07e1ulBEXnisLsRROq+ONd8bzjFS9wukvzyoXVPf7cVtYRQJRMc3vRZK
UPfKvNEtFuIubC26ZMmlckwbHGqwMGJp2Z3TmyfS+D22tSmCrgu9Gug54bPsurRKnG26fWtn9Elk
1yqHqLSMOzNhk/Nl5CSyxG93xM07jq7Me4MDZhya680RaHiq4amkEXXSWvYxbGhZga6Zg8aGwh45
rpm5tjO8Raa0b59I+7WMRCSmXUBt64PVQ8uTtA7lvpTAumwbUQBvQ950e14QHNksT2VjgJs5pZ4u
bAQ463ql+VI9fHM0tfMGwHvNnQW4zrFhAkgBrB6s665o8yfEii5gms6TY1TXUiMhWmnfkES7I6TK
yrrlhx2s1otQqTXBeIO0qVrmEIdO7Re0cSJjsoVJTbSgAidfCBLWpSzoOrqPogDcZxxNEzzPPdRv
9df6jx9MsczrmdACwySoSXRp3ICJUymHXZIC6v8IEydgq3tfaAJiGSntbmJaKy01UJX/UiPVUoLs
Zs85ULG/VRwDICTERqjwAGdIbgFmduCKx0JgXB8ahOUd1iLQ2nfLKD6tzFVfDK/N6qDC+W5eagP9
nudWeuH7Cjz43lKKfcabMTy2vQKuK0jeyOEScU/w8Z+QiakFW3O0Wi6U+5SxYV9Ww4CzKsu1OmUP
p8fgJIkTpIAHtiP6jsl+5lvia9YCWE3Sv8/5ZdRJKC0tknLTc84FSauAiXEwz/kvEFwCNJgOquhA
Tu7gFY/WUMgtB5Yhd87O/FRlC9m7za63ruPjImeHYlu1vnUyX+nwtEMpl/hw6VfC+Pph/mTzlgra
4vMos1qiDIn6fTSvWmUK94QS16C3UaG5w+Aq5RNHRzr2Mu1k9Rghcv7Il/BOXcpQpWVU1H7TIM6H
c1iYSfsXsXBLBaR1N+KIMkgPsB3IlghssCT3o1VtNkvSeL8Ms4dPrg6TNZWBmh8oR7z0KpjhLHbj
9iYmeDh8tlr+JhoqecTzwp8xxeV+M7Bnc6MhLTI/r17S+ZtJCBSDJM9T9H63TdCgVPVk4WzA2KA+
8uIw8T4OS3bHvA56rHpwe4blAoaiPzDL5oH/Kr1jR0JFQR2wb0tM7SvR3BvqYzyie1tl1t20aOUJ
OAXYiSuuZm8QLZQw6YQtRnPVozXa2TMFjPx3GGFY+UCddkpeITZhKTXbamgvtq/sK/mtXvaYl1T2
4X0g5Nb8i1HeL6kEnx6VJ/atvCCq/Pw7Ok8PjBSrijezJQm8gwQZHBiYUcZ4X7Lbs71PvvQbIPXp
pMwJVdS/W7h7DA9N/HduzRW01Kshe2eMjq4MYhyNCcOwdn11jnRU/GcJzXzYf+3KRJaFyHJ/aCAT
+7b4dxQScFgyxUXoo4h2IbcmpzwKgjXlLRTeLwBljPJfaVaBP7xiaOnJRDfdde/14A05fuaRYTxm
cSXAt0i8zfB7i+00QBAlbIeMgnxQ2mFBomRZA77Rl/789tEzt2uZOlDsk4DXB5e9mXQoUUGG0F8r
ouLqHR/L5lyxDcwR7eERkJDa1SCm5E+1BswrdaOmMlj93M/CPMvyhnJtiIPpSks4TcpyQSjwIt5u
pBf+pxqf0Du2AocAMTe1E5rSYSfPmgqz/UefKvUjg2F08ySXTL7SVHa21xrVjD4ZtTVkJJIg2rD5
WoxIg7J1rYV4Frby75RtrrncXfQt3qplPohbnzY53Ncl6nOhgRM9tbbCH+hKbEFMNB0LRVEblMHE
Ad8y1ICEk6jftBE3OhyhBe0/BiD8+Xoxy0+RcaS4hqrPp2fo3TnqED0k5ttcwirv3nGeehvmMHq4
bzwHjR+Astf1JfSUrdtWjz/45xjafhRw/Wqgpn+uoBA6Fb7uSSHHdk2856z/ePid5k0atvPNEcpi
HOt24RM6mnuFxl+yoPeuGvvFp1yLfDNWV5A0VqHUqr0Ms1gAM81WlKal36bzCASmMX9Eklzmd+1p
E4pQ4SWk2/PuVUJ7KgrBJBNQXPh1cyHr8JsFUJDuY6506j64xmHmoW3q+NuE9RzZe/v73WiaupYQ
lp6+pFZSFmJzWmMc2RcX2T7EUhzJzGlG2TGzqpdeeNS6aVThtAIEP4el8IXntIO26YKK+YJERMpT
VMdeXhEJplw1fvm6utwlFfJVTe7JCyW/SE1WqNyU9SFHn4dR/GCS3OTgs0ww2M++qjFN+p8Y/iRR
JxpNmZxv5CNQTvLA/f3TnusS4EGJ6MXFQ5vSuhYhNGD3/q5nLa7zRLKNKubhmVbssBZdRLhnRzTQ
Ne8LXzcLvWzF60ASRVlr2clk+dpALAfxvJJdTczrjyiOpk4qGWdOIyid0La+1jMEaOKmhxYzyrHe
ZXlmyE/lyOVR0EpFHijDxla6K3FUGezfioAyYfsMx46CIAYQp4r95Yuii5bcnuKfPJyPpTyTtV+t
iKoA5vieS8Ouh3V9Pdt0ZWicCfyVke5yIW06thFI7zXhSeQB3mvQlkgOnRs1aQgVxBr586k5KOj3
c/7MW/rle2AoI6X1gAnysyx0LmDZ4l3FtipPLXmsOZN9KjNJHIAmJwIEgGGdBLJAu+6gaErF5Q0L
jrq1iRTZmQPG1ZG3L3VwVNPohB7rmjOHpTp07Itml5UgyAJU4E+SzrTIzCChbRGG47S96IDtJi6v
DiMrIFfJkvVcmB/Paw5ir7iOJFClg9HeLDopm/rwcEP/uZYkLKORR6tPFAur5H7jkgq5PnnQXKi4
YT0rcjmy7V/6PQV1rTDHMM6AlYWK6ao4ZNqWsEhNgk3hxk2i3XPNH1/REnOzYFfXWhs84qZuINyi
Uf3fvAPnx8+9NAfxS7atz6OR2Ii7myHmgzCL5VwpQm3yXPv8nXSqvL6lion+l02pDr2WLBQYmCOu
la9iWnq/XX+aVO/fpgT1I/WR9zPjiTaK5ChlybP8WeAGjG/pQjb2rlDilH0B8vfe8A40WvLcb5Ji
MDp5EaPoh0/ay6EL3bwdbd+YoI7X54E3xwkNcEywICj6eKeGp1j5Lj3SQKCtH15GkiEJTYEjt8ru
+hb5A3nFOHwsY2IVz2TkmorNm6mKkoBt8f+5v0PxK1BwbskT5Wtd3zsZU3UNckIms3kzGVzK2UcF
fRm4s0/Id/nrikl9lGs854HKWQr+LpMGJ99vb7OzDtWhPQcCT/ZErPth4tOnY3DzZKVQOyb/WLlG
pmN+2RQMPo2w4Pxov6iQgYIQUSupv+MyOpBBVmtYifJqY9LjTSm4bcKVwRWwgFxX6AxeD1iJIwKU
Gel1I2fQS7JQ0bb/NAn2pWdwAa79tsJ/avCGg8gCpXRqmzvQTy2szoHh7gnm2kdxxTUd1CZMXD0X
7aU5IJOMXm7zhBpK033fhpqEeYyMYwLksQv78UdI6oH4UtgKXqlVJJL2iClvypqNmeJqP+LJ8Zu9
+n5O+Mc3zskumqb6ovVODgsxN//EB/22YbzRqy9FgG7Rb0OvWObdBIl1b8vSMv/gCsR7FbJiRBeO
IDSpenG7gou8My6yHZEMdOUpBt0mOUSqJW3jJ9GY0XMUtPnkgoqKC84o3gcQGQM1UJ1BNPJ4QKlc
iov3EKJeS4VliXy2bVzpWGWvbwUDOTweR4UfA6zrfKHn0LBamj78GVCTwnZrHCbOyB1f5YaC/eGJ
kst7e+JL34G3s8pBipy2vu0Q9Hn5N1Fu6IcMnfuW0RDSQ/Ovy2XHm1I5PX9abPxNTjig+V4Elpis
dLZcJBGxdwnyGELeYDPEU/peA703KOVQYEDNWFRb9AOHTCRtyi3JjRaMbpQwBJ+0cRiBBWLF1RzS
LGPkHHB5/78DY/N/Rna5b5P42OQsmDaF1P9fcIUhxx5ZnH39E1O47pbVdpwjTrLCw7pVV7jZpbvG
/vEE99xqjSV/vsHAIq7By/ub9xlBAg2EDmzoEES/yOHBWUR+J7+AF2PjLcD2WHZIpKb1S57lsVmc
dQdnyjdAxZAfvEcLUwr2NpU+ybHdI3DSpUeC46Xyr+IlSzOOI5Q/YDLZeeRl2x5KrgxSlTzB9FKH
RP1OZv7nO1nx4E2xEBgRrrz/1Bss9LXRZUORyxtcpb18xny8Lh5ijmoVIKMbWJ0EI6e7PVtQpPMc
k22VsOq3DWIQfgjtzsecJ/yCG5tXfbE5RiAzjkGGyA8H+IP1QMN55x6c+05eT9VKcVdxR9dr/MxG
7YDTgS18shjDfvcjPEcFlr1yZ54uND3ZYk3L0y7mUoE2MLoH7xwo6Sv8zc/Yu9wsUIG6cSQ3WJtG
vkz1ZdjrVKmBYQoDk8pmWsCksGg/A8NJsdf+TpkaGxuuSHTF2jf50tFcjyF1r+3OM4bhoKwVLybV
mA/7LetyeZ0Rzn78Cvfb3iBUpZRN6AcDPD/Fmt1YUBl9XkML0MFCGr6QiJwLT4Z3Tvz/b+LoRHo4
hRoOoPpLMCQv+kQ4pIwCQC3491AM01QfPhDMuoNeiEz2/Nf1/zIXe/XMOokrTaVcFzE6LR0xwrdv
j2zHqh2P0V7pILg3JKodsxHgJCTVhNcCXdfOIH1iVSu+o2PWaA5S64aLFZbwnexTkqiGxj14wCpZ
kisqReC71Xx/wan2w23XIpuENPfeJJqV47w8Kgb7Jk+pZj8Gjn7a9Ajs44+pSqcSyfRRP3hGXsgt
qx7vecfmCrPhxELiAj2b9+JZ88yjyeIs8kBRWM0i4SO5VeYmeJ1ehI8YNp7ezD1KNM3uQAFmBdMq
tnXvG49dHlWkMoKzjXsa1dVXcrAjK8VG0wYSM91K9hkWiikq9FpqQ9Fjm6GedSSwI3CalyaH0iRe
6VuU5bX91x42v/Xf0zOjiswI47e0ldZQyweQGjyfO8QbPw4ZoQZNL90j/e1+xHQx5ctTxx/JZlyP
YP02M2FMmgUgq3aiqLtXRCsPa5hdMqXKKQPw+88NmRyMjb16yCAxWr3sEXI70sBFNfV7klDep93g
+y/P4zaQW8YLAiQgzLLwvLx7KjV+F7DIhwzup62kyj1kj9wlgQvfH7i0t9krySG0jDAq7lCIDe+2
aSN2+syUwq7eq9BovADEWFkYAwFDwXqLHTv4Zf5nX6Hzwp5Pr/Hg9CUJqTIF5ygzHboOh4byuATW
i8zdfYMf0TTb4FI/BIZ7p6E0bNzX1LEBKg/xvVt3fv3RzznwLCLUx7XJ48KLrvTHKS9LsSuIKk0c
uQUkUeVkvFrOHNnAe5pqsqEkhr2GSVC1XTuZ1uNyqAPoqHqKQld4Ch3p1x0qjdlBwxbSL7rPkZX8
uEWrElUPQzNdCIR4KWrTWFxNzd70SEtHo9lUjxZYr9cWJLzefV4RqEvMY22Zm0lIdrncPgtniyha
frQKgfvo73SOS10zCRgc6aoLIbCGLliAfLpGY/K4U4SYKoJSHXbB5wFTQDeRq29fDueMZlI6I7La
6sxSg0eleM8BnaZGm+NQs274+tvMGCy2JKqEMLWvO6qnztCXYcOKhNCrY2R9qzD3Git+gLkx9xaL
xCI6RrrTTvB3q8sEeEmRpVuiVxrVXbcaRHxnDaNLLHtb8S7fagPE3L754GDh8Y/A7lLEJd+vaI3x
NUTg34C59LWa4E06CKeRzTadY50+NHsVGWXhgerzrlWKZAEAdULN7dIHl4OG0K+F7McjR8H8e0sj
FzdwPxsW8XsClKBxr8SfxNOi6AbSXIBzvMWQzpNaGJJHJjY3pDEpRdLyfCnpz/vzo9vFAQrydw3A
7GY93z+D9ui/PGkKjBnYbxcMvrCY5x8BjxbJX8wnRnMTPS1mgo0e+cecnMrd8odGgL6KkLKszsdX
4+fsFPCj4K8xsdoUqVMXkGFM9n4Bl6T47OLowt/K1eBBH+ubkhKtLj5wLFEo1Vb3bCju0GglsiE3
+b+iz751EdbUchfCIHBQTVZzhun5ZnH1WuBGa9VjQ9wIkSFvNMgM6hXQ3JaghlX7Zpnpu2el2ksL
WEp6+ryICi4Aun+qLU9yMAyIIZWzsVcmucQmwTflruJJa7aS4CHk89fKoOux3gILEzS1KuBIXxHr
4lXE1I6jT0AIHbGJJZLuJjggb6cgCej7w9HaDBSWgj6AxdsDwkiACI54aBU5ynz7U9Br/S/XwojT
jmLwSiAPA+Ed8MXKrIfQHWfjz46yZ2SBcdnOnM8O3Zsffdo+CJY1ZiISXumxpcDx0ll93lHBTPST
fQz5WVIZucY4nPGsontscrND5pzLak68Bf4KNoAE/pDvG1Bg/yVJE5k0VQpUGU5aWceSARtXOUqk
NoylrM33MnxlEpAb/xcfCDxqUNibtzbUvvB2jcEkci+8ZmRU9w4xNaGhnITekTzEGHoiK1RFPlaX
Lmnr4EQ58FgG3xtX7wE208nlzTpVOXLx9buwIl0sW8ZWaDf0yjJIB/lFKSGrA0ekj9eWzHG0rz0V
dIwz3Dhx9B2H8n//GNy8O8Xbv0kDHZEbMe0wSivQytynS0UdImMsOVTzJX/YoZY6VYS+7qZsaF+y
zjXL0QI9ivj2hJA/Ki0BvVd1ft2/wk2RS0/ofwroDfHMVpbPO1pIzITKpCTBEhSheSbSjyR4EyJ4
n458uFZkfzx8l5xwByIdbm7mjzuNcd50a9XOY2mtvPDqhhd++sHR1Zwiml6Tz/EjX0BMn9MGgwOZ
S5ke4DhQlveaO/oPrh4M+QfG3MSlOtlyLQkBHetWp1o2o6ccPJF2CHeH6P09SelXQnWFSjRUFzEk
ZMwx7lRXNvVpxmStUam/IOI70QJM72kqaD9rr8uzugZGapztXblOLHnoDrUU1PyB9YTLRX1R0ldh
VMhNkRwVWwrjEGobT5zbPvfbjrov+Ljy6vd4e4UVBmZhdOtcv0QVXqD2DbRxP6ltW+GVqENk1TXe
14O3q6vykYZcV3u04eKY3FbWFrjTzCkENaU/YpyJWLWh9BwgoKPIHwsXj6Xk0c9PC2B4ngGq61kt
8G4SJD+FYwoLkhfBTySbcRNlYQ4YYAHC1lXF+W48uPHTsz+/lEAKAL5noOhZ+UuBZ9MOnpgYCpKT
oBN3w5apP7JOPjSXsO16TdRd1mcuu7q7fhV5qNrGLgaNGIWtMjSdN2cf+WfxoiFnoYKJY/MBpbP9
zrIlrYP9TYtl6D2pFTVIMHXtgTJ4toQrhdpetRqO6JKJjOkS4OI2N1EpCTaUZ3MMpCEkcZZqK2iV
V2LsXKSNmGikJWGRomOFdz0cBu04B2tAtBMnhiJzsVEz5JHGBLMMTo4QJiQX+KCiPzeKg/Fkusj8
BoV0yGq/fARk5ZhgVX0iDKGDtWaAtb04Kd9bUZLdluZBbsVgA4KP+5FM7KH9HkCnjX+DiG6yjMBW
2KcL8CEtiEU2emGFmiBk5KAw2LdNa33rddUKoZCor6C7faP6AWwSgl5DFq3YC9DFdIpojxHR5AW6
qd1DTRwgcSQlQ5vH61eQjnHlDvP6S+YliyBZD3n7hGypleAlOI8cR8IjIriOVUQAsna5BgGUx6BG
2AbDl0Ds2jAg5vI9f1d2a8l5aJV7mtmZ+2pxRCu4h+OhZptEG3T248R6SO58cO6utUh4CDDgnKOc
Fc6IUJxgjghya9qGdzyA095+lU0WnG2dq/mfQZDoiRcYpN6oNnd4ckC/gxg/aXbB/o6lO7Mx9gp8
eWr+KNCPOKI7BZ+k4jCVCPtZXy284W/WgaQgoSBjakVnUOAXh/uM3RUw0+SA50u5Fr2WCvSbCHSx
4H9/Qwa8BWkI26LVSGUtDheEsoVxEpBNe96NwqChZcX6nyyGLHYXTMzZZHjGma+hdNemaXOnJn3b
95LypmdjViJR7HfmJAX7KXejbfjp2c3N2vTsPu+B4BBnSk4j/WqPnLzAd7OjNagoLV0Q/krdh+36
O7JdgcTB2eDbWVjywSbCzFxrdRc7rDR96n6A8WdJVjsUNZZn7SBWnhhNCcOYV9DKdC2wyK3DabHq
yxc66CimZrsUoaHmxjSRDsagky0yC2pJhYAAg5b+o72tqmxtE+JfvxdqbVVt3q9OA6DLwQ9oRdOE
HRM28cEM2GBb2ynZHXPdE9sJ3v6X5lub/phQA8+r7Q2/9FpjdBksljpCGWmRqRYuQiEuxpwH6FHM
Ki1QM3aDFKcfaTkktQOWaep9wbXcxJ9nzTqZZij/OaiGEZcYtbvgDCHOTG4QOgsJQTxA9ps5ZHBN
JK07XuIVEdK5DXBgCJ1XCbQeb821NUeIG4blPO73De7mq6Hs267KD4Bs07rn30O7AfQsSlP+1cwH
j9FQih0vYMTssDhDL1+KeaVty/E4QnXM9LSYiRhKWDnbUlTje/1gAobJkvrZvBnLKrd7nMIg8xHF
IluaPVk3BtUthDurBMvIi7M6zcwXevOQsvo1GNfVNUM4PU7gsb5WeP0aNI5EdpXEAE0B8cSEGHyS
bYEs0q4Xy3vEE5y6mDjQMDpNgCCv1uba7QavXPZOIPn/JFZTTqCdRl1Nq4N1hl+dTZlsWqvnRlGl
nrgi+WnbF8t6rgL8vdtMQNnr3vHyeUTlcAfDjRpgzlFJQrGpyu2XdXwEL4o8fIABgxPWNVWMipfq
8I9PHb7GPm8cpfvW2JrOOcyIyZoijxb07Rhg/KJKgx4f5SYL/zVQlRDiHyh0t8icyz6dHgynvE2l
o6PPgOD8X1BJu+Fr2bTGsC4DJmFQhDJF0uCP6wf4ZkSdEYrP+En6Jh7F9jzIq1BfgOaGxcgCFeOr
HRwo2JLURCtJLbxW/0Msjcrdoewf6eRuOj482K+cJ1U++Nr9ulwwrj2Z9ZMLaXmnVMGyA00Jbr0n
zr3Hl82Sw9W9YNlkHTGQ26N04qQ/pE0dgqB+7L5cjyV5sNZTG2WPy6sYcIxk+M3/LihxPQD3KFiD
P/inMPjbPlsXP2/3K10PJQ56dOlxGAY3aT/NLYcc1EzYs187vglsSe0bQSyVwt6rTvj0Q9IiXCGv
TXfRfTUF9v4lOjFtGtfaoKD0vY36dvWLHz+XvINUlkbC4/zxt56avgjlNijguJqr4jO9mC3Zb3GX
j2mxdGyV8T/UaysASQPxOcPf5F0opVVBaHYsr8n0SSeIexjvK7Iy4CxREsHq56ngXWq8DgnDx72R
9aetbl9ZfvlHvkA6g0lJim1OY8fsWngidr6qUK2TBWVFDpC2d6aiBhxSqeT3QGLqJPSmw8wsF9sB
+DjEOyzzYy13h5axA7ihw9ateYELNhHFcQsRiqrmN7R35wm+XNNhMY6k+72U+vIJFW4SLnoCnDvF
wCTnyM+g73WIJMsz0dbRVPpZSwQR5e2Mm1CxlTkm87zfjYri0zVjHg/cheFQhGUidaky0rR1Aad7
908innMTnBt1RQKr0+q/mQzC+zgLcrlnGsN0fjMXAYkcVOG+yN4vrjIJpvq/rVLu/b8ruUzr/Dv/
cyTHMZ1kVQMz+kOfD+LfZMDQlOw/1Cm1mZwrs1EH9oDtvnU4S84Dd5Zp3evj3w2CL7mPBlCf203h
ziUKiXppL45nHM3RDQ4/gXyHy50Qfzhzf63ep7K8v8aDIOBIjcVxdjcwLRFEj90ehHIO+Mc/ZaUw
ls6lc9UO6PY4VNPRQdcDMK+QtmK7Bus09BT7R3Za4brbrLa4vHqQW2YLJHMpfgkO0brrz45zmSol
qJTZuU2XoXbADAe2vkBl0S8OoUcE+s8j1uZE17OLlqXfWG5TQRo298SYFIWJ4UIQ5RGp2UclM/IO
vah8rUza5iT8CGxlnmO4eAnpPdR8YdSzmn9U2J50o/d6v9nSLjDPXoT/74157EFN2co513s2Z7Sz
jAwKQoVf8WcubgpWUzTf+DWLsE523DE/TZz43ft/6dyEM/5tk69YdWxhL3x6l4q5TA0ynibO0F8S
5j+l4gxi79Bw5BTbTUTi76CQ5YQsjZjERmQUzhxeDzTK/XCb7m1Np7IQlcf7aItZFEhUaIhycocS
W+L7x8R9gtMYWJvrUrpli8RzYxJMAJVfPkWS9d5+c5w7W0nd8glkDOTpDNLIdsV0MDgE3sU5Pxu2
AgSx6UBqLYKatD+a6oPiZUXxt1lUkSWWbxunURpA1CXOI+YSt+oedO21zq16IcbPBiez5f8TV5RQ
sy9r8t/r5mPA4raC0IiAYHWVMPCiLuNvL7+pTIYpWj0IQYaxD18xdyX7ftI3a/02Rt+AVmbY2Kei
A8t2lOlI4q7pyZfOVgRfFljlCoTh7nqUPp4BvWlJNHIr4K7cmpA3QhCu7l0PH/zXJrEj+c+TuCh2
/BpwX8lzC+bVnXcD/QCC5msQ35VxARycbEFDp+xLqDNrFspBhCIFCCc+ZaNeIO6f2gOqeMRD4y6o
1O2864nGEy6Xf6BnTlRYPmnx2ENljBs6cw2kzZzXgVGXgD/Y8+ue44mzpokugqFTPHDFg7yS9vfD
//tsMGiMQRfvC1aV6VrAoUGwzeClGE+NQ6D1zlcaqOdSjN6JZj5jbJ+/gHrozxqu+FojCg4wyVLX
l13G2KVOOKoVPD3jVWLv9Qa3cTwGL1Iq7uxrqjTREE8Q9VfpJovlbBv0QRj0P8t+9z452mPzF6xb
cTykzq74TSjgz/MFPeaxCBNym8FVYnXg7MjwoQ0+IPLQxqJvPRCMVTjIogVOZS9gWAxRO3LvGVch
Dr/YWJSY6jpV0d6/UfTR9R8P3HALy+xWkLaOn+LIp6I67XjjVNm5acTZCMY5mzn1PZZ5yB0fexSm
rwVeJzknNIJhbxseqf9GRru3u5aJWkeYhlT02nTg4z7duQkDJ/LrctrAbux90mMf8JnmQwJjDpNh
jaW761bDw2A1u8Uucs87hPuhbllJZpkgkp1CN7S5PXF4JRF/7iNTWCKcDhtU76UUM0zTnh1Oy8Ic
fEqaIEju66s3DlUwnQv4XueOLwzpwc0axM72nfH5RiVFnmxubAU19hGdEJbj65qjSReKxNCF/jjl
/+5gFhFgjZMidTRH0I4vn0cU0J0cxoP9XHONZI3QWQRkgbDot2njyHx2gCcm5IcSr1LwrdOJ5W4e
r0c2nSIl1xo4seOWvj/nkSE+savQliryuky2DLP3+6IsrLjdXEfOAMWvg/a3v+1XKwBMRHIRkuLB
VFEvRlrYra1yuPjsfty9NRLwU94ILaWKHnFi/Ekh8jrDNo0HXBoJTwVR0nmftwDeqwTaNExpIgjp
bmzPpgyY+fozWlm+7LEwerkmbkW+4o3gcweZZza9LQmNADif/gCAumob2MMrkY1CR13fGwD1oMs1
si0lvj3eRdEwsJiCA04tRKXQto9znwYTFYJrzcquvZjoyye+Wtr8RKIdBpdOUe8F1V1zA/VIMjI5
DZe2iPd0o98eN1zzG3aU7ceAUe7Md5K/Gj6706q8FNmEUNsYDDhzNviPoBYXvIxMyaMQeFLZd/nw
5/5J7b2VEZHH077ynthueklzJT6PquW8NN+wFjv8RUMjbnNG4VB/YYNpG5rrCpqTRq4VNB7ZXlqq
yT0TOS5lV8E6k8539zNPE1s9nY5ZnK1+O1ZYHlaqbi+RpPL6iSLbgW6WCieOr2S+GgDByUPu5eZE
LNxiK+ZUNJ2oVdPb1P19B9hUG9aWvaUA3joGHwOLJN3+bzSlbigYLFtsDxI+bOPCEx8L1rpzWicF
3youDECYhadL+4DIlaSxjC8pWkoO0fGrPfjb9AbaUOoVRMMesNrhlPLX59bl5bplNWOgU4dyn4CS
zj+0TpjHdecFsKy8s5NyQVmTmWAOgWS1yrjEbzbUH8Mhk/URKy4YovlUt/zYlfvlK69fgC5DM+wD
oygxLoXhavXFL8HxPevCm3h2NnfBZVkxzA5AAqN1OCP6wPaTzfZbqxnIMjrrf2cq+lY6gLukHDwQ
26jlefURu9JwxfIyW5ze35NfI/PJgrVK39LxSIa2Y8kZf3p8YZ6D83CqDCawZJ6Dz+HtAKHSZ5nG
qs2JT3P1OkbrHTJdNODL1eJ3FxokWjHynPJEsajZYwSIdJhCuPecKoPoAp7PeSiQJuR9IswDk7RD
jkxV/M3W5xIMqryeMTUuZYzY+BhPw5G6HiKIhJC2O0GDnt5NSI79k5+uoVL0SYf1JNoSrpDk3CrZ
8vHABaeccI87p+9JQ1Anr0Ws8QTHqzOfSwRfrcAVrbb529u4s81JVjv7SlrSyhpvDIWRTjcrtJ7+
m3M4jwLkNldVGdCA7UbVIM4nlAaIOO2Mz+oGdDbsVA0bSadpRPq9XQ+LMjFjRlhE8BXHZCrxM1vR
hYGDNcAJ3Gu4OOTzmpl6KxrGx8nabhLJPFLll97Vd07M/vZ8bMOa6G1Q0N7pDZ0GsxJNZibl/U3E
g9ZIX2UMYqMZQwSsHtQoo8pfC8zGNzDZ5emBZFzCNXKiuaBNnRH3N7zAtc6siN8XKx+9JlsPlFC/
zdDhkHoZZBfTW5xRv2hISY4oTtCA6mtvj+cWQ6Nw5L44U30XfX/U74FRpmqV8LecAi2um25ZOK8u
ylIcFQLbvkqLjUy2yhtZWkAKyqlIlrkIWjm2hceGr2MJxRNO8Wpw8nCLRh99RztSu1n9ZVNwcdcK
ujtFDLOGcW5Bg0HtqFH+v2GxUeZUIMFSZBxcUsnVwm5wGg3lHwQ8Em+MeXhiCB+L6a2oTONP53U9
DsdKSwc1wajZe6Nk/zSlZqfIOthJeZGoqWuK21DwSHVYuD+3RFTXK4jsN2CJYuUdJVstz9JKFnH0
vmOl/n4iOLhEDhXfGJwywSPTpP1cDraBRNEoVbwttAwiOa34oyZWsrEpopkVBjlXSqnZKPEHD0iL
ycgweeI/2QT4ylaSKcnuCMZL0Jbd9w8BTCNY+Q14h+NYkX5UNQ/NoCgVXWBt3j+dfM/TMHzsXFjC
/48Ipidw+FqjCm1tYYD1WktWiCCE48R6xNyaR3sjMCwYxub2gGrWFCCeHzBQVjxvMiUJ8A3NL/MV
aqaNpgQnEtpMuALipaKfdfvUU6CPrqOqzKJDKeHlhK6n5Sywpqyje/6xGZ3W7NmBofxXQIeb8JBb
m07YZwitoAKQA+k7eupWGUmTi1ePuVkTJCXIphsSZwOrOSQttd8YFZCdly5UeANTM9TVNPn4mx+r
TynS9Z+sr1OcEQ4+BhGlMyJr217eRL7ZWv0snjYDEVq7M0t9NbXe3WSMioQh7DHDeTOxyhXmDNeM
Gv3WtHUdyjRKxJEbTU7WI9fKhlLPOkcLfcFQ6inRM2iAuifyGgltgUkQsZNoJppeH0rT6V+cKfRX
G6eM7tGTzvsCgLlG+T23Ma74Hkv9D81/i2ERANmnSUwb6oFJ8xWSuJxb+jnVEk3Mm99IlVtVnXKF
4uSPMnBFmO3j4/10eeX0H0kjwY1LtMyjZwnTVwtdnWuzD/UB13n6BzP/ycI33sBygrq2/MFNBUg5
Rix4/39U/AZltdhtJ4lmiIx6k113n6+fXCvC9PuCcU+J8y9NJpSaOiH5jVf5F2RqtcetDg8ezjRF
EyTICCerI2ChlvPaD8MGJaL9BdOkFh3dVPRT04Xu5KOcMYkVf+iJoZVKOBHKj7KCQytEWrp1kbFn
vwY86O7e7e2SOWvFDVjle3HWa2AKov8qKRnrUjG+QqdafNVGEkrDww3qw6pIBGbLm4Yw5797+VoZ
3/RJEwn6gx2LZo27Q/I77yhKBehdHD1K8+7o4cYF+vi8eFCQoTLj8Y36pUzU8FA5QVbkQ/X/aISN
QuXl0nBWPxzEW0XoFdtw+U/xq5/heV9ybP1yEUU4s+bd0hYcYpscb36lyUBkdFJRa+vMhEh1Cn2a
0q+vMoImuaalLchp5j3kx/I67jy7dbmhMazHleA/+/TF87jIBd1PWBcwviVd0kzxpeVRv+ft/bQZ
93tDEEo6wKhwHLTYMbS2c21bOI9qVYvyNw8jR632oflgcW8Ppt+XBFy8s1LTry+5bA25ZTx+OaUk
qbXNMD59nUzorN5h/dAtb/rAK42DBs92O5ktBASLv5jrZ3S229Itq9t8Q6kjRASoForGwlaDL/46
tPh3Spr1HCEvFyH7LOnG+k4/Qd6erkTTlryrxSChs4lWk3Pg3rjRCWdedjd6IcFyOAQ+4eY7EaA5
gGmQYZXMi7l8BQQqFGn4azF/tSYKKjQq1xg2naAEomhAe6RoqWex7vTO9xTpIMmxP0OkfaRvRBH7
MQkpNaFVoPhzbHTTnlHsxO3du/LliW+f2eBpudFyHbcuz/lzZwYMTjpXpzLGbm/yI5bZ9fPWnrDp
/muejpL7NnzM212uLfL3fxFRYPfJPIri2WOjmFK0yMOpOsMegEFnRQndMUKPCg8vDbqULGoLEmSf
ZtQylQEBZyVbFvETgkRlMaDITLHIugA+VB9mzlVr3j7mQ7YjNY4z/Gi1HpNIcJS1046S8RwYfCnA
MOATYvFpbBQTSW4hJESrbeHei5K9cU4e5OTXSWC5EhBhUYAmC4nI91j2gvWC2BAUIvH5Cq5mM3q1
ywefFPtve6V7mwbfg7uMAZiA0zLXUJ0lU5u7qjUp98gS6ZuQemgwOu/KKXajcH/jmxCLK1bc/Yi0
2cCWwXujjhv6MCJwPJQ5faeWrW+78pw40HQldzhruCHT/tCVxs+0PwaIDSyneLVswNMlKfk9mPS/
I7Dclc+sZHccVhmilklBC5shVyuLksszH9LC9kuOxzZArlaVVhTq5AFMFtdcgExYhH1TaAH7KQXg
wTH/0ZbuM4jvrH69M7vgl5MjLjGGelalmILqsBDGLxconplGbNFVKi370nG9zCtpmIu+s/sn8H39
lhXyGiM0WWlfi2H8dhlzik7KYMWhkQsLvz5wf2hE3NZ1kozuWETP9VKvBaLB15BUJNWZZPE6MBf2
M1jvP6fK+Q01Qdc90qKglsUkOU5U2Uvk0+2D2Mxcneg8JkfPOAHtlU+bN4HyR7FJM20r34/tTBlu
2oHM1cR26v+yiaQU4sj+Pb9BUBlZwro3tJ3CSteQDlOh1HMlpU+GHTQF59haIEvcBeqhauLiUj3v
CwNJeoktt/69Z+87wzvLNz2hFT7lIZZzsbpL8wrxwT6vsXGMnQASE4xZFon6rJMPsJ9PTJGS+/Ls
z+6aSuwKjvfcG/PAPW+KDr6pFdkwmWaPYc4Aq6jJLKVdo3YUxHEs4hCEgxBXvmVgsVuLeHcxK73R
Ty9Mq9o7csTwbsgcNtXjMYANVcO24xLPuMr2u2L+T+xFCC2wC/5ZUTBAlUmXyJxRyEqbjOKrU0/t
iD6KOv9GX4Uq15ONpDG+bzb/SICQ+o6NPD8VYIgSU/igzBSnqn0snYy8oe+YQhxNrAHOh9tnT5jr
Ov8CW8pxANmoKY1NU+3sjGjRv9CXVj9GbmvLMSorp0yWNnQKGvtt5hkqCuIxg7gFeXw2P/ObMJZM
wqnmRZ692+7zsSktAWcEfibhWnCMS45fajqSp+Gklr4SzKhY9Z+Hh/OYzX2HisUyyB2P0P/4ceD4
CVavHb3rFTkC6AGks73kKSyndnoMU7NnTymP0Ogn9h9gxdqqjWHfRgQTEJ+BqK4PkpgaMHCzyGtn
xoDFsSEpyKvzee3yieV6ARbydfx/GyeCE8NYPJN19nqERP1bjKgRiIp0uYeWSLqBQ3RIQ0fLD7/G
PVni2C8f7D6ujaetvuAET5kTfBuwLYwAw71JOUIMnsd6msGcsqcnQB3U3E/kHtEpJU5bkUF00YPH
Q9BmicaC2li09MSL58Hl6KBAf9UA4SzmfwMg7TuZRqwX5PO17TDpnOyp3agpSTQfq32CnHs4P8Qt
Pj51aY3T6YnnULSo+qVGKOugHdNds7LOaSznEhDoviJ4hjATHPjxthwuzZdqLaRIS216nDt/QwA5
LXkLgO7+KtviesXxAD6t5+Gv6xwMkq8GRBm+GlkQAS74VqMdfcVY/Sbhacnzl79kpvIMLbECpiG6
8HoeytDrNOAiE+sEZJiHFR0yLmYVxeykxxJtoI6T3qPDMlzwRYktyjjTQ8ax6rlHuOm0VTW3R5Ta
Qt/tzq4cAOf/CVhrhRn82xJm9EUGaYEWO/2vvR6FP6tRfnF5EJET9W+DO36dLRsRYlMUkX/iyaiN
YHTkizNWkrV/P4a5v7kSS/kXHr0FqbHYFg28Y0U78RjpkxQ70Or2xhtCIkbx9MHuZq7ZToSAec5l
NFc+kuQG8w4ZT4EXTl3Sh7uLJ9EeYVnaCXrnueOFm8ttz453JHysyH5k2vec37IR2Da+Bx6jjYD8
pI0FAGHxL+cOS5r+hXgGwdBxUc0uYl2gYJMTvo6TBoRdzIwFnJjSW0zb1R4Kw28q3ZN3c8jBetBk
weWCXK6DU/3iS52mqNNIPAlNEDs26J/wSoBHqt5PblXr7rTVmow/cUpX9CGz7uHZTWorBuQrCs68
cwnycPzCvWvsdzwtl/PnTlkurBmIEVY8Xac2zOiSf0vQzUFmt7CLlOJnDdkBgK03+dy36so0f7NH
A5SJ6vsFX1/l6dYUbeZhnt6iZw+yDeGE34K0GOKEPWIYc1Xh2m34wfqTaeoOBQAzO6r9e2yr69RR
xjljoCsz+v5Tuy6FC9Awakh7gk8Tl/QGQ/J+sMwl1CBSYbaSEv41eimFQmR1NPthZ8/WmnJ8WFPX
07UH9BO7hfsICf1GCS9an579n/F1t4S8ZqpWvxyH30C6zBAAfIdvGSgHrYr0sLwpZ7yYFkPlABbb
RE4x3JeZVFLXfTodWYARAamCZXl0aByzbMXlobIUzhCfP09nocfrfMYH7tKvQNHkizwQ0125Dc4G
FaRaJD0iuBWafIbjQ1z8UByTQPmCHEwIUQLZZqlR/gNEBvH9CYSfqDlEB9zWI7yZPWXoHLTlP1Re
ofDw9sIVviSlYLC7Lq1iOmtpAtKZH0oPFYkbAM7mFa/dm3CHjTiACLTmwGo0f8W89XPA28uUFEM9
+nW9iMdbJTTKBa7vu8M/Co/onUcC+CCpXAwEkQBXThiiTS31LFlXWkKnu5xubtsPZ0M/I4KTJit9
tzeKMWTTHL72r4YBHlPpSYhs99zC704JPleZulk6XSGLLDYt5bqUTgDDd19agDWk5WKK4evnTOvw
WiZEc37rrUc8et/oJnz2nF6rJUosAXI7Map8kExtNbkNVPgNJLVfXJFop/i8EDJdi7gm0OjLVDE/
d65CLcPuPpqHBYdmt2iL6cNyN1KQDlDWjwdwmsbz13F/ogJF2hM2jLFyMPlVNp52TB06H7n9FDb2
XDqjUqx/ZY99oLeVdh7BI7sBsRbY97mBVrEBEBXhiSrIGOjZQWqZWOmLHgHPgkboYAxfWV4+i0f1
jvP7yZuZ3qeMtvmNIZdgzJT6+ziPLu8cEmKo8kOadbZCI+UxI7skLzlnMV7gdjyh9jVMpmODGkud
FSxeRl815WPvu+8eZYsmsNoDiqEyRG+VTGWm2XSA1t4XjPASscarYjfInmAbU35EsQfNtUnDNrEX
+Crwx4kGGEC1Q/9TYsBuLbhL+5lD8a1sy4rtCNqN7T17UeFvWql7YK4xtaJU1qeiXmqMyR7eJNSQ
vC5DSlxvNw7KAUmLOJ4KB75q6Q+4LFO28UdLG08fbeF08DhpE2bqY03sMKDoLyRYRHpdbE5854Gp
NeK6fKODHepQsc76LQmMtx6ahuBcwaOBt26XTPaDQYl0yspIzAVf5qCcK3GAf1xvqeMH7/eZYHg3
Gtkd1wMDAOeFsW0sfH7OLyVpHl1uXMaSPO0eYAW0/SsF3RI/pmHPJn/EGtuK4oxCR5od1ftNAwJg
bYFSHNJ9gCV96zYrlbQbB9/bssJhFDAFfZdb3xnN7FW26l26jDBAgdA5EMP5iA/Vok9ZpOS1me4U
8AhCXcIw9yjvC0U6mFV+icSdTJuJ+HhQoaLWgB+PuOhw+gozcOtJkAm6qj0sUzstKyMBBItAyAGO
cYBtIIl1pWkWjixyFqdH89MRjlkJvO2Szed9Oj152OrIq/t7F73Ji8vlkJLULHRvJAzEaw4QKFPA
YY1lRjkuYtYPhb1D4IqCgHKYSZRThsqrKUBEnIUM7hi9w+Cy6DtyjtbaEs/bMCdEDVQaiE5hWU03
FvCeMdax+Hb1w9+lqnWIboHB0BCCnBVWHNgWtxPJRitFfSLGFkUGbjHQInkeX8nRJshb4RdPDSD+
tIFpSn35p5tsdD4RgfPUEL8hJMC8kg6L/Z1quhpWScgVrB0kS1CxHblc5z6Jr6bsYoq/gcCGBXat
H3LnHFneZQqMrW41sdAUzXTns/5u09OWgolSzs1ilbsqtlzJeIiLg+Plna0HcNtrQHqcCAaQwWK1
eWM27nkUfy2/oFrmHUGNgjfaGJwBwlpEt4NzxlyJXjVQPK7UmSNM8YIYX7EeXR9L702mczhZxpO1
rCPt2sS1V+X2iLdSV+5bH6iB8IRw9UvvDF4UUuaV3reOFsq7dm2mdXb3idsVuBJnbI+WjXWJIEft
OUkrVoVJeJ317nMoUFC4UzE8ADVAZT+1dTbkoCaoqq1h4MYM8iz7Cg4es1Yq5FXgKAZeVRYrvYk7
rc3anfOzl8DrD45ap+3MjjjgZcrUN5h1btcKk2V16MdgDI0uuvwr8EedgWlTwbzi1BH4eBNTLAM4
xVCSfvapufO/VdUhaVMz1U3vtMB+hF1c/2frcQcwj5rHL3UzBleHU5maKyUhmKM0NbAoVLoZeFPs
A5v1u7Gz5SdPRvhW9XuYHg+8f7J86PHpx6H9ibBU7D+Tg4ueOtwCyo0Bj0jq6QPQj9bovGNiDJA9
k/Qcm3AOGEQHlxH55kaQOlM8oMAW4q8E3tjlFDLR0h3j3XDB69JmNmoj1XVEO5VsK9/ObIDs8dhu
Ushy6tqS9DqjKY8aqbv1eD/K3J0CBqSHu24eV9GD4lZRIIevpl6diKU1KX06LiYlBLz3xACSSLtV
+yNlZFR4lc8ZN+yP5xa8zwODpFeML3Z0kxlhKvBcLi8HtVERbDVCh9jLm5aZ8/SOb2+4vJfks0DO
tS42QoWNU/PXbZ793CnLh5hw/oWKf6RO2L02Yd5IlLfgG/+25IFXOjeEj+GV8UW6dWlmULtv6Jna
C0gHKeNrY/RNWnW33uD+KORVBUqgz/q/lIKQByhA8pf26EKuxnK1RlL/11S2AzW8noh1AFcTSFwX
Xbif3zjS7oAcgoUPTc7bcou1b5VFD5GWj4GzBuSJXaZOdQrFTwbZWpTE+CJCW5+ZyuuyF8IQ9TJN
nb5IpEGcvLTxVOO3plEWUetgZxTuIoNX2KD2sHlGxTZPONNvg5k+uIlRVBNXLDP+S26E1ar3yFo1
WXqt5bjVBVRLCvXkCC8IlgZF+UyIrNpYZgS4UxfRObfMEiGoKbS7Ol1a0iIfdiNVoYXK+TYPSBVZ
Bj0hGQ9yw22qFMYKrrQvEjaAd0q5ioez26LA3EXOqRZQjG+CT4OJC40INtCn7SCM44mkO6RAiZmd
4Nq+Wjuae7UtYmT6Un96BZo5tgUncKZF4nWOBXEGcBgQoteu5rreNH0AGJHALuGkH+SPHjffecNK
2JSMpPWCjln90ZPdeAc+ubg0t2i8nbAe4aLNChNPD67F8IuwpMq6h8cKkPTbHh6nYM66RK32kdmR
0JvqNs6h3PqylEtpz1TT0AwSpmkg+Y859PTHtZAnUa6o3Y4Vy5UJQh1UwDYOre/WhqF2jyORWXdT
JJZT1zfhA69sWSzBLoikmfsUqiJTCHYPe/1xdQ/ql2H22ua0c1Czf2KC+e6hazj42oMxwrb+7bbt
i/h3RPW2YnXoJ9gW8peKsThd/5uwPjNsyV4hOauJF4gmz/bCVmpeYxv2hMzZUyy7PxqRxBTuuNLY
Nsu/gWbfjtCDtLVbhpkbafIImqb4zh4zaXeSvDvMsjhQ6Xt1P5Rc18OA7djXL/L6zLr62NcwyY2Y
6WmQ/CLNu+BVsD0XmiY2xTKfPzdnNtyeRW/XyAHrWRf1u77/9+IpK9eRzdlqIFgf53AtAAAdqNXr
I5tpo/NXqK7NdWKdkoCYBTUAA0yM+880SyW8FU8JLsjB1HyEYO98+aQeUu+Y5bcldVkjHUJCx8sC
llMUqsLNS7VJvVVAJZYFZJoj6GEcBZvHzkTRwq6KQWADGsVpvAjFuZ9HIwpg7G7D5e4P03EsPVDC
HWjwRbVnfGkBZzgVb/hgD0pKhjASqrkXVfdBe16SphdCQP0NC0YNLTLlkId9wnE9q+ZmSeLfAkQA
wsxdFey52Y9ZyZ4ljb2tx4jc60KBShtO668QHXk5rG5N2JcNGb3gL26RIFbiS278PLzR6iVcwomh
F9/2uiY28EEg0vKtQlFcaSoUtqKhefF5Fmdph14BtOWnvW9UAyGFLXiEOVZXvMS0ubZdf9hX1YTG
eF1S7+ypawfHdXr//gfBs+Xm/U3MLcLH0hopf446cpN1biVLE5Gp4LXhp4i3ilJpWNTiHMG/dy8Y
/CsaseKYQxizEf4JWVP9wozuxKsvrmt9O5fqPd8++9xZG6vbWMxhx8Tl9OWcCMBj0H4HFFZ4FJed
pW0pkAnkpCDK3DmrD3O/MWovi+jIMG7UOwICkmkaM7gLdwRFtktPJurEI+rfMGyvhEaPBoiWPgCP
zpvTamBZou7rb6GySZTAxcN0+bIOj9t6yutxlBz65mc1iYTxOdgZiQ4Z8IphLBtn8c29mCaAEDBs
S0NQHtREg5z09OWrB+Yw/57HbEon2stBKxzn+WiPSEj/B+XPuuK6egKFEtUQeNjCna3JfIsI3Syx
+Zk7TXUoaoVKtHovy4FB2vMfYerQd/bgFk0O3GreD8WJpDmTlyHJ6MatQoagEOIVFi+34SohOYA8
AA3j59wqfPgPolMQd8tTIWCR97/tGH7P0AkQj7DYSKWtQIfojBdtjdUwZ0K2Nan+Jsp/zcmkjefP
UseiOs/8i01HB+4dzQCO9LqJlcM1mFNWtyx+HoFenHEVdU2GwSJWDZjsBHZpmFZXiSG7FWpvzSPO
Obu4gZ1G/a5C2vTKeNaBsuLqnc16IXJQRY9qkAxAHaE9CVytJwCQnDIRCLQDI6xXMe1cmoAdplTL
/7nXpP7eCYxXLmZGaQwk8hdQu6UTpOgggCMKTscb+RM71r5gQdSnYlF1xkv42JpqK/I/+ZlAphXh
FEvD43f6AIkD0JdNoT4w/rOO2X14AdDf0ypdAB70mNM0GcUrcE5MW0YgTos3Kk74lW5G30tbmByb
VyxImsBmwrUO1fY3i5scLrLgO6U4ja8dgrebeX9+2a/YaSyhK2H01okdTI1wGt6dHSReW09ws1Yw
VYiWSJKISOb9z5oxwipRzQE2t0VqtttKQ6L9rL0GOnH+a/dPk4qKXeU/9Rb7ehvRQUz1qEPDXWPq
2WUFdidBHLq3BD5rD79bqaZ5oTb99S/AORpbw20hSLziXYBR0T/UNsGHzQra1n/XhixDj/1CZa4N
QRGRVWreclMz3MABDFz+WhxpFFmLAU81HYcQPHd8u5M4fTdrTTN/9mKbiP2KOjorsohfwaeB64pf
VLYMdRtVghMLWlovNQlykeooGmspc9/uP/KNfminTCZZTkUuZJTG8aC1PB4vG/UqViAYUZ7ufg6M
ZyGXvGcnyZv9otHXxUCJYwx8fUeoBRq+JA3pUUpjZAfg9ASn0+aN/wHor+4C6gXGIoaRQbwdnxX+
ZpU6zb8FxqklHUHJ7ecFNPpypbgWRPMhvbjNwRKR6BGH8tWO0UQoE2HQBVPDIvzgS63Avntanuct
334ZrzVtl1fHyLNhOMNWkavdUdd27XUInWxjS50cU39Iq5t5DCGKkNsNGWqqeZps+OnmLWvLa5et
pRtRtJFFgOhkmxtuHuqfQwzuC5HLMTFwcsv0FbDGKwT3kbif5mBHIhaDNr0jOHf2XUCU7wnjRudo
6+85sxQD7Fn03DW4PZ+hTo/5H/GNIlCTNGS8Yx/q9lw9x8AEta6A7T8SPUzc56+GE1fnbrZPryWv
8xVhqfkW5o5t77BZ5yz9+z7wTIoVYp/G6I09g1F+evdO0U7m5IIG7rMinSus1RL6XIgt46256yQk
5eNFo4ctahaHVtBYbRo482jv9ZA20adxS0CF0RlTx1bGKXp1UurCPS/3W6aj32KFWiC29wrE5hXA
k2s95xMXMAlVIhwxMundUso1mcKJXKVeVnWKidQ3z34/kvxFRCGCcIzt0wM53pnyCWZ1Wb/+Dkpn
SoFNV1qOaT++OwHg8BLXiuMLwKp2yBk4JCuwL93e69G58RSHjU0kHhuuBu270rhk1uAqGdtRpKG5
bl26NCzObfbsg0RHwMbxe545xh+63cnhLqYVY3ePDQvwWHv6TB8CEnCW2RiJ16WzELXmS4utta/4
fVhhVf7c1n24Ii1bxPu04FRL2xvtwu09S6clJQy2qWuFa+By3UZTQGUem9fMG+zGHuqjKOrWR/zj
iuxvAqwQF2B5Hdtag3qeq/wXredXpgIXAjVnrrlK80tbeVqumAPaww5+lA9qKq2mx31pBkB+RVmk
bkob/vaO1fqEkV3YNit6FYX+p5Fd7D/Ifq5ODMNd/gid43tH6e/zsIb8T8UNi5teushT3diVnqmD
BjO4O2tdf/iZZykkHRDJyIKmAp//Zma77VIkxaszTUa/QYOIMiAd63rWbgga855cGXKe4OHw/rZ1
Kibn0EdSoaYYq77vuOAhZxJvqO11WPYzvmK181etg8mIFlNnWwHpuj00PhIh/fAec7MJW/r9vioV
R00P+V1/kSeee8+sX647EZMo/a6NHJMZ7z2c6jP4g41yTem1TbDtHl59gEtTrHfTBCgxFIXBFU6S
qfLdDopbZHsdSplI5AnjpMlBN91gwUoIrBdMoel0YCzBKUjlxbgpyMYI3etackmCcTB6YS+3QWQ9
izFG5EwI5p41BC1oUzxcmRVzFrREIefV2eIUv2xedit0GAZnnh4sblF2zlVB/qt7Kko/hDF624FH
nlU4szHyXTxZJk5wASAQMFjapEEPCYk9oZugnaR5gcVFsnCNAbDIyN4p/0KXD+ZK/NP0Ezp5KvAt
a/djFDg3HH9ircuz4IKBDO74GzwSj6EYBOmyJGMS3ZZ6lDv7t7T1h2JKP8WLh+dNVH6O+lX++a/n
ln6PPQFz5f/VYaHjDoJB5bUPLhdjUnr7k3dnew92PMnWD2zByJ8hurqLOHZa9M0oHPkoRiwtdY42
bzDpqwrCWqI352SLBVmqNJ2LeMq7X2F5SBpvMlikTVyJtwXDmw6ipjUVNJKr+WpOJO4dGynnasVg
yF9sUddRQFhMP0WIYNvZlH6dAQanS9S+sE+aNM7IalH7U9DZeEWnqnFiMVSbDf1w6Xylyvm48A9i
AI8UOQkOK3uovbF0EYFV/MzCwQq7H9+52VFl06f7/DivY+0bii+qtO7CpjQaC/kiLiW+xasrgtp2
hXI9OwEpmwhJ54eRbd3xAC0TlHAKI836O49X0ZHH1jV4tBIVq7OTi+ZSIlckKHHWA7l3Mead3woy
WLq/Pc5fmrRNCtyRlkMkldSQyTvVoRNeQebm2d7Eupa5+nP6Raltb1ep5khlmKe1HuEMaZB4V0Zz
lfuoNMcJtIHdkWeEbxfqxn/RU1zfw9O1my+YM4XeIDb51alvX4rpQ7fakPu0eRI0+oh6ZJ1PkaGZ
m4evepTXtGIM8xk3mwmF/FLNMao5330lBmYgerIzKW+4tf3C6qrmrCEKux5onV1nORAdKUw0Slku
N5OxdYUvpz09aClZ+MfgWZuUJK+7fkf7NDAS1rvE+h6Z1C6NZ8Dp/0eIYTIVN/7TA6GXK4+BBw28
eLCLoYckr9meVRHKcKLwHZSsuvjfma41dKgEWYbIjFxpDBotBbQ7vfeS+DPB2UpfG7PsgKPOq+im
YThGPYY8jT+T3eHWv9uxEbV35YF5cz4UwcTyC2mUPO2/KWx46Trx4qoQ2gTVatcD+eKjxpOzueE3
Pq3gCjvxuBXMzlouLD1mmoFyFFUi6TwSwPefnA2O4YGumL6voYx8IABsdtbNl6P1ViNTvA+1N6VM
zFPMnRJZ9n4To9MgzwAO3VIOPXxCKYpDZIgwdAR8RE1GS5N2yjX2/PVTNF+iBUwB4zGozT/Rb/h9
B+9IssD9S+mctdfXmKrX+T0RBhYYoKMLp+j6BrF2BoxRMHXiGC1zEuNURgnXjhYTUS8y2/SYkgJu
GblFGt4PRVrfMTdF22QyA2vi+CBklROQ+4k7wDAjKVeN40HGyib61YAsh6A+Y2IFqY5wlzVxKf2I
23kqLh45cNsA2ZJfkLuu9Yb1stFR61vpeS4Umg6qCpdeHPSAEqdrw/hvoUVwB/zETv/6VGRCQWmW
6hgp0csmiJawdgih9dtvC4c7OABXvsAWTnT2KdDzOb4TkiDa4sd4iS1HK7hbuiah6IcI5c1XBVEx
Xof09ucE5QNb7bADQu8n2oZQ1DkBgOCakGVU83DZyYoffoLn5iAQyET6ocia+3Mw8Sx99e5a17oI
JGlUedgbsfYgIoOQggI2Q9R2q2Ad0ZPADunZefL1ySJmhcQmE8uN3NFwJdO+FLsW0rW196X2OJwJ
uNcuw8Y9Uf6drfyjhk9iPOFvyzWzFwT51rVeQgo6pDrxHnnuH22/pUMGtNZYdObfLm9c48EMIHBZ
4ny/CvE7NhzVL/WXWr48XdPex4S2YVtZ6pBca9TMAzmrmedbXvoi2sExHEntSUQwrXPNtVHPQnTJ
yi0ndJ1/Cf4ZCHM3vO2YH+ItwLag43H6J8ZFDrU9jRoJYh2UZXJdpinIfjCwKyhnSA5Gnhy5KKcP
ftxkLnqLFa0pmSxFYp/xy77l6Pis/jpsTaXeVVk1JEnQqb7JuZArhNYa6xvxo3oASPLDuSHCQ+Sf
Y9RmR+8J+K1338fPh+F94hhwbklT3YNbKTjJmERMCzXLYvj37e6hvVGjMWQAoTYfVD0AC3H7PSij
R1VXrQhWaSio30COAEezezSfCwt4OpqhANt+WXHRCrCtR4VzX8V48YfND6IgNvy2EhWV0kl/jbbi
ahgZSn6i2XY+otXu+lgpoUHK5pgs3Fe1Uase99qdKvwTeCzx5KZjff4XxftYUPr+rn1umKQhDTE3
s5QOMyNuR2j45V38zpKoGtNUSohRJp5D2sLAQwrWDtkf73/1MQ8IfC0BtLjR6A313ym+lfpl/mal
nR3rUVym/0VYt9mw7qF4CTUfpWic4CMUZta4hjDumZ1c4zKiK3mWEV+Wk0oz/LtuMzq2BMlr+Udx
GI67jLPeufiJyXZc1OqL7jM6FLXFx7UaY3AAh9X1xVtMloc9y6aCJz+6SHn2OjtHH/r0Jc7d32tg
4vy1kPeBOym/8HBohDL0D008SnJP6RSGVEp0mks6LFXWIKvP+Ar8oT/NYKCwi36avgHdHTzxVPj9
XMDzAphe0OmDVlJf2YMO5SHcxUBVq5wITziSOwjSeKMcB9o94uxmPP+teneDF4PxT9YOM0HcS96S
bjhfr8pnThUAVgjsDHkeJEEPunn6gC/ym2MAKoVIp785laaixW8fZ/dbn7x0Xo0C5i2ojfTXvonB
xWDih8lzFTIeT+1blVphQxxeilrxX2IJWcgjO0SwknpogpuAf5kJwmAuSmxCfII5xIMgzOnYh4Cq
fQ8My6OHIIYj5i0ckHNqndSqgX4/L/RQsjz6N6GVt+J5gaBHx/MgxwW5wBRkTwkAuBxBUAXRl4S7
ApZCYwikUP4UoO+b+ZSwIKKbb0uHFqllFhgQeyT6ksPkSyfwrcuMjq3NUbGh2Omo6cqktjoqgGPn
gPOizYWEGGckNjDCYqzst/VHt95FPx6NFJG+Bek8kf1PYEeszP+EQfnHd88pXsLrWR7CJdqB5DX8
p8X9+RtY8oNKmQ+Q2XQSPH4F+RQG8OqzrIW3MS7JexS79Btiqq5KlvR4W+d56B3ThDJaY9qcoApo
F0mXu5MUFYZz4xuqzBMrImLGFyUwL5Lh1ppUfGZ6Mj9rj/5oeUp4uCrF1Fu1Q18WQyyPaxu3mxIS
c3ZUfW2KRwzx4VBvc9IWraCg+O08VmHmle6VCSkihEKtyn3rc5/ze+MPLjRcNtRssZ6tjxZKdD1a
JEsglDqWHUf99bXQq/pZ8ObQP3vDn2HULqhLrySdg+0PXW6K+KNNT5udFhjoN2Pqd+ml5J2eSrP2
gemImn1Jl2/vkKIQjviXE65eOrR9xtt6Gz+wQDOzDjkR828P74dcduDgQG8Zjz/1VpjOb6BAcphD
weurREFeMOh0A85aKP1uyWyW1xzVxBdCc+HBYyXgsB3yM+b8vFKlQGscLYI+tlSBXi77iePE4sMT
ZAlUjFw4oeUgyJWfk1XVExpe8fBiaJewovBBBaiTEh3zqfGb0aAyhoERIuxO2yLtxhwCB7xUGMqW
Umknj6p3VamUyl3mse4fYk1QlMojDMMYvAqwwVRQBytANsm3ECHWhub9CfGkf0J1/p3MqWmyFfZv
1CPTO2838NGvkd9Y93/KeV9WntAcIwl6VTyDwN6X9Fi6epNBhmIsPaEkP6HZZ3Ug356QXqo5JTch
mqtXlrs+7i51q0Vg0aYvrejmiQlmfi8QQOYx+73ivLQriL2NFg14pnRd9THRlbzpclInJk6SLiEj
PcW1w9nNSbHQTYPHO7K8gF+t0YFlk0Fj9cTY2dUskxcORr+ZTLxTF2V4SnERq9WzM0zcBzlFVXmR
KpuZtWx341wEEdsAAroHOKL0+oTGr7LvDARrtEncIXxsfuFVnosgJUg/4pbyizpMRmzRPWZmco2X
nrvO4hQ5ITCFc0mc0oH2N5dFstTwyloyu/RTfQVH+AAienmGIXu5WGCOS4+PvvAo5Sy/MEBn0ThY
+09MeKbwn6KTF+Vk3FvlUzESuAD7BjIlun7Ix/FTu9412C5p+HEwzydiqn5oEVNwcJGTi0fzAYIo
+E+PfARhEBwzEFhER6Y6MTo7a/MMX2TSIlVfIvVvFOvvfeWn38NwGvefx25m6F/xkw6Vb8i0ssYy
uG3Z9Ymck26T4mSB1cc2t2PLj+DVwOwN57k97SfZdfRzss3ZQhxv1WFXvAqeNkgwvMGev/rweG+T
tEr8UhEPY48MlqI1Wa5p4Ya8No9WShItCXAUwt5LSBcK9ZiPrTd32+3ce9O4gF/xz6PVNNgeI39U
tl9SZnNake5zWwtQwOzNquih4zmkmjfDBmoMlV1dPk822jy3+Tn+tUj67vn6ENONWDadHNtEkcAc
vYBfEeNfHMhnZZkxQlk3iTtcMbZaycJqipspnLu5pmjRCEBS0CFt1/d7NTILon+cvh5GtcPdqRVx
0XoxNlpHoYp3Ba5LWwyAHCOitVBQHYOIHGvrMgrBHYFNM/LLC/mKqxrGbiTxM4Q7WB9qcU6a+SJ3
jZliYZoUme1yldZQa6B/mcRCCqAoBnLzPIvfmKiyb/wYvBLClKWvrEQWYwNbNl70EzpmGuFDrLlZ
aKwudA+KlcuP1iArXX5thMwrXEEfK87j44l7WC/SVH0pr/XrjjNIFE6cVy5pxA1fE6cMRstEMWrc
hfubHwlfYtdDWbs4u7lGgPyHtpaw8VM3ajhg/DZRFHU4h8gSSBkm93mG/0bItFqpNTMzuSsw1Vj0
YW5CksWrfPXYiZ/96NZcD409dMioXBYwp5w6BuU/0o5OOAJkdzcjeu201ncwzVsmqP1hv0qp3bq9
bjRQH3cmzLE3plqecmpuOUJ4PFeXuCvYG0Py6UQGTHCowKRzIYPRt/4PJOCJjy7Q1Wjvh2TJKJcp
2fESFOGFJmN87sYE3+WKfjwPqqjKec/P8ZrV3J66tQU7NTP6qwF+xB9QWWj61coSFMsigs2vzXWb
KvInqOalloywn7wW7rWYeWUALwXLmgHv/FyQlDAsu79khoxQqHlmY/q7tcLN53liTKQSCkIcRj8u
193uhKJRiwE6vgH3U8zMEfl0Yev7SoqJ4QEm6iGRxL+5eJ5jyYmTigoRB2FxkagRLEUJe/IFJp1o
6oXS5w7g95rRTTk6bWP8cQIUrBmevZpMJp7AuCaZdqxyq0qzlfrdhmszdwYAO/rlS82CbK+btTP4
PJj4l0P5DqX4BZ2x9TRPTXAQ7IveUFfb+SxrJqFQuhHDopk57rDzdJcCocpSEQSuP2Sj6GqFXlIP
QJv13qtjrGMG5ozWtyRd5AW9+17rlHEG/a8CJ8hcvsadIkHhgVYnKiXE9WJyzQQkzvhYC7udSED/
qd9WDFNRpj2e2+G8omNOVND6A+zPNo+W3knZfyu8/6lF8GYJLgyQgpY9gexp/Cqc9Ufo3JDnqEYb
NazM0xYY+grhQiRoEgDbAppbXOfNRCIZftIbvpB19XnYljbzLT+SBAOjYev8+4Q/YwdGUmNQ5bXI
iXsZOHF1+tUov94x5Mnq+bcjTfQf7SQMDnzS22SPAGxiE5eIj7c+mi6grnTx2An+44IkcB5sORVp
CjV1mMApb41F+/HE9GTKIE5WVENs5jzwU8pKvMzgsVIRKkyWokECKt4pYP3a0Mzjt4TY1EcnXpbV
2I2DgM2gZy6mXOPj65RUR22Qs9UJ85ftiM98UgMwR02qAUMPgrhHJM443UIpo2IyMTPOmUugRmuK
CU1VVZzqrMgq0QWgqCQhBHmdX5RTUGV+H9FGmw9OJ8BpEW2H9pGsHzZ53wuYIF8eOcou19Dz9Mnf
sRMeW6Wn5ma9YqG9L0LlgWfS5Y6cgk/96ew/kKzSkhPp0EBqhpSRfKfPeOIR0n2YYsp5TavfqKxz
zOEokWJ1Aw1hvnFoyJI8Q97ED/dHNi9WoMuC0HHAgPK4rt2+SZmyfWyIKU1BP0MHrnR462kausXR
941y+sAWsNSxgQ5P+/N/obLzGC2Q7DQWoX49M/SnkjctdNY/rKSrKBZtmav82ykqMJWC6qzLq0iU
HZmP/Vxk8TTa8dOkZ9ifsNa7/9oejbGf9ToLcoUl1pJLY8QfBY17opmigOuti7xD7nCXmrcj017U
caOFfqxEPMNhaijR6h7Hu8jHSao5X1jdj4Xrge80HEb6+NPc2D0u5KtvKYCEFrDDNnSOMUNXKA0b
aO+IS8vvB4pXnY/q0EmtZXMVfrFmMvnHTPmX9F0rFpsqX+j42GjQ06M/iRzIIk2zR2yHOVkfNKmc
e7D/mQn9oDszj+DnUtOvfY5hyk5PKUfHcFTa0+ye3aKyGkfR0xEmI+UsFGFtavrq0fdTH3hx3sLs
mZo4Nkk6ZvDEiBiJ5CP1vu011xpfbwvd8Q77xbs+yLd6Gw+h+t4UdRJbsV8di8DpqhmEgbGVWm+v
KveEqoi4kwLNcQQOcM0HDlbmsfW2MSuTSh88ISTLniy2Vy61IFDvWxYCdNigrxS7doOVI5JoCTgX
+uDp/9Duke77GClA1fYbp502fJCZ51TTiiYft4/3OGdes5o+hLtx4uw2vZUhKRfSnl/5MWdxe4/j
fE5VRjLFrEqa6lhfp6DJpadFOOpZ2eU0MICJmHqzSoc9ztO+6p3WoMcAmfVLICSpvOLpQ+7UTO01
jml8ffbkDuaOCmZ7rZqQNjq9wPV8FOIGuHHmdODYkaYzzGM9g4EVZ+C/inI2ii88HdrJ9rOoqBLz
5TWHoHoGwUDeAPmVScSv8owh9HIDm0yF7qSIg93VcZHAn2WZf6rLIdp71LCnDnIc85PBCRYW5g5M
8PQGlLWesKC8olUxIj1i6lYVUuCfubUlqEpOnTv3yQBgXGnD4Ru0T2guKDFIP0UVISn4hZejlIxf
l+coA/kiT6RrS14vPoEK8bRj/0Tx5s04/t/QeRcYVBfI9JN96Vt1RWqg3bRgrLIXHFJ+ToqxfL5D
QU8cy9dXgvnx4KlLnMrKUDU7+INaI+nzZAQJ+/komAFaUKmqELh1fhtBCRfc5ITPi4ukZbqmpDsu
W9gmQkFpGizdmzjktrJN+7GmmOZ28fRDypfX02jkDe/HapjMVPutchCpwCx4DStZS9H8oJ6Oo9it
m/WYd6msnCUNzlbfG7OcYcj++xVuiIxlK8Dw7sSmZds5k0TuKGELSl+DTWhLni37YoX0AN89IGJT
lTXUrqYtbiIguYQR1efq+S0z18IHoFRR/usPBkS1s+j3pyMzsoPaqR1PgPVecq+UnYRYXuk10N7b
9szRbmTRhx/sbZVOL27dpSU5BuJi6mmKK3jOzwZVYFvWHuh38u2xsqJ5xQcXpaROmALcLygSoUv7
bZe1mjMgQMsmesK6VsbFMpBlr1Nb1j7huk0VtZSh4VvmKxpb7v5yXDAxh3K1YOYUEzmznERwkoHf
S7iBlXasJJ5Z/IJVSHcWc/A8KZ2V5jdx06a/kTZE40CvrdCPg5udzx4gy168BU5NSSwih/XgLTl5
xu+/U7wLL+qEy1J6sUC8GVj+Vqv7QLtr9y/JKjKi5UIfaraLbWHV8cTUwR/8wu3LLIhLUeyWKgiJ
2kvR91sgw1ZxPBokIteiGi21jtS5JvkGLADGY2/Z/cDKQHP9HQAQypexx36Ubj6K3fJeFq2aosOJ
C+GbYH8vHPiGf7bDfhjoGiK27t1QEeL3vZUVmEabeTb+KirwRW1w++RMFc351nNWHtCHcPfs9b9z
kMtMP0RWx1QQlItkZqUwyOJ7xMuNnepke58s9mYvNPmmNsxJqVL8xyNQymGn6Q3x438ubmhl+/Vs
iMsh+k1AljzuawB6fobH1xZYXKT9mxOOyBtZ9HTpqwp6ztxYiG7bM9+TjSMNaluBPFqosHk+Fqfz
OxANtHp8uw0Qwadz0TpWVXJrKG450o6Sdmc9aO1ooPKQBnimEM2kBBAUKinM6Ct4+wXSsemT1t4O
KhyYvyFmrv4CcKdjGnlOSB48h64VRj9OsSHMQ+TnGIoqbGupiXe+u4zKZ5jgu4oIgDmTjA6H0OJD
mfGknO9Bs1oZm1a8da0QxbOE90IQvFspYNWi10ZIQVRghGWR9vInH3G5D96vrCvUa3fEZFNAJmH1
td2o7BlWP9QfoVNS3t6VkNvmu1S7tOsh287lbIIQl3ZLaFLBA7UoV8I2+tWrw3HfaK84+2RShg/t
jZoyKiwHFpU2+pFLeti7Y6NtSMltr2BRFXatAGA+lfXWsp8akrkNyClMzPeGpFnKHYRm0KLPtDe0
I6KEKaU0hEgufw2LQIxwftVmiSlIIS3lf/j/xeeBk4nfmjFK8N1maugjLq4O2sKXSMxDXAU640MT
aURM5IXXefqopwD7smF9lxR4zhu+xw+urQkHYMtf1HRDkdyyJIxaIxtY8qR6DW/2p3xZkGGgBrLB
2m5rCzds9jj/MsqfDv/frf+zl4c6T70raVV8bDlCsEh2dWnKNk5N/XpyBRf8k7hrpo9iJpY+c5ow
PYo9fH4vLC1rEKlLpXGf9HKIdqyA80fxNJ/GElQhtGsTnKR0qbMy1xcp4ShyPOUwM2CVBnhTl6s3
269oCNhWWfkEFM+gap49yP82WMzCrN6UfKMPcZP5WU36lrnhcy/V7daatOY37tRwg7BjYVjpd2hD
YhusMmCE+9iC4XWSZf0wuIpBJX9mDsTcDUxr5SnP2MSrONMKjlpp5CxC/ECcG+bI0fCmzDpLzW37
wlPFThcy0+9HEuMnczrpzxbiOCXtauBs1dLtnrpEohNA2+f4xaSgusrEOkzYWnDEeeufcncpfY95
y9atScwn6h+/9W7RPziHxt83fX5sDP1yrsPUgscIFAc/dzBEW6YH38q0kEN0VYwDod+d46m288Lr
jiJmRLJjRR9D1gJnGx+Uvak3sdFJDN4XOmIUCn38KaAN/v2p3KLHTJAccD4f6p7xXd93Zboq/iH5
Um7wGVNjcsPQ2BxSR8qM0z06tlqSLLrTLDFj8IP6NkGlHdJTM/8QiaF9uYCDcDG0eM36N2GNhgN5
3vkwv2D6oEZRBL5aAA31gTCqKvrZFl1bdRubflOrbH09EVz7EJ5CwOkgY55FnsKAtnEjoIJ1rQPO
QQTpl/p3NO9nbsXIDQkWp3yihQzrF4g8N8Zw+RXTL/o5TL+pOw8OcDnlUapx3k8qLSh4GI8UFJLp
b4fBmwUElpJPnIiYKTGioT8pTdiG4Pe0IyzODBXZ0mRUVUrhC2U/AwOXDVRtZcRrBXP3CB61oPzm
QOuj84e0NOHv4SC17ZbFZZZxJ72YTrBQThqLHww6BM3uD0bRuJWsMX+luxpRZPATOn+XUVeNWb62
GgSQruBqZoK161uO9XUz1G2HShM10GNXX9Sezu+NPcWX5T97YKAqJhhuxGd3EYlOy/WsggYDUNGT
SGfN8kO4Uk3U0nyUOJElmxN/e8hDmwsOXVc1BjSFSHQZbXAlYXaUXzo+2/lF+EVGSW1vZvqNBl0U
Z/U1tlI4EkvCxMqA+St246olvpWjl7LkdMLS4VfmO0pJdV2KXrJAfZKM5M6qH1Zn03kvSkCjf3Ty
QX210xLJiWk39fSiMqZmqyBfXgU+ijczrJ6vILlYwuaQCtG0vbGkqhcsF6xrmlGbV0GzjLMuEfcx
scjhnxPoVq+8+cihHU5DSRqWcE6gbUBSXFZJv37nX2v2ViGXJSe9OGAbU1N887daDXselM8Eo9ap
I1yD/WFgG7QP2VoaTWdWeIHSy/4iGZzDjB80Iv/EDnf1ip78HwY2mDQc0lgMFKJyJuIqpaX+HBjb
n4r3B0xPo8hgdtcqiSLQZcRmMOaNISXzj8Sxz2PFGs/8UFYc6OLB29If3bjFAkkPxS/vvFShTBKc
pIavZZkAZ3LGBChr2Y0O/912b5XNTItxQhdKtgQxr76OtSicfTdBiESYeQSjkv0aosBz0NL59neB
P13RUoSZAeFyAT9v4uL7cTWavut3Cb2zKEHA/2Tc6R8zTB6GIGyAOm3mqjYVnDunAFLPIHjixy9P
C0BFdSnTQECxesEeQD69lsroYUn5h/iZWL0sH+NzuOrkVzWZzjLRWzYriik9/lwy8iCn/6fBEQLo
uQs2SDf1kxIJT0FObHVsAOIHtxzW87ULXp3VGBCOxTn1C9qCj7vNHd1RZedNFy+eTXygwP5ibpZV
SYZ7xBSYS51sqSW6bfh2OOuNPZwr4JStjQw/7f3d8O4DgVMemaiRq8v3VzjtGVlLZqLKlbQUghuu
nzaLYkOENY0QcRIlcQlrtbRTtD9rns/Z+zKezOmKj0nbYjPvQ1MM54RbStKVHDb2/w634p6Wi8CE
YHSmlsVg436s/0HDtD1+nL1YmX2PJ0GDPg9HDWmVTcedyZtR/DraQ21iHJufZWPCHDUiVG3SA91f
L5yvqlZgUnu+RcbmCR8VMOBvTXX7ZnubtuEDcioh3uG7JIvuXQoCYeEjjjKO0i3DLZXWBuLNOjr5
+tFP8G9cuHdWdLqr6i6VAWWxnECRIU2gqZA/dsthNidMfAMXRCo9ssiAWCpa5lEHlrjY3evxF93F
tKlhLxP5YZui3rOOwDtzovmYu0YyX567XCgEVJXTpBtp+LcxZLOqNnpjXWwduHwpS+8ZH404/GwJ
R+b5D+bkApe2NxLEKgg/T96cgUUqLcxcLsHjGQPstKwqrkorRMHxquEeamTBZcDaRlf70SecTo6y
wLErzKo018pm+FpcnZb1FJLuuulTKIUAQkb5Kt0Rm8qdl13Ml4MIMi7b0iP4BSsKLeLvJcN0uxrW
XKf+SE3nrCFe+ZgFQwZTfL83azQPUU63YPcQnNILuAXHMLYenYGe+Axt0nZXqOwT5M8FVzpst/Ez
iBRa3ldGI1O7RRNYMGqIQn0WFe/uODuDzyxrHFbdTDIXz1Z2jOtUTXklHZj3WFuDswxK0UknlqUD
3N/4u3A2ZTfPGsPAs9RzZBxCaKCEW0/s4OJLlMZuixBeNSej+T/EYBRfDRzZd1XB6qrkK2QcXyQs
8PYQaFWNJa/UPxwMKKdMiurI5b9xaycUwGB8yChCoK/G5mOUFgKE8tyduyzwGKed3hCkskGETfCO
S0Ep7AHjWB3mTmXfMINgZrMAkwF7LYCJHZW8aY7eo8emma/FB7e52GLdf2b/JHrsnBZsFcV+nBs9
eAfuK6ZcGA6sFU0Gjl1TIlZqiHK6oNgRR1JqWhrP8prHXOGv7UM+1JmmCPlg0bocYs+g0EV7/EVW
VG1xFkSroSm0wSbCvqqU5gW2VjDJ0thXQGYCzZqldEklPefzy9n6Inc2C3tXZ8SM16ZvLSXNSZSd
w/ePaebJ7vrumR2f4Dhx9gUm5qeClwYwb28tM+OBRzsVRK4BfOO0HagxEPlgwbzLV56EkCeWht3U
2zYwkGiKoG8WudbQOlHqCgjS2ut3Ku5XVZ8bEyguhgaEEDhT+hBgz/ZzmOjF7/tM07lkELnEbWwu
a/DLlkHAf3xOO0RFwT3iVGdg/YXuPXvTTbJ9U6nKIQgW3Uqgqy4N0amW9fN3e/dgcn/W99bWYUwU
5/GQeABgm1CrK2Ylk+o9x2/5nx0Mk20vHj6TA5eLrpB/xHtS775dMGe+s7xmBXq55EBYOCHJvtbA
qo9vNKELyI6iiH4xshueqmxkhDTyJOzVS88u2EjIQcXj42gF52EI3OVT6k5qMdVNueNj8sPqMHQB
FZU0Kp0cJGgXUw0Vquv2LUvLEgItu/m7XJcENoRi89GsQvj9wsbsSGfLytjDwKHNjkjnEPcG2E6t
U7etE1Z7ooSvmvhCJQvz91l40MRTd4QtVKSwmGzCJEkDSG2ZKaBQZkvv2X0UsDF+IscqDCGrYv77
X6gwE+rQPmw47G+vGaIMYS3KinRo4bxN8pPFyp5CzK75EIIaofiFEHYZFDXzNHn0gDGQ7I8hoEBt
DNpkYnPAOGK6Zzhpfy8aWFP4mlfN/Iq2lsbArhwIAQ03qcLq8p88/21hLu+/F9Jhf3MGPbfiorc7
1W38mIifXG5B6KlrKzMa6Tid/ukF+FIvTY9othvjXA/x4pobVTyimo8Kvm25wUWXM9DT2DMdjqqi
wV3QQhATsFrUVn0FqW8jJexMmOQMfkFK+Et5d2vseazW29pa0ug3dntp8HD/n5JHxXM5jvWF3pzF
Jqft/vVXnpD2Aya8okLpAAaiSrL/cPJ6TvIvsmCcCUpOr62Hd65qJdsdZ3MMJS4iMmj/QZrlNSkn
wKFYU3AyBjO4o1baq+Ho4TP4/pILz/Uf9q884Q+LLx93w8kT6LrGY1lTxZMOD3kQV5P6lmjrFzjA
BpOjHgmIGgMs8ALo+wg/oe4hHqgv/8TI/uqbxNUv8CyrtxyjZ740ZAUIA9T9Qh1W36BOPo1I6uTD
y13HF6o/2wgU5kCbJfRjJPIPefhpb0W0vhqRejoCwyQpXO+yoWb0PdcG56EfaDAeHPm8QV1+Bk4/
HYiUFCmJhUJp8Mtqcnpp5MQEc2Uxq66CXd13LPFVrLBhllnDe2+Shb7kFnaZVPV4KhsF+/tp0r6i
zCMAyCN2oc1IOdJazuFaqHU0LR0bEewo2qp2kYH57Ola6B6+SQxp0p6xDTxJl1V/qLvXzQgY5TcL
DRPhqfe9cMAPisv7MBng0/kSuDcs7EtFAuz9nVjBJyBDyy8QpvoPQaaJFdZpHBSxufoFxZsgLZOh
dR5B4zLHZWYHumzRWYBKyU/lrvvXmB1HdmNXAtLshljI4iqO9Lewd8OIDym0gaFrhqq6w/pru9Et
gkX42bRZOFmSy1H1intu6chbYK5HLedcLcj+/5eiiKF11T6T8EJ1wZJPdKVD55wNSU0Xv/t86Y3H
5UsVl86BhlhCZMGvHLeKH2XActPmPWf99/agzvTDC95uDwMNpMPuzgl6p2aSwF2Lb7J9MZtprZQ7
4XvZfNgM/jtRUq32lhJSEiHsqS0URy8WW5R+sy/3sjOPdnpzci5ezckJmi4lHphdMSndD6fj4rnf
P5oiYjrLM4S+xhJ3khWw/m9syyc+/VS9R/iviMsYE4ItjhuHIQsp4ERcb1UiBP4RSpmW2017uDLL
AjP24wr+r+GZ2bdVw+G4vftH+qzuQNHs3Qm4v2hCrpWlUXxMjPVTqSAL/5L5ojY2BRJBs8Q/Am1y
/luuGUldO1wFReyWNXJgvSypZjW4pf14Q4hedRrOdY+o7dz8KmnVO8k6PF2dPs7Z9BDsM7kpfdXn
bxznLmFV9mVoQgilZgvPNbfeLk4+N1+DskZXzLHUUodliu0tKsy+YuyxdYr+OdJS/8n9Zm9hNSdU
csq1s5TDZZbgzLvxe/vMRnnT1y51W9ReOkFKa4YN6mAQk/pEWxBQty6aK/7BhVkBKgpkz4zYhoBX
szHqxF2Wst2qMf9K2zTX40dMv1Wusf7oMZ/qizaIaoqhNIuKIDpJwwLTSTJ54eAsA5B8TbYwsmMT
09+dl/AqEbRe1EMvXdwTsNy6Joa2clWg4CuHkKvGSA/iWHRHHGXUEk31h0dAQqp5cKRIQUet2Nrc
pfB1HjnOGOIcAFs46w5g/DF94Mfsqh8yUx0gLI+y68YznbNPB98firPcrYW6pOkA5yYgyUT0aZzJ
/20+WH7wsprlbPjE5OjLCzRZKyXxxRZ+h1sPoRais4yG1sGVHIkfls39ym4FcBKoDLtiMmihwlTY
oBuEdy66AAegh26eWJSEVOtZZdEpJpiWPDt2pMNwpAk2GudQP/zlR+WJebScDVOnxOCH409JUWwh
BoW066aezmAlsxITrZdpllcgl4pUi3yX7hjG1q95zUFAU/FVi+BGO1j5FptM9mnSXa7QcLBicbB/
jrgBn4O3D1nyvPCHgyTMBVElNGr4LAFVBVbwscz7ujaHokzuNieQJT4zz/GOwTnyzZaXYkO5ZnBW
AVQQn2z1G6mb3rmDCfHPNAcfcZtiE+7UwP+YwVN2ObLGsdAQV/bm5BpA/5eB5uD/FB6mKxGjyoC8
yv8XDoh2d2rfnhU92O5CQeKCkNlgssUn8D6vIEzNK29S+zYZ//LW65xxY75GnSmpGk6IQ7vph1X6
vTCKQCBUMxwuJFnx2VLHFHsRboD31MyVhL23EDQiiUtzpgvE32fdtEI2BXzol0ZAgHWWcSwncQ5p
TzAZQfH1MNBTwwr5S9ujTK43gApBUELlPg82sXxft5krQIVXvfOukhoXVWi47Wf8bs8pT1T7GDGq
W9RFhWyvB0akyT9e3PNxFmKHmfO8eyUy1My5rxX8p4bodwtnr9RHT7FVQVRKrY13Af5H1A/FFg0o
ifLrg9GeBv5kOo0+HEqWJWplv+U1mPfJFugwWaqHc7DN7/OuFxoTp1RfmO7zJqQXmJc5sJedH7j8
bnpmab0RL1TmQx7LmPwv3umSqlRcwJUZbJMyyayw8k8CLhIvSfwneuECeZ7QXA6PQOVtDVVRZu13
36aNIKT2pO5niJVhin2wHRwJNEZiRNRhUZVymUb1Z4DiRWvdGpzzVxoHL/MLZfX8uM/q4ihs8fqS
75EFoAdCn81uyY/YtUb9Urk6D5/CN7nbem1t7bUqvJL4vrtofs6mnKQiaDYNnop0Hy0KUjcOLhEU
d3by+jOeuT2BbDEKC4f4brbZSm5H2NJfiKXNV2VxvSegEKYYyo5oy0D84QWpLa3eYOr1bXlc0tf8
w21G3RXmVBVGBW2omDIzQsDiBlt2OfFPfAkhJyNgsv15bne51ay3R6sempDtCTUyuHK0ZuIVK6/2
163CNk5RhZZT71j4eoPRY/WztskGTB5+R3V6+xnOPV0qw961VrKKB1eypRwz6o3N/BZrEyswPCxv
OfDFnflKSe+H70iGg8MP6YPpJms9ly2SrKPvvLAGY3ql0xWESj5Jtzs8mxVFUBn1l5wRYjb4nGod
eF0Qw6igejUN205rAsh58oFP0r4pQ2//r/9SlYjkEs01ZKhLtn1F+3Oy4gU9uF08XAqaOX23KbWG
cpkeslPRHhscfYNoT7qDLEz/Bz8xNkgBZCvLmCxhsMWrAjznQ3iyZxtfBWtzJQEfZy4oni3rl2Tp
p33pNSX8XvM4F5qiZukYT+9k5ruhAv3XUTE4YoAO0w0pzeP66JbDSQjh9hqADI9ZugmpcL6QFYCb
ycJOHMHoBmWFvyi3qqfgb7qDdOdgQD7hczTBM6D6Lg7Otch83mIjGFiovJllfCUSWOiQPgsYlFY/
9m6yIrt7M/0OUFhiJzDuTDbLSXb0N7X0QAPwpA1uB5fzjK2JBsGybcQvM5qM2Z2iAtxC+kwjIznP
xR7c1hpXG0WrRmRbeg35wkTVahZgLTd7OoOu9RFp3If+BWoTxe6ISilyyCnMlm7TneYlGxJcGwdi
5FwrGvCnfvSp/cXDVocDog9+Y/a8/RRbEH2XriVbjhbX03f0ZojwLr7qL5/8MX4p6nhN39rHiA4m
cwmnWBiq0f2VSuYH2I3UwGi05sq4vxyschjifIUosMYRwQafiZ+IXRsZ3A8GFYcrD85Tw516d7kx
sNUi/jOkYonZ+PRwVeWym1AuxoBGHLXnzX7JjVNCth91hBAFJCiDhyEK6s3jDpLeyIgYWzTKhrsI
HmVm2oMVjB3t6fxKxPh11NCNG9ANCPnSi8Zzivmf4+JIo8QZCL1FYKh109MGMXgxpe/zOkaKirEU
CmdvsWCbo7Gdkv3g1xsaNZTs5lOwezoBYYDaxe0qgrlSKIp9/CLNZ7dcuUtY+BJ/b6Fs2qusn9Hv
ZgC/3I2EHuNCDGghX5+upUls51ocGcebL1QicABJ/mN+Qdfutj4wf14Ex7wolW/CUvSWt2hvPiCE
Mfy7iRz08uPIbUOOSpUMcG81rqVSgPKH8d0Rb/Yu6Rg31uQdHq0zkD2pNcnzKvQBpf36VF0AQeYH
9v/swdgNUk5USHJhr0ffP3wyBuoK6/QHjXdGOg6qP9rGC223DkEsQ/NA3r/LVzJaLY4E8Ad/qiC6
catwlGPRfZ3Z3qFWd9cpDPMcLgxppoaCPSQCRb9tfsLM7wYGK6ENgldr8WN6sCWA2BYzkqXkDwDa
7Kz9BM9mBGt4lOBOH4enxv7vrr7vi0BeYvUaZ8pq8YmC+dpG3HE1Tnb0b0EaoEUrfLVY3PCoV4rP
3dWgMXpVhvePe33Cks/z1pjMywadkGkjLVpW5zdOhF+MQkaMKDKJBLaDyHaAT9CI0rDpmuwYy/TW
A82dLNc9iY46pNDQaZs08shAcDHuOFNA7+gEC73CtMEc5ZB4A3G6x4j81HGYTTMbG2ffj/TYfipY
kISMxsApHdcEwnXNkoyGky00zCtgXd9S8gDGTjgfyc0BjRsPTcu4YCS3p+P4d4k8lWnP+FSXBWC5
b7AQoSUofNhgfMmTunydbt9BsrBy+TA3GYpmnHGypiB2JtQhtzOiqGtIO5drWytSv1sXeHifoz/X
fQJe3XWamGN/l69YCDLjqEhyMMDJpxKMxjgTg1puf8mV0tKiZ1BmB7i3ZDW6i3jntnVQNDRJxQ6a
2XTyzJTzvMeK3E0iy4ZsAm4NmpmXYirV38U/MLtU/BiAypUCvGcKvJ13dfPkMI9nreCH3fGZC8ww
YGM2HMx8OqAMMD3TGubZ0SBhnsG61DZbYuTvBqLwWdO52NU3yfsbcqZ/FGdtBnlVIkpTkNCCbi/z
TxW2/NxJiAplwKfUC/61P3G0rDH1D0z8HbeDCcSvNsevBaRlzYR5GZkZBAaow6DWj28bmKlx7N6T
bFVycyBgV8LffFB6Wvm/+xS5YYVEQ0WsqUsi4NJNBkkruMY1qnklqzZWECM2vjfxM6KgQTxM6+bE
77xWjMhm+YgIMIvg6Vu/GD64mLwKwKUMTIOEPv+5Fzpa7vvzRq2Kuge3y8SHp6pwhWHb96s55D+2
wdEcOtbe4h3WrqzirO33JttdsSyw0daUoZGjQ+fnrZsAcI5kK9zN3pYlhkG6+1kg9XLReXQ9FgGs
rb3Bpg5khXSq6GW1CswVGpOcvDsaL/J4Y9HWIjzNMz/KPh7DfnSNMUS0AnN3jLck5m4g/GcH9XY0
lBDqZ23nycDtEP/MHZXYftz3FiB7ka8e/jy11fgoW/a7XJbGSttJMYkJ5kiiFUZklplOiXm+Dn/d
CHOMH+jNOpQe1Okhi+iXLJTyfIxCNuqQPWFakjFPaD5llRWfBAhjOIpG+MhAqYCENHN+PPUpgrCM
rSqG6u/VQZ7J/SDLMBWveaYQpRuzGtKFnYVdlmMCwN7WncxfVu2TksTFS45RvpbTn624LB9ezHEa
DHH90gNB2TMA8dbulRHTLyco2BjxFBlpXgw6NFEiaZfVUv1xJ4omWjYOj74UROa1ryXUNbehLYcc
KZm3L110DTG75ziVU58qKl+Ca62IksGu5OzJEri2zifjlG1i0PYMQv0hfSHFEl2KVkKRpeOPCEMd
hWHfAiFOSC6jGiMCznJn+a1Nq6h4yEnwhbn6gzGopIshoaI5rMjfM17aAzqddkfsIKnX8fkEPv80
T9KyFSWGteVi+pyU0vazglSkVHIAvp39X2N0adxTDTX0tZkVuS5sOi1WzwZyqFdMfWf6detS4qtg
beyLlHIVaKoGNuMeWuhIP3wbtQ2veBOxPov5kj/MP+wsnb/sYrw+brT+tHq8YxB+t/mX0zc0OAEC
76x7NSvqCSZZ7pI2wf7YeIh+WT8lAO8Fg7XYiFeN23eGhP77g/kV8ZmkWeWEaIASjlrI8nw3R2rn
OdcNi7tHCoM3PRDXvzM6VLtcOViVGbkzXbyJoVe3r2qGpBuko3DMT+KJb5GaLVbo/eLeLkRZnT8i
67gNkJpEfUhijxIc5iWM4PYGZkoyZLlDxgVqtUBj9GC3cgkDIThd1w6CJ6vEUX7P3w0MWPFm6O0I
i4EiC3sYBnlustctqXTvHRrFHYiEfpUk2jsT35fjvtogmhu+GPybJDHsi2SOxGpTS+djKg+b+bZr
PxiQoUQwYyWAvUTisuhEuk1ZyelAlV1wLIa1/FhL5yNcCJySVDpFa3RNBsrGeEDm0TVUPbIKc8Vy
o6k8JFqex8o6Jcbk5GvNmvP7+Pulv9aLkq/tX7iYnyuKoYtUugicuuhjmUnH8rMvYCYrahJs5AqF
iU1weX5zivfziHZVfy8eDUnaTJbcm+qoNa1NQLZAbQMgGSYi+D0VCzTvjCQbwY0BtPF+xEGfTkuZ
bZmMOLeRspsCF7I/v+t7bik50PfDrUTG4fMHwreuTANFB5AUupvem0mvRro49i15LAWeyDV1x2zP
TWNk0yRAts0wDxzl7q8JtVogTEI3EN5vwgkukwSi+qd3l42FL7I55yOos4wBW9576ehpf0QgaepI
i+URsR8jh6/nMqpFowqiuH95WA1lBHG+zLKbNwgC4d8VkpwCv5fu3WQRf6eHkhJY7YK/eTP9OGPm
RyO/gW7HEB+1nojs8jzfFUTd0ab55jmis48eIK3XTCgKjH8OOnY045D4b9qNZTzcLm1Sj0MV9BSE
aoxiItbMq5dwv78jhn6lYzkLyduq5LyvxulIzOetz2CbQR3gElsQ1R473Lz5GYFw2qX+yjOu2vFh
jZvYz5ElA1A4laSCek0QQfvLGwtcUgYt2lF+OpGkzS/YPZrwljqQ0KqFs8Jr1xCPCyvqkdXwqs+W
0owx35hgCJOZFLNeX3Je1oxMoJE66Q7ruR+HD5psGqJ3ya553OcZSV7LNIAOo6+pRGZTGm84pVuH
If3Jw0qs5P85XJd62nL47rImUsHPFlFqBAKywfMADbPn9PmpK2ldI8ZYwqjRH6iGgt9YmKPjOuba
OOvGDpO9pHzCs9vMkVQseX+mUUEl9mdtVKSxeQt4wOu96fSrFcuacBlPWo+lJpfhcG5o4fZDjHQ3
0P2atvroP6cy39yXj/ClOvJBRplJjVE1FPVVniBS+vKiL607XhDCuqomT+Fw6kXOGq76tqv+AXMP
TZdkWFlMURGPr3ApnYfFO2g+U/b6v/umtc6W+SN26mI5laT/F3wphCmlgpejqMtPzRELxZzN1mHV
M4OnuXVeCHaOgxsQM8QoY8KeScOw9vNdSLQM0QpykbTLJOF8v04iTA8Ydt1Ph49P8Co1WgpQHtQp
yTzrlKvxWrbGjonvb64ZCPPXdnwdYlSfFtcFJcAxtCGSCsTLPvaacRpJrv+/G0tAzaLspdLSZ1GA
Pk7mH+R4YEAcgPLJmlK5NrIVDJEmydacCuNWTypT7OUBtRtPB+ah4/60aXhZtPq4S69172GsF19M
J2ZhyGIo+aiU0zK9F49oGPGoEUBxIM9qhLq84GZa25eXp6XdiBe6p4gI3aWTNBHVPHRZ2+sFdn3Z
KSOMOC8/aZ1dJGVVDOtq6ScnERxe23leN54UqkBFgwwbSgiA3uC0QfwUO8xqFXejJDZdLvytdCgx
sPfwvE3nz3x5GZHnJUShtYCukggPES0iHbgy1bbyL06JH/jhzkAkyYYCcHkk8pky8XeAPMq0KVmG
JlH1QhzsBuyslSMhB23ovpBMT1E22Wacr+6NC59tZYGLeY4cw5DaffWBhs2AMKI4KRjPRRc9qfkO
lx29qc+3q8T29veURknn7KP+Kx7xO6OuAYU8AWDlqOnpEtNRkrym1L1Pduu2ZxEz4pUv6UBq33Xj
17D/ZZ0ebQ0HCEjc0MrfzeesCyAxOkLx2/7dAGPFpS2YeHmLLjW2Q/LMmT9MtDaLRT/PJZO14P0l
ymMWjD1fSqndhdRjHni/smFzYK9UZHtegZQ6XdfNmaEzx8365udN/l5MNfjmD+sdWRqXKm9ne3s+
rF06X1vjXOSnZZTlc1+YDjKN/K+nVeemQKWgw22EEdkbuBWbVk5RfsWXPRBtzln+hMaS3stH2MMH
vz7SEifIsw8q8BJBxTL4aM84NoGur9/rC04fSMhU/qVhEfwe8lZw5sV2xVd2+DpJpL+dQp9o2lJ6
WWT806XO+DMPm+PMYY/+5ooKbS6/ykfa9rmDyDbnYSQrs/7J4MV4M8LaZU/Gsc+xuo0Ded6ohkk0
Eh8I1a6FAYwKmI8HxmPq53edDMzlga5c5l7P0qUOSTjccAglY3e62N9HLX/vBHwDDOmjr8qpZBCa
o3DXkEoI8/Cc21yu9qOygVyoa5uhvbgRl15NH+D+1pu5E5hwZdJhG35ZiQjyiLlCcI4OzjqW1XwD
lixGETaTBmF6riGdnT9NifBBEX3rJbrxREuDmDaOLoP0tLWHTsHSTd1jT0yTNcDFBr2u1i9wtlWR
QQyYthsxTZAM8zrkSjG6UwB04VBaYUdBhWnGt+3yH0MHI06CKOm5IJtJICMrU0iK/vSdZWBMOzqM
w9VZVDAHGKpvpETVwLYx3esiZrtug5RuV4bSLIVrDpsxV86JrL/bd32BtOLeUvLrRgUrQZ+oJLxB
hfLrPM9PPWqlVjckwe+Lz/IXv0cgk6f1hb/IUZXCwITOfDG5hQ2QjmUa893NQjaLBay0+WqCVHN5
sfpkZOGLZkltp9coioIQWRLm3A2oYrlo4nMBcUpfNZylH084pa5SO7Biq+CYJihFtSny+/0YflZD
GWqb+fRVUlC7TLZ2KPWx/1kF15npzGEtoHWc7qb9c5Sjs16tG7UAQEAGvOvqb1iD2nW9zgmioVu8
+eFqYhD/653j2esg5ALfukvOFlxz/nCo6TvSpSJzbN5J4F6aMRGfTwPQYOsFekfRc3+8Cyd2Zrxo
y3YdSoLeKDd4GWj964VP34FfQnyLJatAdJbe+Pwvlj9oLjALWj6LAd4EoQVhQGgaOeCtGyxWUcwF
jm196ndf7BqQ/ufvDsopsLRxRv25LT4ggBG1pgBttNgkmH49X6J2uUT50VqrAhSD1TXjgqm73Ogm
0tpJms+Ytdakmy4ZMl2x0vmUTy1eK5bTiUUehSvw4V2q0mx6Z8Awlc3WYk7uThgUZAzGOxtinU9W
z+zK3NZ874AyHecZmSHVQRjgKoup70elQr0TVRwTUgMFtMvgPTnrs5a4kWQO7brXdHeSKbK2ykw+
I2YXsx0VOvUqqLS+GiBAaZkhpg2MWvja6iT3lRu55le+sRRTLPCnw+ia3B7AmgN6Qc6X4sAuoNWY
iZ7ySLVSlmA5dVajXXthxOQY+tXJaxDy9ugaPiENjejluUOjRgbenPjWCzDzVPSz7ai1MC9GGo/1
cT5oX+kss/uMwBQ3DQXZ5kKq23b827JKfZNWJ3z3W1yUKdkoGy8Xtr9OYYy7fdxdBKzpYqAtvy6K
Hl80NWYa6KYTV1fmNL3YJwvyW92x+c2ujV9xaBpIsRawIwNWOa+YvlFaz4WYnd3MnKposj3tDmXW
PuvXIvZ6j4A0E/YxKoFY9t6hPdJ5r4yFfc/MMVyidnqpz4W9GZSiBP0Ng7VOGBaq0P5VvR64tUzM
KxSpioLXvpgHkrXk7XUXyvEeloKTwIG7S6OMG41vgR9IzoBdB6u5fIDDr2UrOmkbY6dVRe6flDH9
AVuAQuWHteqdwKMYJoaMk0hYqS1hApdkqxEbGbsZWv9Vfn1+VMV/WhZb4vMOH4F2VmuuRsikGNNH
0XPitFGdExafqLI2gOnj0jC3qq90cyWYgIn2rKSnGV3766Z97fU5vAMr7TdPu5hxTlkzpvK0ZbFE
Cx2ay5Tpt3t5755NirXvzdvuR1/Hr12oqWKPXZhyoimjWBjQu9MRhd0kaG9WJ2n49gm3C3iTOqQ0
HdpRGLkmO68Lsp4ClROHoNPeZ0cryJ3jVM5qB0dvskZ2YGxjs6RkuZx7J2/Vf6KMuXY1+Gu925tp
h3JVtIV90cvm4Xrg/6/4st6JIqfyCVQjRiyJgwVvENZfUvdEuLgeoXCeTz8t2j8BVPmPnb0BT77k
tW3q/bEt2MrBBVhU8qGFk7s35PHDixoy0SQOs2y5YbCVgucQbmPvQpTZP860m26gSDXqRKAvemEg
Z60qD3tKmPjNaGYwYLVSJ2e1KCqrWeDLZJMrz7ZoPxXPbVrHYLjjIIllWOis8Tx8YU1YvDscgkcU
rUwUrZYrgM9OjhhEgPSNrlHBanT64qxD7mfYgkPiBRbCzEpDWLlpnJBfAI0FtLFP3jVpf1PE/JEP
hIxqOx/yBjMQRhwQ9FJFMRY3E18jR8WAtoQM5Hc5m4SToet45cRhpjMWkxntmcAIq6YeJ20dTyaY
ssbFuefOunFLfDnleCEXchZgxj1aLqvLjTR2N7a5c/cYoRbSgqx6IAPJK/fVpnWqtqA0VqO2Pd4f
3B5JPOu8LcabnLwbmeeSF1aLIQkORwn2VuMrO2vKDi1fz0iz7bcPdnQRMZtRk5IJvgauJqZaMnnF
ODfun4l5R6ndTf2BBbWKbpk4hgn01VlM1BFU2e4WJg6oaLFJDOz/G1Kwld3jZ5JZEaMRF2w6mDhT
unPWSFzdNt4hlio/0xlKOruH6C0657SAnv3kpYQxNlYBGeSTtSzteqKkGHmm6S3jE/yZ3EGdre+i
rxjcvDRP3aZQhLPFMFfe8TGwj1HULBkBGnd59g0gtTW8cOQLixb5uzbJM166HqaT3xwQG9l40rtO
2rAQCBVq+vzPHeJLC1urbEJWeF2lQetQcwl6NAwJwvw90+A9M5iytdpLjtvsU8Hq/7EqFY21i4Fo
SAVhynbuaXmkUSw5/h5jZzR1kYo1SpElfnfZGNEEYAtXv/vAw1z9AjIkxC3yBUlmXloJgkDDdUck
WZweZNN+rfu7LjgAB2uhtS2HWDKpg04XpJ4nysuPb0GJ9nW9l41+Ivf5ma6S66loWRxNb3JlT7zB
ooWIrZCb3qJKYZRxAnvCruPp0ICewix6rSkA75ue6axfqiGQguKi1WN2AkJpKtYC/L6cYrrkZ9Bz
fqypdVWvQbM433O5N0OZg2j1uuiJwNk3zOU+wqyomJsIviusVXF14FkME1wmv6/BCflCZMWHo5Z+
LqZSZZI7LoTddJgy0mqRND7LmLA7wf5hv/7Zo/P0L78pTGOSwpVlDe4fny14Q7Ac0vs1iCZ5tohN
DhHRIgc1OG0ZSmk7ZYDoCZfpGTXxchnxw28BvmLwkCLED6+oWc7Uhagagv7iWqktVNC9D8BAeE7F
qIfq8gYQxt1Rx28f6jnppiUIMZbevudB0Dvv4N4f60J8T+LQFtSZtskT7RtPmhWTZe82D0SnKRhN
pC+AY747STy7dKFPVjqcCPUrXrFBzOvNb1PVvPIcD0hneLD3Q/aDCSDVQM6ZEv5G2Ju6F0SDxVsn
ire3VhSJz+eTS7t0oTgeecrqCu6tsC2p2nNd0/YD2s22M729baTwlPCHttNYzo0bb1A97AFYaPKQ
pmyl8NTxLOwLRhnIL21Z8RN/bbkQVGHq0BnLdgetbF33jKVNvyC3ntcg9pVWMK2aA+QrxQd+Roko
+iKAid3oJ9zMwo2Cg6SIGSULQdkjnKJFylaMMGY5pjUeLlKVsuWwznriV3oSO6ZO93GigRGlKUqM
p0J18AnljtyORNchf9iL+yN5wB5HXogIqSl0Fn0ssCjTyfSMdrcCmrQ2xdywXeLIvUPl+7vkogh8
UWais1StqjtD7SKzlGpLvd5L5F/jqiWhU8Q+Z6ERTp5IUASbLhdP4srjKbsI9Weaj3x4aX6gws7R
UZYdYI1+1t6mhdF2X9GWistXGAKYTDR9M/MLMBsTLBhwfzPD0siKZQboipKzkINkPAQISuqGlH1+
H8a7ovKRK8jYbAdwQI2p4bN/TJa2qdFDRcjXpcwimw2NVWUHw9C8/WfOqf7gBiQzY/9TDta9t69P
rNbrEFTrBLPmaEMTYtbffJ7KRAOIzzAGwSWGlL2WZRVrzzF+1KZvkSOSHay8NeApeQlhD+wJAWKp
DkFp57WJ9EnZmin6qNozPZyiOwaIj5F5yZlVLnhDJpy4VzQ55Xs6GDe9QxgrxxawqtMgOSTuR+5d
WSn/TrN8rqo6kNuxvztKeHSARetQBiLJrIP6ONoiMtZ/ojW0YPPvQlKsCoYFX+4Tu/taJ8X7oXEn
KnDKpfLMh6oPY0IDZvCCvjk4aarYBmLCbFPIJarToYW2SwmZgEDYsK+XoRjeyRl20SByq+d/XzTC
872c1M+Or8mq8iVtestx8ObZinA2+YPalb43pLcjkOS6tsdnASeBmkq/c2m8OXFgYxjnVyvtm4Bx
feErhLrqeCO19qEVo4I7k4eXvZkwahLCha6fGRn8fEKxjBpNWpXwLaBFcNkepS6lrp/rl4pqCR4B
q284pIRX4vHyqo2Jri95UUk4NPZ1Z5adkzvN3tPYrdapzBF0iM1yeQZE2BvIhtEWdOdkekhXQD58
vzAEUwCosmdRgquoU1LH4aOVARwIBHaGZ/K5Vgr/KLkrSzAb5B7HIcVM0rruGt6ZRzM6WSQZaCBw
zMAj78Jc8gPYXntC7mqhOoRo+6SLApzParFv6SorO9oKA0462R3vjOl+r7b63cJV1QM9CR06y060
o/EpX/WMdOgi/s2qReQIP6L/AypuINMz2JE/ndS4dzEACZUg4H5jKcABXIkNuqLJxjJtbGrzthso
hwZRFCYSOBDBlEDChejTMXkecnQhAJ6kqVPiaH793SsmFa1rj/4nq3nfvADFc6G3tVvUmxscqq48
glfA5zbtPBZhfWhWEP6C/6J1SvIeijVV3NmEX+PapmvDWs21lPP+b0OriAAe3EPm/xOBrPdTcwju
QHNV1s9sczdq1C1vwZfFYlVfhEYSUZfkxoPVwC79VA9T+Dt5P5CXyRoF7TOzqY2AUMaKPYMRwIan
NM07+16qSnsPbGb+1QDC3H6xK4YXwpaQlQl2W8g6IwKWWjOCgkYzecieYJ9f4HsulqUho+8d0PB8
55VAevj/OXwPyJCuskqgHJ8wUMtYdHLvzr6Y1B6uKyGCF5azs39BNHGOSc/o4cjn5iLAKxM+s0jq
4pu298ZjopPyh3EbJPhDYFLAHDZCxKof5fBkU4N9cHWBFC6vthP1XqM9SLVKasEOKKpBKFhelpNy
WZzA5YtAw9XCRWsY6scd0xvNGl/7n38SxOegTgfNvjxBS/rykBCPheUJvk07W6/vVrZNYwB3eoT6
Zfr8R3AmQ/ASDreHnmFhs002bTl/i4o2sQGsCYvzmjxx8BiXaicQUXSai/anHtOtO2TJFN6eJ6I6
vMh0OsqBdXUZwOSfD5ZfateVf/TuY83a4VauDt6AkqFMhwPPVyamrnW0pe9UgrwD85gRGaFpvzKZ
SOA4+DDWnb+BGhQc28f6IDXh00iSgn5/paGfU9mRUwKt1RQ8vP/knIYS5Zr1NOxQNN8VD8gUzZIP
S2UtbxqiQU66gGoB5Z8ZLl3hG1avCo1UNnIiugdL150sOkvP3U1uKWH9aB7Wi5MNu7k6ifeP85VB
Bj+YB9gvyiFG9w/RdK7/m4W6mcDlDara0HwDEVw9rymni0QMaPTHh2/um7nyZioPFr37xCpPlcQr
U0ghSsq9CsXcR9G8xeS1X2ZZtTowGfiUJC7aPoq7sDAJQhxio2x4lb6BTRx97ciI9Ps8y8gM9f7A
AnOryS7OBnaWkqS2vFyDs2noBbmCZZFfNDRdl2jGGMlGM7qJXI9XHW46z9EUWVIR29dEYQZHHzuw
Lr0XJ9yUTNb9vFua48jP01uzxFooy6G3i+aI1ZUaUdmWQ7+PXuM7USPl8a3xd/edq7o9Ekl+WOO3
2kMBItbOR+st+X6JyXWoHY3DOHDggg87vkGy4SIuoE2XACJrgUPof7kQupU94bFhjNBORxxBNTRL
FsXPFJj0s6/YcHIj73dS8pxaIAgM9veHOqLtFL5XU3HmKPlDF8UVOeRw6Vmd7YIVEXoJyU0mBPzp
cRh8l6K/U/fSFzDnofBr8TsQ/mVnisMtPzpb8rp1Baib2ULf5SXEuNFfbG2NmAC5/Tb3H+EaQXY9
CFgrPJY7MzgnSHY+Gn5g2NKW8MLd+G5A8qK7MxblaFFV6L9jU9d1zCr7OgYFKRaLjSJwdYip5v01
/SuQ0g1GcpXZa0Ynz/s+T6NMLAKS0ImSl5X1L4v/nJpWGPDFPMp9kDppQLpdUDfsJw1xcgdTPCDM
kR7fJCCCa994LUrzpXziMB8r9VGk2DT0hHgOCgltaL2hvEGcuRvIWbXFjGPq/Ur58XjAfMl79yQ6
IgSSzu62tMyL2AitEm9I8bKPi8t064slUpQcXWuNfv9/Th3+TpvKWM0LcM40p5GDjtp+1g9ZTXkk
c8d+3W7iSunAehOQjR8BjP6m0GxC8gOr13lfzV/5VykvZ7ISmarVYg0RP84WZ2sPmMYxjtwxxWze
sxtIvCmwSbVoWVgg/ho6TerNDXn9FuPGZA6HoaUtnGAZg8OYsLx7IyFMra3PNPJ5dt6o/P+NrjAX
pcwk+d7UaGefAoelqsWLOYXEuvrKtUXb4xKYL7yfL/AyufJ2APE60iPOH+wjmT7/hvviurAcnpoC
HmGeZ4hfPht6cH+O2rhj6iCqigAGlmv47VRtmF3G9+4uSys8vk/xOpkHuY1m/0H88HYaPO1aCtY1
zZtRywRrAaFZLdF+0AzfG6OiLFmiZSqWdbKGWUzMkUj/aAZaBF4gUNMRoqTI1JEr3ErWYeibEqet
hL/Fa+XCLmQAuU9b20BPPlLnMTWUxzTgzSww2wk5k0RYPw+iHKbnph0EICzkgz05zDPEFmhMbJPl
iIU5QnkO9kSszbdGMRZdaby4frF3CX5831MZkgYAypXIxppuG4OhiDayHCH2bIsSfg7ZMHsZQC0e
HehDEx/C/m7F8OZetf3FaeUrhFDY9R5cL775f62oK8ujPoqORb+EumdKJoOkb2OauuB4rQFC8X9K
ZzektvMi8uOiXtv0dpxemF4FjO9+F/Wt1QmXkq/4kwfDxfAZFFv8LmM1EGTCUKDH7lD3RW65UM46
AGjGRA9gnLXDFj2uAAlei+x6A/t47uWrDuXPxBQ7v/WdQPXICLV+8BcTrqy9nRARLcsjEHmsGr9B
bWdoMrpF82/6TSGrZCWAeDkyhBEjpWMXSCGnAJbqZluhv97QvdorovRC9ujMr4mX36MyLk2Gswza
/dbLCO23Ftzl/14x3fWW9D1uQZm9dEScOHsHg/pHar30RW2bHh5W4kvPRw0lyCnpTvvrP2thDhzS
/b/pv6HBDs8DdR4HWo4ZVTOfLNL5UP5do8qi6RwFzwNCxM8x6ZUwvGxk6UXYFWVQDKx1vbUhvYy/
jyqpWrexRg4pakQLENRUSbcaLjVYLrHWUm9yko92zNoA9NGznvqBmyOL5/D5Hr0qCZ3gaMh3eOU/
T/kuOZakglzJWA1yjWohwjapbdJfGszhoZffig9o31HwnzYRHAomVrGS6IhVOhlFK+4KYrOVCGaM
XU9vLGEUup2CMkzM2wYWtf/lAPOY9aVoMb2r+PHlKGbKRUVVyrWit14OfRSu2YHGY8PW5H2JYEmO
2xPoEaI1v14QyNYqVxS8vXzq37pDw2KQflRH/vbQAafWgIZzqufhc4BF23i8zMU7w/kzrMrJ8SMO
efz7OWKW2LfjFXlkKWulG87iOWNWjJzhG+Utc7Ynmc9PYEA0FF1ovmSRyqcO74A5SeXgkODWe+IX
Dr1apCw2vlZeicaoPMyl1oSip7OR0gozPOb3UnTsquhoBqtWAs8M85hFVbsJ8yml4t0B9qYFTuG7
2qLuCYOTYS4FfPOvU2SFJEKQkcD/vvRHbK6EkM6mWRx1arZfvDdFP6XNuVhcwccnUP2votOJtV26
yxr6rO61RiPBENx4hbEiA2zs3JvuK2sFr14FSUp0BwH2gqPyERZCaMBVYgaqLiZfWpV20RuVYch7
2ivId3WeNypXjUyxTBeW71MVAc9MRF3BNbV3FooXZZ7ulBktp1N4FnRoALpsfebGet19eqJQ5+vy
Op2HqqOz6lddmX0TKBXwYMRKFXA6DlEF8jGFbEcx8o0/gY0E2aMrTpTKonM5hBlJqL8Q6rHFApHj
O5P1uc3Hl0PaHEkPjPxtsiJulOLy3kk5yUtpOZP+7QLusuCzkHiBwD0+wVsYf1nui6SNCadeo8bK
RWQw7HlAMhU3jbD4VCKWR1Sn/Y4ExE91IlEKOyXbrlwU0BgYmoHTv64OCAMMXIBpWy+9fLilcvLC
kziO831EFUZ+92kc0zAeWfMNz1VU/YN2aJyIXkRaxrttp5VtwcoVe//6ogTcDr1DcIDO/DABdP6f
ndBPjdHFYBBZWkC4N+hp/JawId9z/DS380Hppp5jUidAaZHQt2hsEmTgnOqVTCUguvCSOxqOpfVN
bXp3JwFc4Mo1Kv0r9OKbY8nN5kqTL0EXDIr41QnRMc6HAXmXhkiVsVagowc1Z6zNtvPunlU7e6ez
D+3ljLnn+fZf2eqrRJhMW0HqoZA2Jej6D0y5VrIIjhO091+c5JuHmxSi+KfXy26SENwnKEuDqZ3U
OQPLb7qAnuyr2NNLQOQuhICdTDC18kpwSUd6Zj1p/oE+p3iGZ0zZqk5IQrnBT6TE8jTUMe3ca9Hr
Ecsyef4045fbl8VBgtzse3XMLuJl5CWHpco07kDunpefrd4Lv1VUxqtvaEgkMeuU7YErm0Oj81q5
yhM0bN3TrYhUSZKn5h+ynwalbum9/b1i30yj3+7cv9dnOgUYpyrpdXAuZpmx51ENSfp/u3j5+tdE
lAJr5XQkoCTKHGOecklsCbSXzDeDZd9jfE+KHzX1sVjNdsXDf4nQ/pi02r/IllJNa+QLZOVPixcI
g4JCpfEKc9BWM1pLWASGhjj7pJ6re6HMZn1NbHidIt+rUgP1dm0W006sCQzQKl55i6pbGNTIG88i
l1COx09UR2zU3+wps4/8WCqewLsffch+LIaMlPAyCMnKOxP2+uA2dr4WuOQMHyjmaiWvYDht9En6
i7yKPwywFAAD6Bm/Fx4ai69426pU7/F82zo2Yjvg7aMBymY1tVxT/FD5ORdbr7acuV7tBguzhxc+
lS7n18867C4lXB8bJACq3gSsqZkNtXhgmdgg1YJNRP4/Hx/GcCDZgZGHfMW3uLrrv3Hf/OPZaZJq
zOKx98pdT5REyLSVeNxUN5TVeRjTK3mckqH5JmwWOS5NNPDdi2u/SOwQ1rB4vLoUAMu/WkpSYjmV
Uaw/uDsiNSheJa0DbQg6hiijfBZi5m0xF2pCT+AsKSLW/KEt5PL8LMJZyXc/C58vkGP5tBnD5NgD
wkomKD2zTR0FKFPRA0dxmLcAbib5hdPYtrZrKfjEVV9gFSHI7inTeDlmdBnGTorj8KvFMVKEtbtd
KRvHXdr7NVAJ8sfShuZV9Fhz7KKHVtaUpLHWNUK739o5fuicQGZN0da3D3o3vfM1o+z+OHbROJy7
fU3sghFQxmMyFk0+phIKH7KVz4/X/kIGmC0XqrPmrLoS2IX3tto+mlzNSb9oo1/LVUGdeOx2gYZ0
841uZxo1hk4f2IZP99hr0tHY42FZVIA3I33iPyPpoXeY4gGSdr6mg5QsOaXalz7La4la1sbJaIZc
nj8QsAKRHp/yK7v4dyEA+MyKOCRDssbdNVI8HXsl/xS4tbEsFwiA8CMtAXgvU2yXlOMo9x8ZuPo0
O7JNyW2s8TO4skSEt9ow5idPE/sd+5D/5DvWDnde4yv78WNKLzwR+Q8gOTkVuaxA7Uyg6N6kJvjH
by/l8MXr9gvDegeksmIS0psv5J+5LGHugwYx9kyvRpL/RmyIY6vxpQyodqiSerlrZ+IlSawcvN7G
v08nAx4r3+rI/GSzltKAwfIhCwR+cBBBR043SG0FOM9t6eVkN+JnS1uvZb0vFUUrKGPW/ndmBbcy
wprN9bMzk/9I4Pst6S/TAIBXPuSAQ9yWTj7QMfEo0dZfZhMkiI3dHMR0fO3+un8ARciNrGhsTmBk
zeJwPB6Ih1k6a4lUzSqs+DWXaKst5uanYtnAU133DGp5ZW1ZkN5LbXLptgdllAhWeIpA+FaoNp76
R9PdIrMdvfwL/DdRs1X8UufZGiIgqRJ4CiK/I1+4jFBnLPO9PfCS1+m3fNfmx4GEsqIalbx6F4TN
L9hEJgg99W6bOQ+HVFpR4+LyLH/G+XBzAyKRoPudaGecMOrv5iTZ0H3YZ+vP+lJuKmUivJD6p2CP
Z+2R8CVR+9bJ7jdJB7tAanWfHQAImkcrKYfBSNa8HHHgyFSyatZDb2ZJYyurt6hL9ff9EqDfupUx
jWNtIy2qImxjreLRPgIkklOBCTNRg7VWAv17ZmVz4r5rr/c0EKpvYtTpsizlsgG4C7VvmMQvf3sc
Zy2vngY4RceS45syL8nB0o0rSENvWG7LdjVk/bhg3Y2ty4JGpxQ2VPxpRU/2pan//gHqviMskouo
MwXsnpo+SLwsKH9xA9DTpLf6vOIgDDmDwcjSODGD+2UyljhRDK46IwvFTMXZeoZCVvJiHORk+7bg
Uwv1UTLwwCUq2b5S976NkgcbNkEQCt9RVpp2KFYwyeoIf8UYmlc8LiKdP90/Kh364WHTRacEph1N
OEYkyGlRlIkEmcNi4kRs+2FNEMvTvjRGgRWgteNPVrg8ASJQOMw6+S2swq31mayVJ/LsDh81PLNf
Sqo28iw30K4+NjlM2QUZZTshRZfvrpe+1PzCVHyainnPB7ZcsxLhG0cym97v/QhyBna+1LWcwgDb
J0T1nGsha99sQvbvi9yjqX4vHPitilXZrQRUZ8TueZ0+3PWmfyxcEfqLZWXMBO+yc0UwVTtFNgOp
BLcXimvMzL6QiDjtDMAgiRoTSo9kScfeLaIjfCDoRf3ivd1QX4auEZfCB9OezrqyWb4FOOj6mn/l
oFarZEQrhs4mwV8jj75ptsSCNKI5v1uuO4fTZB+1egTc2+5HnveyL4aboe/wK1+lD0mBmitLSu92
oh/u4OrrPFfQNVD/LGD5t3l0KwFDrauPv3GYmXzW0qClfdyDp3P67tgZ6xrwFx7n4cjPhedQmPfQ
HEbJO9awWg6SRtdWEf8QcyyxJvqca06tT2U3z4VrRiQHxSWRs7oZdAdWLrWlw6/ijsCDMkmnEtqy
QpDEz5DZ6SzkkDEBZG7OaJPNkrE78TmqrpfMqwyC/aaj2aXbgGLNmVj5jv/IL2rsbIX6M745U9sM
U2oOcQDAXLA6yJH0aScOlsMsMe9gLWJoMLxRoVdRT+zqz14DT8mvHw5a7UhSaA9KL3A0jl2pioEh
8Ca66J9TKa7TB00o/vSnSYcpbZfmUnnL2lhXMYqoM0OaPK5meRhlEcQTfExZVJD+pRaMAEYSXfWU
UqTMij1AzvTHoGzPeHlYHBYZdSqLhLRtQIbGMR1pQg7rsULmI2G7UhupQXwMblJBmS9sdUExC7nv
PGF4E0jmsTcP8nP1dMfrgnO8dxG9vG71i7ptW4MNXOg7aqvdGJf1I2Vj6ppFOUsKZcFMg5kCw/MX
SLvN9Za1aGcS8NHM6VZdHHggYq88trqxV9Rc8ClR5oX4tc5QmfXBPSEiq8ppZLHvitC4/yUF2Nls
vbqMf8xl1hT+HqrfxcWPOc+CsaujnbZEhEqYXWlk9YYpsZdpS48ydCnrCXIO3ViirP9OU8WMI7/R
BtZHypUMMa4eJGOctMpE80NX4DCH2XBHniIpcuSEyxkeCruZnM0ktrA7MQMmwkrJJM5luI0OfN/V
7ctsb75JXRfCrwARwfHt1qxJJxW0MW2evTig/n4RHcV2G7g7uLl7RoIx4rgtue7y+61GAYrXrxql
JEV/p7ul4zWGBLxUCKjko2p32ixRfo7nE4vfObfAUlcke+r/oZGPC6IXqBnV2woKiad7xy/mYaip
xDenFoq+rupqoU2zQZwX2yRozw04ew3S2x2vnn1tsF8iy/uJdd11czSqJlRGsFpym+0q/nLs7PNU
h+ve/FM2Vyy1dAwB3u8f/BymMQkQWlF5DDAzCpFL+zGNzY3Hj8Jg5EQ9icLc26pfNRa+gkvQ7NfI
dwqr6LZZok3yJd0sD5xBUXb1QrJFt6rQSr/Pke3gkQVK3BHZhjqBnxzJOMYf0AuIiIeJ+sz4x+iN
FPQABjpMqdXe8IQJWxWIkQBy4vnumfF96p0cOjYloTybbJ/2BDvlBbLtbNtXIsnH2VIVRHr096mL
jTq8AXCcYRJJhbQyBNA2pSiqsPOMnxS2P7ynCvP9vgxdv48Q2PJQ5LX1Rq4t0nollYBlCZhboce0
THS4oiKv3gisXrHRCkZ8hKkbAL8fkE8CTizIq+H+A3nxvpQs/IJIYc7PAMsLe/k6eZQFpDzs/0+Y
Lj0M4PrvZ58RNO8DgFRN1ICot3XvlIJgJiEnkswcfe8+mUGpTvpcKswIZ8KNWBrmhWVZ2IHmCqrN
q5l2bDsOI8L50xD0O6NjtjS7yahgPjc4S9bV7VhKZH0cioZEXBS+75rNp489lLdayKNXFN68BUix
HScRdHj8LiDsg0bkhoHX6mQO01UEI3yQAKizSjYCu5cPpSUCOxXexQQTNC3LeRGHwSAb7V8j9e1m
PuNIM2vqV6RDYDWFygW9G6SIP64mY/YoOdvNqSJr/xMNgWh/K5kYFBgXn7GIWAxM9BOG02pji/8y
6YoREHmVv+yKcMSmakG0T//LAI95qtqJCz+rL57c3nKwiosMYykksPGQ33cBG29l+BMt3vdBxI9s
Xfmd9MluhZ7womS9213RSwn1Nyc+ccgwVdwRuz4Qqs/iGeZ1+sAdyJAIv7RRXdAzsqXf2KNcCHd/
inDkQ/tvbBI8MbyLXfUE+TmUMXo+Ie10xMLGFHGYeyka4F3GLl7/DSPr/AaAUYr3kRnl5SUMJbas
IILqOKVr2W4q5UVEtx2ctL+SksjssxYIkt25k5qEbf5lzHEEF/ZVdlWZYaFOWJ8fM9lzmwKR0feV
MBgqfyBtFH7hRb88FE6q3fKvO5hT9PMV2juL4MzJKyX2N4Kbvmd0F7PGvB6lhX6H+FeeC5ttmf7Q
7t2BPVGuxWMt/URNz1GS86NHccUR0J6+ChzypR4RFMZYewVon0P5vcgjb8aNNL8klHmaiygZKn5V
ZxiTnB3GSs3XAtL9P7yx44RwBkDK/ftspKjOmW93V+8Y9wVanVNdwN5guJbxzsKjvFiiHXFBoPqL
BZ8zpizwoaI6r9TixEs/mezNmh2d1xVkJ/wgM5Hq+xG5LhkEk3yUghfN6D2TYEqkHFhsBWcpnUeI
M7UwNRvhidMH6bPw741OUrUJioXjPPRVHdHucE2Lj2ch42YQ2jeYCSPpeFUBTYMtGTGCM+YYDBsC
aZv/l4+jbDA9dnWQYXVkkUUUfd1sLmlXr0AcFIMx820Xv3rNo9Qnnl8/FBEydhziDxpXnk0cY3Ou
iuTX9vqMYvD+12owfVhYJCog3WQ3gswhYLfElYmE5XqLFl7234TZbmFYC6Mc6Iusd7a01RST0+Iw
fM0Zj6Fw9rbO4rVPr8qVrEXQ2s2YHyP7F8WR0oZXiWG9ZlEPKfnfBV+k2jflj6c1lLlmovJWgCXR
/bYRh9h8EhjN81apbZjPAAsENxcokJKMUs0o6imJ2uJiNmJ/c8bb9RxGzLgiajZDb0oWPefyuB7P
A+N50wkacuAWDWGjSSuNh8e3CQsbUgnl8Ls/4M879/fKYKixDoL1l9v50mreo7kDPFgTMjUZgS3Q
sZYzIN6/3IO459u8b0wTR3S5xnthdJkcK2aXVmR+Cc4BMLQ8nrdlkiyMENzlG973NdDrkauojLul
3AB4sfngz6PCK0/YjwNsz38kWduGlYcF5pP9LtMQsmWB4VjoPcVlnqEcP6kzWasTBldeVh5CzzkT
L9l+Gn2wUX7EZiRcOWSSq4wUq5UM7ZcL2jy1R4J2HjidMsYIcKOf4vypJ9W5RZnBpZl+tQgAImRY
THCACCpeGGEPsLTXeqt61TD6eCk2LG9llNviMaVfIFLTeOXSgVu3YZ3FZnEGdajYnDntKYTW2qI5
E9PEJ+gcg/ueTvU0cPh+BYUgEHMeH1FTd45hHt+OT71uA7bkqJh8vycTIdVpDjdnCL7tVP8dZ0Ki
KXJMiYAF54T5AibveZ28L90mTpzeKQ5mzod+mKYSCgfBNOwgeWWyIqHxo0toNok0zmKloXUQvey8
rPyDgsDWcjQgLxb7NFnXYwkLwOkH+nQUvoygQNrSzfTaumOVD/gR6w9qV5uRAl7KMbiqz9Xf60hO
dwG7oUjIu0noC8TeVDG5OnF5HhWAv8OxEZlIh93MxtB1MHG3lFaF5gBXHiZLGtXfVSelA28NVn/P
8uJw7+Nkme9rAEf9U3CtQvoRbfQ1FfuldP9O2MMywo4Xpw+qCBl+1E77wZhenXRC6K++sijyVOjE
UGjQCN8IBQpr4P+TMXJ1xQVl1Q8GxeDZ/oy9lhDYfkBS/jjmg5xMvitPVk5tgDU3ai3AUG1OBFxV
p+BXc1notApNVukD7LEMy3bYXo8YAiYnwgGdvsPP3EAZsQYGi65aEN65KhkyXaLz6REVQMdNqw8q
RiAZ9ZtzQAevjkDHC/J7IOlq9VN4CkYz6NRy4i7h/CNI7p/EPZrniE/Tlgq15ImhX9pGvRk1ydgP
pxQerPQfpzulAc5Ura6nwvoEktEa5M3wjgHeqazrY8YFXKc3i0q8WBGd18PhOCI24knh/MK4YVFL
49ZsllzV7vG28sMB2VPXu5CoPF4cWVMZhgTJ55e36Ff/UUkvcYvh814WMZ3JhJRSvbNrWKy2iMGX
7M3RJr73sycVEuTIEVGbei9BYUUfyKwrk1Up9gXLxtXnRV3P0VlJhRO29zuHJ4Vvoif1e8We5amY
Z0jmyVHq4dtA0dSt86PTlJzIF5I3ts1ef72CR6oWceZVmT+uzv9Ec0CbeOZoEyX662Ws1caqFo9c
++8vJFc/u1lOeJ9GGhkNsfdOHLYXN8jH32e4p+zPGMU9z8cwFa2MX0iTh8lQyQFwqKCNE+ku5J4x
jmgas/lWIPTFbFm9HL6ULtnSjZWH8lzMs/z0z28iNQ+MqWrjSEpXEn3XxIQ16t37aj7Pi1GPCxiD
ci9lNcgq+szH8iqJT93vQzovlS3D1E0TL8kA4Mbm2EK0FYO7VAUyeLblKWutR9xxLxvH6I/eSNDl
ymJAPNcQ/0Qu3vcMmgAb1U5JoaX5/jelL/9EsvscVRlwD4TFcX9WCWa2avx3bOuwOZ7VsEIMSkeI
EQZEMO02nglIinOIQLGdP1f+xSkX04Dg96SUsudlU8XM6QGlbbrz2UIT5OLhlvexp/nyKJZ35Eg6
nunxa8s+sDmpDpHpSPyuZdr1xP++Ml89pcCU4wtcIL8gDId6HsiXRoZB5KDHy3HMd/uMDau/EhNT
mfOUF6mWpb+md7Peqxwl2+z1Pj59Mocg43/OBOn4KYYqzRGvPel4WOu6RCRdhWrArUoGa99sRL5e
plxH2yKreSM/pWCj9eE7Q8jPT3yrrnC8HJc+qeqS7Ngebi12xYP3EfU2CWVI8KtWrS1ICzN8IJgb
GpGv302l2iQCCu+7a2ejpY+VT8UGYfREs1QaLSok0UXALqurmSoUr1al21YiES7QnYCiIz8E4vWm
zuGS2Swj4np5wlCcUSN0l1TFdcjlwyLEBOeMRRoC+l+Aftet9+zmx7jdKJZxNM2s7HojrWfN8pll
1vaHlH6KyNeMXLskrl/V6v/xtxIZGKIREPKVdACy2hiZGqt8Uv3JZhGby8fgidCmFqKDdFD/bmm7
cW68haGnfy6BjVB9kbDXy7Z8yJimdRDmvVJnWGK5cX+7QEjQG2UJC5JJOEShKGVmDVgcGUwgg0sp
piTjDiB/2SP1HnGCqWQxSxjxudqAzyl0q55l13HEQE6asxPTx+ziJh6EtSoF8pRoywmYsucAHD6b
LkfW1jVtFR78H7yyMlU5oZm66gKe9Ow6W2XntWqvw/U5cjnLeaTvxVIaVjPulY64fHerqfiwXHrO
iay48jjykISzVuPjOhoeMYni+pLrfQKLfzo9SQF2/tmE7M35NoDnQSQCToJD1XDml/yP7a7vYFU6
8ajcC9YTZOzcwjOxniYLe2egmuhXGklFIYdAswF0TyaoGKQLOe62UHzwLCbCgUzYjA96ZC+tcHec
E8UasZ2oA1Y1+iKhuBsohJrCWBt69jQAB43P13xM4hNbu6qtjQBz73hAd0zAkwE9BSPx4EfFckOF
KFhZUVgOBMwuNx+wsLjrVtW04gfPCZ1caS28ZuP+S97ibWrXK7fGea+EciNjUaetgTpu4sfI+tUm
qlpkS7VR1bCo7M+N5pe8CJwJhTHNhRSFPtm6bCtoga7rR6AB9FiABh46EEcYWzkmXdCQZrhZuYne
Dc1BWvCsZhLyR0MDOyMirLiOCjolRN9zTKPypsib3jF41jSCwPu2qfW4iE23WsslGOMacl8X72BP
QwNCEaxuj4JFcQFvzwqvOgWJh/VQdoIbKkU9GKLY/N/xrxlKI+NPLBukNVNyGFj23SNDpqbA3dVz
bYb5zHp2+gwpsMAHEhAv5OdLXuLsR/Ik5ems+qAkWnif/Ad1QomR8liF+sRMJqVU/ry+vseGHcFg
uVzFHqLJDQP/zi6nsrIQkgBlrGxiu0oc4VPRMMBKi/XtXiVrOp70fYwgyVrySXKKpFiz5VPkkFtF
NqjmYEoNcTwqGKl38AB7fU4P9s69x5tRfitwa+vC6TnqbGokIboHcmiXNgVP5XwGIiIZYL5VcNqw
3451RI0dQG+ENcN5NeZhfeiA6zTm6Tj0KUY5gsLFeBx6Y1OzYhNpzgpRdeyPu9/L7a10ChDkFFI4
DpqwmiPecAteCif+/C43aDNdWwrwvxomCELpME7/o5h8lpZYFUFTd913MEQrKzmRLTPIjinsc2i9
qn5DWu2Da9R8s2k9t018sdnICmdWIiX7C87nqb/36Y/QO0NThmadMc9CvPkrpt69WhUymXZ2FPYA
UBjllu2XRpviLeBjnKU79Kq9MZyFlQkmE2YnGbGufKFmbXNqL8FXpwB+4WU9JL9s3UFz7d+B20BZ
/AtF76LUfSTMpllJtFTfG9P+B1XKto3ZepZqrMtqpf62jyKarpCoolLpzP5rM3XDoyf6EehcJ4OD
+rohIjTBkWrmnZ+gPBYw/lJHZXtFkpgpkPJs+wC2f1V2SbEtKblR/ED2MGF0oMsqKgZZ92tmpYM5
SgARfHsu24pg61AKk+lSRBz87B4nnGH1QNQmC2g2PZZDD7BSK6IQ/lgc+HaDlb/abTegx/Z5RS6c
BcvgjiGleDnSDYjndPsnwuiB+lydttHjuMCrq2aVymWvrt5yrdOgBj9+bTUZO2GhdZxKkv6LXMF/
6S82MEmXmKb6RuSMQRPgqBHpkc/Gw01TbePGdDK6/A5FYyWAMDqeyIgeTj6Ft/Cf4qnkAGJO7eXd
R2/sDl8YvSvQguM/5+L4ECHKb8WzKQC9wwtsOHRZSba7kjJJErOF2bvrCImLmJeAv05BEI38X2LB
6l+NV+RJ8Rqn4b6MtnbJdEbmLLIpOaVBVL3SdbhLQqq7XAj4cWaBVCW5al2ICpjsRvrLrTujxQ4K
3bYClcdXyHM8nrWWj6Ezd7g7Yb/jQ/IcO+jNp23J74EvouNPbSUZAMH7Y4frSKFIVyeB1n5C4qFR
BYaeV9ArU9nYFQXpHj5A/lkgk5D24TMTebxNz/QBSkcNwiUp2hJ83BNOdT7yT5A3L5HErf3Qx8Az
Zr66v+KBa79XgczFhx9NsxdO6H+xG745q9e+ZBrRuP3TFMJVhDZwkB9R+XBFp5ACOU/99k2CnyYb
hCp2MghOJl9SX2Uua6MXvDJcwMSwKbSPD1I5Ch2IaLugMapg3dGMIZIkvRIiVsd7ObLBKBRya4Od
EIqNyugm00Sbhprd/Dv0A9caiNfCU1bIZaoatdRHDK32wN74PrcBtfEPlYWhTWTmvI3NlW8zRi6C
ZO+gdTWHt1H+KDhz2ojsjTgynakY9z6QtUosQkLoKIhuSRr+zQDwdtwLfEB20xol44xzRxJ7JjGy
glwZqF0AXG3GuWTbvrHHMB1GBwfeUZ0ntkiGG52SVcp1uc4i28a/rLCkM/5A4KRrrNIfnXML6B99
iDHChrc035fo6n47Jt1tDipsBF/WPUnocLu/1rwX9XSj9te3+LvZ02IddGcifTN5dHRHajcGzDi2
4uKyb9C+u+DfMbgQ5G9M5hyVDf0vAauKqqmZcAcJ7vmp8d2ljD8fpLrro4jTbPKh5eTHzFnWC4r5
ZEpGFURtGyoE2G+M5dvt/p0Wfse8NAbOp3+jgZAZ0FC2aaUG+4HBVNa28/8X79GFW/Ii7cDwnhVU
s38kRv++WeHAFqb8OcSg1z2l14/XlqlyckCOMw4c+ocN49EelsJuv9TKq5nRouTNYtlJkY49FUR5
ovpmRM22ScRXH5gbzOBjTn3jISrRq2xakh8ibVHMsHEDyLGknphJe2+9qAnE+zBgdBqzomiOWoex
0k0V5VefCrj0le3NQjl6G+4oLtLBfSexJcAZKFl3vyaNX0+uuYjNnePseHyldg0yJ+j0CjPGiEFY
qt4Azq4/W5qZCU4jjgFzN1ldd2zY0+RKMYCOE+9XWIL7Rrm95an/F8T2cePKt3z9WcAlM1j78xzL
OOWSqyjZ20spMNKVKnN6E8w5ZXx3uUzkpF7qfUzC0L/ztRt54Rm1IMfV62GtqWtv3jiE00Uu28hy
ulDACTe3jPLGwxx/0TBQ3P21QZ6aX/9YNjtBt87Ac+RktoOxzuXkL/O7IxwLn7BPX8rGAkxSg8dk
g9gBla81KHjumHhrr3YdjBFZqKW4IT7uyA1cW1MnrtLMYKjLarzeDM3kcu/94E5u8ooPfOdgNKgL
xV1BF+42+PvXmjAlBvLD+pnePOcIuFFlAd2nUvEcBfMMxLl4Uga/ckpYRYjQcVdymi5LuMfqvjz7
og/jX025qwnrbg3GRURn43Hp4B8RZrY0fFUdJR++5z0k9mbAEGdMG3uqX+jkeKUm7KMXj7WB/L+D
EQxsvZWPMZP8veOP849f+6oum2Hc2ZIhCLiLAZczMzO46iCi+/0ooSSbT1P/vnt4708WsCR/9L7T
ot2ny4vJ/J+D7K5s4vbWAuVsVrtB3V3+sQZh1pLTKeJ66vUhfeSVoC65Dhc9rQAqOUE+3UwBPgE9
CmovFam0F4UAG2VDATabByBJW1AouN2XHTthk46yEd7RaahLrJgTcOGfSUGXO5haxQldRalqScIo
c0OPaZ/iuHgRoi0iPYcJHnoY6hWvUmlHE0OoXrjMXaF+aL/eaCny38mVZO++5+vpYjtW8TZ3SMJB
FdiWSuRY/qYdWnDtKatvgIhaGUm7JmU8UgEVCwlGt7CsVjqHSz2AqhS9Y/8t+fPFZ5+05yLVgBBX
ofLsHDb28qKzrImYxx4zmzTB0LL5qfKce0Ai4yVT4sYsM9BmCAG6rg8x7F/bV+CqpVUqa9P9kb5p
RjbZ52bLKESZjsMcY5KXUQoNVehAtBP0kjc3Y7E7G1NPqJ16ddsF3toEnrjb+YSQDFLm7oT7EQkq
QIH0LKv7Pq5vsHcsqkmADCEBlVC+jKhJsGkxvfteqo46hQFXzu0H033Az6Do4tw+gmdnUHO50P/a
0szo2n26BrAOFIefQDVz9OrxwdkGiJUxNg6X3gyASeX2OXbTJDv16UfCbMtNsPnnECnyZWN39b5h
WTlrhJTG1zLWqrjp8IMWAkh8PO915h1VztShm7MgGB5dIQwGSz9z3XxPYWmDrOwlgkaizpIaHPGZ
YZxozQKM8g9qRqsLYwVuzNeZiHS2sct5agp5htTPnJppi82qH5CwBAcDAITrfbEs1nEBAzFflvxF
9XjD/P6RFjUwRuj7fQV+Z6VnAlOaW4Eo8bDV9//XRLGaR9DvlltzUc0x9Ma5kITYAOD9pW0kdXaN
oQrB4aZIMCnsfT/WBrt6/MXKr89d69sIjvjxHVWCuuyOicr4NQnHY5Vuj6E44dOJX8seh2BlQb6o
Z2SRyzJb/PsqT924LROYNAVVIJyB0WxknTcg5pWN7WGnDfOzWryfsVze1peV/ntox3ZlmnP82ztL
39cagQ/F2wk1VPVaWTHvtG303BT2ExsRitPFmucuK3fAxwTBC/dfO75q5UcGYgUfzJ+W33JzUhq+
Yma10PgOFPLaLdVipZrJ8KQbMTOrIUE6zSxIYEOGXHx2mE30tQWjhDRhLk8QAqwhSAwfq358MZrk
SIhm5pcxqGpJxEgMV4wxotEPKT2AWnix/R/deZj7i6VM/bhlq1kLIQpGJrWbT91vF2vab7U73T5K
Vb502tPUg6MhPzg+A9JdGfjQxD4JPgQ3v/3ioZVonFg+FM2K5MoBoYLAKjHp49ctZ84pkORM+WiN
U83xt+lz1+bJV5QrFN/POtuBw5n0unuG+QYbVsrLwAIy8K4OCe31+yMnaW4eLD3IblNy1L735N77
mWKb3Hm1+OxnVQB5xRBKmCvXAEE14SIMtuNVQfTMzgw5CGdO/gPQKAZFTQeZq6pgQrMNzUE3WvcN
5w6Fw/lA1e4MEV8L9XFu5Zp2J5skR1uoe184UD3EsIAS1iSvIxnqMfoo1Ap4D3jBV4PX5GuAf2U/
usTrAwq0RkD9ukDrKcbzTc+8O+1ny1yJQx4HJVNATKx8xb37cwH28D+2Jqbj2UkV04YinnexHKGs
9oMmcGZAu1BSja2G00vThrDAr4eatda6xkPV6d4ql5DlWr4cGVSTIA3S0A0V7chs5Wx9m7nWs3oz
HpB5gHtOyaYI/5a4ZN4LUHIPmN0uB6GtG0Zbw1wQ//1ky7UrrWRdqKhDtni1rasjbuMWN7psk8pu
j8v5JRE8vu6tOKDxZuip5lt1csI4HWpLW/mAbGiuXsookq21P6B5Ft8SBjteEz1UPG8gMULXLb0S
ScSRIpgAtLj+/tVKeCXmVqLU6Y5ciE2l8cnujDrGK3FSn2To2vypaFC0SxjYYz1InLwvjNM3HWBX
lAaC+dIMAGD4MMGfWfgR+amkbnpgs76uY8ptmsq4dPpev0drRpXpQ7YOqzkXPiL8CpIJN26xZGr6
/lfnbZ9LJ+nK596EjzoZK70tdcNLx20tFcFqnOKIkKZDDqxF9yVL9HnSgnKAF6Vn1vnzOQPQZGuR
b1XY+WNtxAlnISfiBqnFwFbe1W83FzDPP4QQ1EeLu9PI8Q2arAdax7C06lPLKdUU0zB4gQ1NvIxl
fMiWvFXUjm84Z35x/5JKdmx62+WHuUkXmKvk9MeFzL1WanbHzA48oMcCBAg8BfIzlnUS8s0AlEpS
I1kWfgsT7mTrZjZ1LK7X51altR9l5Q9LY36jsbmC0/PxrIkLJaHwwjqUtAXgUVPWThrJFe6q4na5
EV1vlS0S41dB9156V5O+Fy9nVUfeu+KJy1vJ558Y8KOJ9C9D722ZgQxtYgXOn3cNPAFQf1sYid/6
CWzjDJyCMgNj4423fijzfLufvi7G5EFIu9qPBh6hZZsQQExVJZPT02zu9jSK2/twwYVQWN2PF6KF
p3tpQodeGhpGPqG5UAlF1jBSBsbN72VDQNeLU3PxFXi8hn+zYG7w9BncrwGcN/ZQvtrK+gEUrgmz
yCrsSfO0YmLyGmJVaTJ6+T9u1Ab7KPH8FSj+0er0wT9HYumC4sxQcjEd0IoIg/SX6/0X/iz25/ne
txU5VSyHq2sedxQ3WYJCDildQK+lBQNT1sQnvz1iewf3rOwenl8bFc9iQUIqrOaC0pQutG3WpHHv
zV3EaqkZlxjKonSH++k6ds9noy32SwpYlsfZzsGGQNdJd/upwu0v4k1s12UXw+tRmi3+Ehs/a0OQ
3ej5hgA+PRUKHjRhQ4EYzsLijdwZJ0RpG7itpvV0jlJ9LKR5f984YEdqlsfEWYQ4AAJ7fGiNmrNL
fhANUYZo2LIW4i37hUeaod2Enxkcy3Wk7Rx5wKZHvNzwqRInT9pyh/fexGS4DEjovaWq51M/TeRl
jk9/9cAxPoRgwi9Q7XOQpEq0j1127FOA6esd6zfsFVC3RQTcKC7oqVaRffZgmAmXWBeDzXpYepIn
fDjmJ7mFzrRrlxuqVSNWF3K5oBORkHGzY6aa4FZfEMVvqS7bgrgQjt45Tk8wkQtL/lYHwBAmEpCc
as9mZ5NZkJ8MwvsJD6IXm0tRluPZc+XxPHRTcjZXzgcBzJuwQKu0gt+jLDkoCtilOiVQyPpoMZFc
Dnx+q88u91yhiVcGUCveWcFi3++P4gS39uHU6fYNBCkaF+7FlD44AkFTeYBdAFbNrzL5OBxP85kN
C0HOofU4ad6OljyHEJcqzlhb8/Rh5OpMfYvoWoaVMFuWbY3eLPCnDaIK97MGljKCk5GhZU3xr/oe
+ddf+TV1z4FEV3tAg8otmrYapyPIX/vLfr64diXrXbCye8QrtdArq49H7kUrCjp2yu7Bse8KrCt6
dIKX+1HCd+UdXvgOYF1IaR0RKF4LkILc056+tF57dUiTBx3lZ747Zk/0a17zri/n/GNkOf71nw1K
4+sruBe6cd/SVvPXCOIdNhSlSibEHQ4LS6u1m2mlqQOIr748uuxy2M6i+qxmXIv40pX+zWHjSO8Y
uTdZ52WXqK2ufFrWlUX2ytC3WC1kVA/o+Jv/iwRYv/nc1AXRS5B7jS54YdWZPsjZ3KoZYHiJ715o
P1zdsCQxFURPaaAIIOoCPFMo/Jdt+U09CYbJe+zpioAyOWJjFPvAIwfgeFByJQfNdX8/qoB43JeS
w5fYwK70yynTIm7FYUr2kX02JoEcu3QVrwihFqFWtBLjFw2JjrPPC4Ja+O3GlFkP6ZvfhyQSgFCM
cRGxXZ1MoH7R9/nPHXSgIZNL3LFRQ5JAva+J7A3AA6SvwUpuKABXHgDuCPPyFLWmI/QRHb/nK1tB
gACKoZ/EjDGrpvuLUhY/kPU0Fu39ElYP49i3Yvwmn+01IRvTuRV6B97royY4civrQ/H08DdOyeLH
eAo4rP4qaXllAOrFYOjJHGwwzAyNMohYyG1CE+AwwHZW8tvwysHQd0nhm+4hTq5MUhTxzUP13jAD
u2+N/B6G6bhB6yWvqpfo3yYed8pvunNwfpBlJHl2W7gjmClqpH9UEwu5uXdeAaBAseOtUVWzpZkJ
diavY5jGrjcvO8WVJc0asahS4Pe+h9VWpE6GREC6sMVFzJJX0p7+bTxaF74QxvWDHky115ucNdy3
AEP1bC6Hf7ve0E8ogQPvQ9MjVuIcH25oTSA4N2Zdp9gz5At9WTkEIsB0iiIwS2Dq7EDfUZMrN3Ny
NJ3w1zNKzEpXgL6IW6vLFJ1PZ55e8VA12Jl+Seb2njJ3JsaF3RUhRfqQgvsneBMApD18xTBbL26K
6TN5DtaUOSEucgkjHLOkETWAWF1qT5JWoLXLLJlJyArfQJdYf2eEg9ie7h4JFv2ZzV2UgzQ/Pmz4
TNWL18YGavYCg/x0P1gYq+Zeq6MHENBquxBISCgQ9YuIDWDD/hQj7Vo5uoBxZQ8Um9Rtfu8He4+7
SYfG5f4AS4sP/UXsbRnQO7sJ/4o+ghQsolaChgAFxmbG2vS9plYpHJC/Z97B7SnFFgWbNK79uhdH
5NM5q4/11kMKDJeDJa9uxIOFa034DNbc4Qhj6RjglDUcdBsKe5fI5GtJ1XaK+XZTKx9avQYdCt9M
149rh77KyECIaOGUgqe4+jcCMSu003hbBZG8XagTCHs5tfaRquj8Gn2HuPtDjydjWxSbhnxE7jsL
qOqb97bffALaBXJhBUFH0eeXO4i9Jgxzwzo+vXaBQjg89NbnaQHqCGzz7kGFzpDMMoBWNH5US2gT
g7tdxBw9TtxnCJiCSUzs2gOPwZRWnGpYSXIFAjmZxivP9PTPxKH5Ip2bKmlg9YNJ3+kwW0m+/rjS
L7RPLnMvzmtmPc5Wsd6zoSKxabigxBMqG4Vr77nIYK7XBsGEjzYJwggAW+KVZyoWIYfaPGlf+sOw
IncCdTmosnahs9Z6prHa0Vld8AEJSJtUNQM96JTg3sh2DcKfcy+U4J5U9KX1LuS9GTKJp986pKCe
vmPNe/vdLWYEGQdyxH6iB0qvlorVhLTVCuuq1pt4JpzQQfi4Q8iY+APDkLpb/5FJAQob/n+j2u7m
bRXUWqn64FfNzRhKF8v5mD0PWpN3OtKwptyaq8eTpamBGslf8Nd/lThIe1+ugjaHNUogtFsQ5Vfu
xnhIsVUhIPl51hUdRii4awfc8oY4ueuI5l4pMvGZ32tbFDvaV2DrUnhxk7URgPmV1uXh9y7uo8GB
41VJJX5A4DD9wTQfwR2URrkTX6xs7x/1EMYScmuDSBYhfyFl4Y/HRlPkTmKcx8yQhlttWQquj7/M
PKx8vZAS9SLCkzRdR/dCqPE0enwzAv5zYuReQRx+KxAsKHsC3Yx1Eh18bEo6hxaScEjRKpJyjg57
QurRp2Er98tbM8gKBGMqyTheFAKUNk6OUznrjBOejsG52l54PJTa3bmWLWIvVyeO/f7QXrrOTMQT
jqoG66N7UOmoNQfn3a+3LorHMckpELfYiOyU/VuDdh5Q/rDAdYp7OK4rZ72IWVTBsbThzLcAxAz8
nHZXcc0aNLyX+PQ2pwgAK+XWYlanAawswRZhxCD5JQJi136uo3+lzva8U01FJLoL8sZe9Nkq15oi
iy9of8U/4zEHpEiBU/kiYvDVMz9mVFLEcqowmG8bZCECgbAyg42w4MIGAkg7Wjl6sEfsJE0k+jzs
Phf9gSPEqNiJ+TUF9SdDDeLAzLZTL6zMa+ox3Ehd5b4XKNPffYxKF/hMxDh7rxFRbhLJlVdMzniQ
gT7qLXjVJvvy+8P9pqwqn8Duo3UumuPDClohkar1fLIbrnvkfuu5D9qaSmnGYqY/CGjALjboiRUq
yIyx3RF9Wr1uhk/8tWagqJab3EvXkLrLnseBkAUK1U4szxq6kvOaxxd6TjADrsRoHORMOonciBYp
yQBcIEcub2b9ijlRf391/K1tTt7Kt6OvtBILtRmkQ9sZKEvik81hj+71pIt6+dBWCrVTuW9j3Vyi
zglIZgOtiDzlwTxH1kzx87G/rOPd6XSedr/EE0xAutSE0sR2qd3Nbjg5GM5M7qXZ7opOkIHt06r0
nCtf9AlfOGBSSsYcQrM5CI/wqAlk0F5bNbsokFJF8wgTpN6/emHGky1PWl91IJ5v/no4n6LANyEU
OWntNRi+TDbExZArLDpf1GPx/WT7LaLO9D8bEktCNYLaEPOU98JEwfwBAMY6jkHrab9aDBWhaVzh
gSn0QFews/Aw6R0egWSvEKXVhCBlPZxdjzoemyeJ3q8hzx9zAqcF1LaHCpCg0HJizc9zSf/tnJUn
/gnuKzkOSw8sLo36cv+FkTTzryRmrnvY5EsTqn+68Rvhe3LMm1hVVGZEDlA0xpz2WhdjRWd+ttlh
iSSgypyae/v+KxM/XY6U8U0irB1cSXCEXJY+3SYFDJ40XUpf8tj5RfFX+MIoYeSHit2QAo2UF+NL
Zs2bCH+ghDO6NOR73bM+UftL71HfM9keOHkCf8dik7798ZebwQe2zdVhlKazk6x8BX8iCVHHK+3G
n+RCSOh8PibhmGRKnQJEBCtgJQl2SSsNImYd1wYx/AN9T0hRmJwxkbwwU62zn1KGYpYuKibLmxDa
pBtttN3FIxISfVN+nJ+KlFEFCE04dDMOi35rUp80fZPMynqwcLHT8OsO/5um7QoLrBS4Ygq5P+ZE
CCn8+07HO8/KHtS09e+39tMBlOAPYqkc5nLdqXeYoLyVwunNB/hF74mQIQBOuCBWi3bU1r0EsC/Z
sjpI8UNdJ10KZiSrFjHmTR3FO85JSEhSgkFTKZUehY1T2qGCTNEMVoeXUD6LGlCC2qRU3qdyRBAr
O5eaTyudFrsvtJaBWoi49WQaUJGAdF+gGjWh+q+TY1ehNsxJBOYH9ADdCnCbEPn2o3u5vliGUjkH
gm1bpsJxFyh3QXR5rv0av4COW5bgCRCBuDlqfdNrKF3EzrlXVbDqP0cs7Xq25QhhYtpG9jnoIBUq
2Z2+gQ1lQx7aMSTLnJH+cVthg6ddKE49LPP9l+v+ATxH1tbaMPNoifIesITjTcgiE2Ftzu82iJBZ
u2nXsEpXnXiWsLsM8Tvi0t02EDjagGldzoRyqDDvYxTm/+0n634jQXIGJVbJxrSi2Ec6F+3xwpEz
t7VY5ibd+UlGNz2I0SBBqcw3d39gVbi5OenSpj128HoYe70gBNtNyuBnm9nP4UPFH0yu4v+4CkMH
hPTl7cZnBUu+FvWm5JZNBwrEU0IIb05+JeYFHzlJ2Z4Kmm+FOH3QxR5EnIPCCOHEHR7yNfXdH95v
tkrINge6Z01S0oe5Kxn3tXKD2cJ30x9R74JMaap2chz5Wadjrvau1zaxeM3UNX22Yi/0kKP5gJLN
Q7qHmEK1wtC3aXVEh8jcdcU0uW71yswsJkmL8JiKHBP9/3U68rDG1vmNQX7Bc5R1TFv5P+uZV1Wv
axJvf8Rce1fXb7fgpBlHfy/WCcqb82Xw28tZhWQzOyZiKdk9gyN0WqsWkvhl2/IQCzDoQa29q21G
O+J6HLRMG13RCmdrfxjHyQRUoulF0Od6jFbvlX2OLZ8kCTXI/iK3sk96OyMIJ1zT4tq5Um5U22M+
Gs0+m6kDMREHd8yhWyfjQnYGSDOb50Kb5AJPy44SRVq3YWgrcX7CREs+TOI/33zWWP8T4SLP7rww
/j0rzmvhCqDNGAyBKWM1qotiRmyipabGQx+cavl0Qn8U5dzOen6epJrxDhpFseXBER+zvNix7MSc
P9Kx3+Vt9sG84VbziL9AOmeYIJZ/ZmlS1KGuXKhRorxU0VtTRY7YlOF6FPyg/yY7pS81d5K6YDY1
dFhCI6MPOXouHmKQnZVVYXwkXIpFj/XPuI1OgzXK9tQtBUw4X2MJME8wBG8s6M3wuS98Zc6/u7kV
34gfRfbB2F0qR7wB+o3vUSkrwqgKaR0Sb3MkDf34WDIUmQoYZLzqtBylWyQy5OBZr28QtiqGs3kr
ZW1T/RrxgSyB+dgFzZlQd/4rnB4caT0vQ3MlCCdH6DegL8M2fJSd+62a8j2SgujviT0fz23OoFe/
qRamhYwu+bPpu/NdpbZoSDAn8ors1y6te+lIuttXJjLlhyQCd45McNZMRjuJxwxqkBvuSJQuv8s2
Iq6SJlZju0OPKbIM3RWFkEw3VC4APeVRD76LCeeHJOMKjIpGE+5EF6Jocdf1Zn2nzU19r5Y+duxT
rPPE5TbzuzpLqDnyyO5V8HpY62IjVQLRIxGgll0Fno0zNU7mP8bPFyrixUt6n02mHkIlFs+Ci9AG
GnF82tiztLuNYbfwnwUK1KWeK6bGmDbh/mxOMeG3QoaRoD033GYE6QdSigw2W2E0mBoY4dc7nr0o
/ynG5wwBi163UAs+ARs7pcXDcT9PVx5mupHB2Fs3oLqPk6RgYjepVkgi0gh3XcAVyjiRx0nKUVXV
8UEh4uVJNVSr8KXx943CgTTag9LGeEZ0EmgBjEBzFYU5SilsKKbdraxT6dq8rU465UmAiB5YIsFZ
vnPVguosCIFiKQWh313VKpPtjJQi9Us2rql9OzpTOoAweFUP5sVLjJ5ZDZF9IwPOl39K2UurKsDf
Ulny9FrPlJmRTsOP0QefvVv1rGdzFxHOtHz0k8KXoesLjbwqzD00UNIJHe7I4axV0H31aY4MULCT
sS77YoJ3kfALJvHYR5pysx+qRNaIQQHySFOiUP66k1WdmbYdySVWT0HYGRN9iqDV4MpL0+cTy/Yi
aPC/z560ly2rTB+Pj5PkyBxIVshX/duo2gHiN4v2uumsA3uFeRZ9hZ8f51ybjp94XFaLHKNimH+W
wsUmFrmUBzsgXsE1v2La8tlVEp9FAjaZSYeNxCpLl8YbeWfaGpaIot+vEDyaEqMJ1RBkBETQmpfS
naO4/kg6IsedHNxm/DrgMmgSxogVzFj2Ac4mQ7M0cP7/5NoxXNv4pTaBI2rNTTaSmGSitoul6nHJ
IUQDirH1T1QsC7hgGYVOv2YUCsg450l4UD25n36Ib3BY0S4IgNQ8G/6/a6A7FGCh+IpUR93R1e6H
WY7F6UcfUlNGRXNSJNdM8LVYQaZ0jxS40Mnv/Uy3sEjIB3X3yzkXvRdV1oWpx5aqJWZ/T2oIZBGj
Qfry07qjGTS9zLMeB1MOXK9vSYHoHOMA/qTLEtQkycuWDFnlXNam+wfIR5zbCVr6k59vuW09fXyp
f342YmSK+5ebdbF9pXgJUanU9P8tBHmLa9ixexbLAPfXe/PbJRykYOZKYht1i5lcQ4VOF4SF9y/o
r+3axjHHEjfCGyly1rc6qBvQSQhmblNKEHnppcDxKDlMd2IaSjEESwK8cFuvlF5qXHkZQsCHhuYM
3NrhEOn0B4+xAB+REVHBfSZ0TzsJPzzrInFp8/HCl5kImYSQSaa9JV3gx33CMXmiz1wMPxXhZ6Rj
LubN1gEVsboQnnKEQt/J5YqH2Yw+5AsJMvTVUFzhvWstm4maG7jhO55l95J46k9RiW1zWcLrDpAG
2UrZ127V9kO2l389NKWmx6znJHDrfymLfUO8f+HrIuFJkEWArxQojLqxllpdpyA8OCYn/z1GFwun
Tc2fwaUxpRSG9Gqg4eWrNSz4MGlP2tFWsttvPKQIUSpnFRWVccky0xrIXhLsDQtiA7qTJWg3EEp1
uKIWHkF9kOKxfYYNiw55obY6djEhAQXJ+cxZHcSI0CRwfYRDHU3wDL3bJT1v1GvB76CqYc1ovNk3
VfVp8IKqVXRd6qd3i27bRZtUabARGxXbclckmXKyiShRSV4ETPRLTXfQkP41CxayFNC4E2N6Ggbn
zU6AKsTiF05otyVzdLFeEcT7ULA+jMvX+ocqoXZ2hq9/REAlu9/Phnl9J4s8n2EsJieh6Sl5+TtC
BMXpqSiKdzgzZfqHbkp9G1bi3ge0EjGoZO+bLreNt0udCfhWtynWBRp9nATgN6rPfMYGqNhbbfIX
wjDpaipXTnBaLuTknzN0i3ADx3VMNqOadDcg7SVPBmtjcNxy+io9DKHhpBZeHevoNJdDyW16UVMA
/oBD9qWvVYlNUvwF90nn7fb82LvbCFQ8k6eU4wP4rI7thtnUgUzQDaOf4+yJM84z6IL1xRJx5G2Q
2ABr8L1Njo1tOjIjuOnxnxuXG8NdSHkgbCIozqwXCoOnP7+sBiX5JNGCsR6R5JGbJ9n2uPrTo+v8
rFCjlvLZJyTVms5pggvn+N5ovAh6MO6QLcytCxHIR2KQiCuhpweBsnVZA3HBQDNofdtkYNz0EZg/
IoRxbjURgKm3gp6K7qFlvBCJ4JOdA4QXL926iPcl5J9/vfjqKZ8GzY7/Y6ldJPSryk4FRtGmVetj
JAw00TDwdjA1DviqUuuCRrJ2A3Q2WQJ6Ud480WuPvpKW+o9vQLjVCmj/VYELCWrxuMv4arvscuwK
4G5M2B39Fd8IBNzKXP6wzCmwccRtzOeIdWMDnPkzYo8WWdvRnd2IwSBymnag5W+u4lh8wTNbg2DG
YQiZrspkSoMAHcYuqB3KkBK3Bhk0CDhzZFi1X1GkwI+YL6v5ySNYLSOuk97+U93c1TpT30hoMeCi
631iDjsNXuA3G5mqWlLktf13hCVqlPFqlfJkPeRXQ/rhxoRzFgVXuAi5mFbYQ6CwhSAflWpHCVce
XmylyOUfjICNV2X2HOxu5OJ7QFqaBJASAMFPSSkvSaFjYt9CXRVAqhTpH1Zu/dmnnmkvLAFYt9Rx
NVleAwiIjb8UqL/G5iQ2dpXLtxyStNUGiXbozRMcpbj6nqNYXDoejSReYdZVMZhUxXe8EtFX5IzU
S5bq74gFUUEDS2qqh3EgIRDb0nBeml+/T0zPp09ZZNX00pOO4+auQ+9f0A9s5+nDoUlRsPj/cNdX
NAoFdbSm930uqg27F8VY8Ki8t6ShS3C+Q6kmieSLL22vctS8ZpSOZ8VoU60ABnov6SRkEpwiWGTv
QEV8J1TehTo4ZAVyIQpl1nS00mMkDLbOjVcYfiB3qrofdE1fLblGSNDMGbFxrJjdTaOkMVvTKSuc
5/pyP2rcxUe7t7N8NodGk5PqGs47zRh/pkLCKfbBpSoVn+GpsAmYhhjLBiF0z9O47de8q+Hvmc5J
6if9Mac8PjUWjrVMnLlNN7z+lJLWLOFudseokB5hCLZV+KOo/xa1gR1h9ILfzrfwF2K0DmkEJG5e
pOSIidTCckDIgppxOCtpUCaf0Mx9JuLMknKIqiE6un/yD8HxDWCqR6EcXMS3ySRFeVQDx/HVSGO3
8gYPZRIoMI/CEcc9+TsPJxLlMPunlbz134uURi++W1WCNoYfNCgwx/qFX916uBsVmLnI7BOKlob2
VWnHnJ2t6K1rP2nl5avRNr24XbO3epjU5N1qrtznW2u9+ZRB2eN8/VS/K+pQX1daD0NHOflAOpF/
Ipapf3UYczAQ8pTIgiJGFsI/F9UEBlSa8CTCEZimWPvWyR4VfNEjzBDs2y9y4N7B7IeIi4wxN9Qi
+7KzzyyzVT0hNahX7soNltb4y4yGinSan0nuZ7bTWRKivIZ1mxMe74wcAbdeSKkVJNS2BECGm/xl
WMLGloIK2OdbHlWFbOJT4yj1dbp5lwO74MJAZVdr+GXUadlRN5lRsRRyIAVOqn/sZwUehR5aP6aI
HKGoz5imjpIsgJJHuPocPxXqKSN3+nz5x33Cyi34Fef5FuaT81LuRd6FPJ9CxigTm0omm5d+ec0R
ep9KQpjRJn1NGxbVpd7Cyvg/GyrJQky+wa6F2MlgZ6orJfA521BFlAMLsqy9/2JEOvDOC7Ntg46C
GwvMVnnFs5O9WjlMAVhVJdoXD5pg/Fw8LLj46tLKV0CMFcyler3UzXzI/3sAloVGWrv9kp1dNZgb
+SNBnUtiPL82t+wh+PmfwpD84rj5/CjPzl52M4RVTygnYvLxhN3ZLdrfhlXhhonOrYpU+fTBFZEZ
KbaQ5VXyQqiQGFe2LoaMnlnLPEpRlrT+42OAfM0pagXy/JkneUGsY3bQu3SJkjGSSdoIm/qFt3LU
xYV0jIOHd2FIKVZWgQAhLfK5as9WgXKwIbWyyrRYQ3qdbjbNX+3Jna4mnF0UnhiP5TI7Is9NvdwW
1lO9t2FStNXWH0jRnacLCQLyOJFri7JOVGQTC9RAeWIczIbpMmvyLO5NXFl2NyU3loP61MyytMlX
rxbX4Q+VgfUt5Y/BvKNMwMZoTEfAo0+7DDrhEgLaRW2UEKyoczmL+ZnlUoeC+sOI9FXVPKorClgC
zW40usV0M0gYlw6I67fgUoJ3cTdf8S61O/m/ng66gzl1k/SSHDoHHnVuZvxEtV4tIcTSYslxbD4X
HXNId4OMi0GfQSTxI/rddv4pcbMFGOt/BQoqF/bQJY8WDYTVQ1TGFiZPk1wv8howY2BYXBYDFgJQ
V6tRnKIjRFTAnTCEasYvQTC147AIRDkpdYba5Rcjpse0NYEl0Sl87Gjo0u9QthPaym0t+0ZbkbKQ
8gePrHAQsfeOVvR8Q1kAjPTY0CK0p1vp0Hj8JpVvoKC/tMbswuWaGpedVvNHbn9chIo7XM0k/2mq
i2Mu9uwopAOFsRHnd3y4URMyLjS0WX5S4zbOD5NfXLglqltQG1EHdBGQVRqJeeK1fqIqvqHpa91d
tY8skYryFw6s/gk/OB66XPxHW+jjjQGEyjsbgNuEN+HeR8HYaTTP9JTsy5RuIwzEVzr2JHZtwIr8
gJUTZPu0IVU9jeuoM4+K2B2yLCFbZVW/wvkKk4I/CrO7y3LBiJVRxIU77wHiHUSgbLteteH42T6K
jrygVVajpzkqvf6COqti13jzKz3iwxv/A/GK04LU/USA7ErtqyYe2Hh/Oi0wGrWDV7aT5QIY5lGH
leBNhVBMYr4anHxjeb/NDMNobO3PM+RkTCvU/T13ZlH9vAUlUMur9vkQT8BsIV8mPT1fl0hxAidW
UG6LYrUH0C9PWTWCWDaMzfcr96KFqzyCvdgE9YGKU1mXYvJWIXUgT0lBGDT0MbenWNS1f/xCYDzm
GOYCC3jF5CAeU2q0OkvlCM2E0ov9rCoSMdA6pfRHiB3p0BitqP1Zerb/9GVxAvBKrBYmgAI2en0I
bnTdjkh7NbyQ+I1drTZqtjHHuZ7SWKJg8HNMEqfLp0liNw82o/MXxGySbNBmCZbNPGsxKB632pFi
ONU/JbhUxTQXgCT388m8sl8nWeFTDLvgTF+k121tmt1NuE7n1K8+q3L7mEtbUVG2zei3+smQLNQz
PpyaYOPKPNfMPfhN6T5RrlUhCiKf+EARr6dstjoiGG9abk5QTlVBq9O1hQkeZ4fUQRBsi/NiWinZ
MIrzO4p5pzbzABwGL5gs6sDdK7M3TSSsfYFnr44rbCCo0ELUvCIGlYr108lM+HksZZFMekQVzSP3
P/NXIaCkab5/AmhPM+UBc7d2Ohg2D51NKJ+d4mrNOunqNrw9OhLOHjPIXzjZqOE8U5cMe9p412qh
mylt6gn3iDkJ+qDeUvKeWScSTLLwnWU8LZDG5LYjVxNL0TdV0PBCqhLYVCsr6nB+qvV1axL5NBqO
REa/0yOvKRomsbOxiEv5Bpz3e0ogq7Q4T7sgnQ+u11MOixafLPOvH+yalJxuR8Jnb9vOfXCwH4Mt
gY2JsontNkhBz6jf3O2onqZgbtj4hQ2/Bvhbpd7HsGFr0dKNdJjposbCi/u1rahjXUMBHK7JCdWM
6ncDqD8TIseJZEkez12DG3AA1xjH0fPq3RkSthZbY+iIk3L3YDUruZ/mzGERMw+24UKX29Ww2Gx6
CsQmdCju3TXENukTPRDn8R2de0+9PjULQlgzNytmgyvy538toGBCZbbXwr8wftYdA01T/7Cd/Cna
mJJaZK98YBsKg2zpqriDiflavzltDkkzDqvDQ3Z0xy2uzNoIKcFsW8ZINfMjDSnIsFQ1J9G2Qxbv
14Rh2objJrfvf5Z/76HToKSk/LoyUzCqLzwm8UleA65Z/M0DvzX5yI5Gz5wHdk2HMW9QL56Nux9S
61aHCSUtHWzgJptMDFGH+Rk0jB6+4XdVvIqAMf1g6ILEyENxd/XAe0o78RryQbVTv9fv7Q9+TPyX
jfzMZzUDTK8jqsb7PLbEPaBLI38TdObvnZePZzfByphZflBckegLyld/x7R+EONRaIDsQavS5C3t
g2jYteQmvqNv1FfcvSRdbgudV51fc9idFriQJGRoWGZiLlBL0z44o0zLWbARti+A6hiERhVK/vOa
N9Dn3Bd6FkjiMmC+jyOzRGw0+mEFnnv4GSGw4RkBV6fxMcFuborvnM5WAw3GM9KvAFKp1HgYC95g
MiyDF74TjN1kPqdTdQ7/VaWE2r7jGIIp9x9NGlB/zaTtOz8WtqApIK/VZiP+VDSa+GH9dQnSKbVL
IA7FTkXY2adqd1AtzGfD342swEuPh+CYvy18DUrF6cYD1uLbW5oKIi7GcXbs+1ujHBJu3w4wsI37
iRkcMH1xgMsat+TDpWH9FI5vdaj7hm7tVLIbQCkPI/FMaSQeDf0BKDAtto73RY6XZo/CwgDjLdML
+2amJ0HvMAiEtyf02gh7oKvUwOHDIlebnM6M+yejdk21JG9lkqYPSXoeaqeFqVXxpp/cArFNycaN
7ZsOaDTsCPw9t9YzNqyek1QPVwaAptBcuKb+shxUBCDWOGDr1gQiOWxA+F6YFEmYmAdKk10qv19N
zKjcBXtkgq0RvsxND2xE8Dkk2awgwTlLRgrhTnEGoLjQAprkbQVOEBNDTSZRhpLgEaP1qtos0TBD
1ExyQif9Ro0c2QF+YTnEnYCFNM5C64vjAKYUofIg1zeLSNAle7Gf1GBBF7bNHHhD+/Lvvx10iVHt
UMALrYSLZ3MpuyFKcsTRCcLzFtOVUQVhB8zhchpFxQtHR/7kAb7Ze4JTI2QZxRxivRMZQKuUIpRS
k7dRZwb5ggGeTw4hqtCXVdzLBQMJgMog3WeRy/trb7yr3CNm96UWou+bYZ7orvLfvFZ9kq8CieY3
fY0oY0ePcNSumhdTzSsWfiQPNPV9BA7gx+rL14rfADaZbEM/RI56trcoW8v/AyWnWO/ga0MQQGE2
0V1Pm0iCL2N+j+ZtIfEHdTtYQ2Et81UkOb7pCQ3ORC5zUxQiFGldWVvArzKgEtcKgofsmQuWxmOE
++Zsc6loe7TpoI7nhaeHXM/7UaooGwveDMu8cwMH9VrWry7F6SafM+nLOdbgNu1MuiI60ozZfl5I
ZZlSzbHTOGCESyNiVM6OVGlwgZSxGQFO58NK54y9jbf++vJs070qmVtqR9fcX6czyqQCS0Cg/i9N
R4mD/mcGO9u7k9x8nmOlPsuaSsvhZWSaoTCSq72pgm/qv3cO10UtHXbzIXtk2LCfdgDbGsTIGoIs
9jGWkDijWCok+kob83sTzFSo/KhWLZKZB8k0iIm8M1B/Hhq1wbPPthg2EbOEWFmvWTfgnqn+zmde
s3heezfBuymZafecQNsRtb8tNaG38GoKT9eFztESeXqyq+tPIfOdnaJt5yHPu5cyVVQyEOF8OPVH
C0rM6/k6O5D/5YZa89vrfwxEnYkeo0YHLPFooDQLTq/3siuZ9lYkGC1SgjjdXlMUKsLTEtnHmnyo
QCia4GHesApjHs/o0Fm+GNsNDRN1he4GAbAocdwxki1MeQNnMeDvLQpdT9gR0TXSOnREDcZQ0bz6
Ev1hcDjgKDY0quE8WQFDPyhLMLfTYqmzIAbBXp2feMAM/HZCklBcuerFLQMf3L/opq3a6uY6E9jl
3x2xHLGf3gUa4b02t5960bg2R2XFgP6eWrsVMuz/eJd2p8szwp6zBl6Yb3SyFiEYjNDWwx5OgvFM
mfevwRMNRbPUeX8bY9vB8gNliISegklx3/t4DjDxsY7bmgDiHaE5zpJ6StVQj5akIlBgya1Hdj7h
9HrHs2jVDiWL9mMAoZJjYW2qPe+M5ZfCOqYgeJzLUODYAFfW0BUSsnrfVsUl7dIaFenLZBJnlZzW
y5eJQolA7yi5ma0p4dMqZd6J2R+gBMqLw8oYcRhboHPQo7I7WOjtdV5Z/4EUEsEvnQDhNXeBNrNH
4c8mprFo6QfN4+rmOM4AaaoRpB/y88ZYtrzjT6cyh9X48CfrEQlCFvjT2bXsfS5ChBYgdb9XiF2Q
XfrNTmxxeTiFi4a39SQ7VFCVI2nrYDRRv3RmxTVPV34PZkgVS1VoAHThugLQfRfQ1DxEYMWEG6AC
lyMBvuyKFDeC8rP3UpaemNQtOtCb0PGknv8NaO4xThXsPwv+IPQ1QcJIBtqnep3KIIUOPvU08u4l
tJwiDoK/CMWPojsMEvfzqe7pi+m+DyH/vI0t+49VUeTDbbkFcXrOht1VJUxY2eawE+vYa9wSy26D
j+eywOEFY37DQT27PSw0EaD10YbEmAoT6szNQ6/JlnDWDZ6sXTKnYDlOrOK0peAJsYFJtj/IOqLZ
KrR0Aw5YAOqm+ooVEDbNva7uJkcnPOfKUHxyUr3xrAxycvYjfhF+JkOvsKwuTbfn9xSHH/5F8b/z
+MzAiOlKvZEM6mNsTNJJFBei+ptqzqZ9dFZHTYvHAKRWIlldi7h2yqn13bYnNLn2vDsz2tOb3S4X
FtDSBpZRtZhzjowIsT3IqpUxt6UrVVMKVdql/R9KLIm1Ia/WDy/KvT+lKWbGUQGVupfk5E1acQU/
oTm4M9PjMi3mTcJBxONRPWJRWiJjdE3/viTx8ayLk+mB0x9Ll3OKaxC3gv5/qAa1mbgM63zmpTZZ
bEJ9t71ADOin5ZKBHcIAc3J7nwdmqchrxAFP5QyHSmo+iUdSaLJbj7glzhs9N2nxxXz7nXfV8NdK
nf68UPzBQH55kHo8oqvgBOjUCr8PiJpuiKm5YU55w216J/Oe3fyudJmcxx6MOY0uL1QriLv6KaNc
8OJdkWshenKR0ioyKus+T5GEs4Uad7XNniFcip7BSu4U+hGiLSySTQv+YzzB+8GkOGK1PbLs2zaX
ZlWhxW2jUIZK4L/H99PMP4Yuv5zw1L/5ovosnUgGW0GJXVz92J+8wow1XthkYPiXn1mPs7afzOj5
wrwnYVuykCy3dxseH+lCNZNpFvDeqRNdPX0ywPih6TiTXHttSCSzmRYoa0LC8nw2bWLFxUxoYIZU
tPXFYORjDPZXONhDKYDrS0iYbTC0I4zgfcYwHEPP69GsuaYNYAcSNZrn8aFIkDa9a4cWqcBI+q6N
QWEnVQsgyw/JZGm+scYWwpqcO0Cx6WsuW43Sc34vVh9uGsJ3xO5lP+uPrZGsQSR6vRlcCTm29cCw
WWpSidpJSDUUknHt5f34qrcEfkCNZohbnLbj5yYk22Re9lzNDFmxCmAx0COO7bHHcL3itiOg97Lg
2RF50gd5rW8sp3z5aVT1LyggFAcrQ5/KUpmAB6Pl4/aDlL24BhwULyC9Mfi6yL5gma3pEn3zunfn
mVZOCVxL5Gp5Ee7lQCa/GrsfvBrdV+bVUQAeZwf3zxRMNJa2gEjGUSuTqNfsknAF1+IGkT0pxoZU
KBejYy0Fh7m5+0stHgXHT8JQThLK9gudk1ozJ7e4m2i6vPPMTdkDSLAYr+ZoLhQvfDAOJJDIZseq
Tdcs3xQnuo8mKaOrc1W0PLp6In5lsye3Y9/lvIGjCvvaH74zQtNr4MQKx2L81D30OMmNoPsWWt7m
+WCC/4uaZ+i/iWi/N4cgSkOZTQDQXSB7t8yDXGl79mjJYJnNeJiBOKGQWKGcYgRens7R+ENuDWCs
FX6kzp6ZWhk3ztlV8CY8ZgZaMqFP1nJ1zP20n3Igij++M8P4xsTamDlZfxvdzscfe7N3AXUxJgtj
fmux4YakayZ6R2PPa6nQj2YzXke0jb6pu+AwLi9Lcquq90YIejsCI4drNHcGmQsbMsyxCDjF5Ncn
CoQBOGzoeSjcKMavnNyKt8M1vIUf7aGHinBnrLVITKD3DYF+2jfbnInWxyWtCKyrqjGWS+zJGa8e
tny4xyfgymeN6StnF4sPdsiSGotyFJhIoxg3S2du63tV3G3+tKSE3hvDMdGjPDPZx/MuTp5Z5w3f
ETuR7SCu2UJgD/psktCSTd3PGM+kZnZOPRKMjknXy7k24UK++sYvbXmTpDuwShQwbbx0Xtxgt6Tz
YvmWMF2pBuuD5t8XemwODlBUumcKOWe1wqTGce1R610YvpaKJSK81fMBz4Cae8Lm3XjzReozeulW
CDYYkMNup34volNJ/oWFw+WFJUMYtXtmGa+7IMc9s6U5RdHTXma+e+XdaaAhOCLFOzNmIIOKqdZa
bNFCZ8QfFe7ViAArX8oxgXnFsqOPoRT1j0mGHSjonZmapEnzDJIjR4qAsJrQ+iQFdEgII3NyJCBb
dO+6YqlhhuNHdsOMg8mbhY3CAB+E/0dAJMX+Wz8J7BXA6SG2Vw0PWbFNvg8NzBkMoYhMhEZbXPH0
xxsGTWghWrKmwS5ETQDIzG8V6rzUOhyQU7t35hWsx2c+x5sX4gf1+XpJP2H3wlWXSKoYAM1iv2lf
CtJ+KaImMlKbN+YiUEdM3R3QbmrACriBpsuA9/hSXqxVsfmlCdWeZIQl4SGpmtqlC/HJdvdJA5L9
LxdqDIzlter6VMVDYKcf1ppPg5P8mVaycBkwlnR+ku61Lhgor+bx3PuJ2GgHAqQSEEdUyk8gfxFy
lr+D+m23EiYBINQLISvaOm7uml2RiaRdLCrs/A/ckRMXdNKowISy0rlT9lIBgoTZONteKUIXQNFA
wAaDh6zatghn6l+L3qW2hoj+2lZXMkUp60V4roZKMTKMXT22/xPJzCKgKCOhEDVK5zmIYBE72fZ1
xng2ghCzcjw2kHQ5PkU6AEujQDWaqOJle4pLHE0HR0c99salX8ds5iXwXJ05f1ocy7jAZYmI8alq
VqgubReV5Cv0U/D0bq+un9QYeLl4KZ6j5rsLKm3rZ5WgNmOWsxd4MaG8RZxknOORIdQI/ISpzSme
djtRFNznJPuC60O0dvduD0sxjRsrOG7cJcxZNzoro1Uh1CYOqkcHDX6z+RPYLJZ+p4w7qr/fJMXh
yTSpTgBxynL8PPSUEFK/qc2n5I8SlyC4q0GRCwWOny3MgUV4QPBZB0/UjmxFW7ZCCe+eavdU2830
vQNiuffCEvfuAFV2aTAV6LZUq//cE7rFXxSnhyXUkaQyf8YGoRFUxvVDSAEQXmpybg9RyO33Nsaz
kYLr3w5R8VOzZVfbkfKtNAQ06dOzsVxX7k6vOR1xpSodDpVLu+XEfy6bmas5DuRslUaYYSWQ9x6C
vwPXXpODlvU2lFq1SgY2UNyIjB08xYsyVLKlTTO5zO6FA4uxgiR0ba8Mak6LO83042gND0BmlD6f
kHMI4Taz1sUQLuaLd//cPD3aWBey3iszS0zpJOIoL3OoGNE7cCxcKGXO9SkIUgG4isXVnHhZqlbk
YowtqDXuw9AghlYrk3apHliUijWU87cZ8l9mkxS5pAE+AwuV14mnkPviX8hOubviCqtwhkHi59Dq
BQNKQ7V7tYs2GjZU2slOZwtLEoNgfrL4GcMVSF3+khqELXRQYD42+N2/YNC3+suANyU5Lk8LFlav
LZTIc8MPeUoH8Ei/dR+0Pq9jEK4rnwyFvjSnQLUn9vfK0nnNKZ1yTZLuwwJVfklMUfbTv4TKUJXJ
1OJsGu0ZGrD3YOpBU/GSUCGtUcuI17e0LjujRqnmYshFyunTB3jscmDWyR7WrqAmsbnRWfj7zTtW
0NJdObW4tvW9gcjdEE551xLEQWkc1UHwR3JUvBl/fKjqixeOAUCwQmqXaOAc8B0mUroeNMxi3kQC
kGp2JIrph9njjfjBojcrKI+67KmMCei3u0dNXa9D5N+NgRTrJb7OydoOCV65cY3A+qyBkjDDIrSU
T8yXPTbc2gUos4CeUv4NDaBdOC300QrWJLGa8AkXcEFk/GPIjImOBYfTisDQ+3HezOLFGG4DfMhO
7hZ9X8RBeC96iDkPg62uiDi5q6M4iErYeiWquzyCRNFiqHW4KbdkqGtcjxsus+wnIVss6dO1eO/l
2m1/gbyyUYRq+yjKiK2zDN5brcLyhgmmg+VaxcH+wnehqrix23C2lWCwHdkuSVLZ7kQ3V6pZujbv
XqdWBznT0oUlyGbzc7JzrSXHqT7jR87L4TbkRlsm2eHkylf+OAA/IdwgzEd/F5pVGiob0+9LuxJt
9ZNRvwVTblX5I3HmzNnprnHZEXEGTdTmcWy724YY7LzCC01kJoGGw8wsl2R506fGYi4JNFeUEYzv
6k+QzIz2w7l931vKDAw5w8LV4NaF70bCpZTA0ZWv9DFjjwRDp14vxI7jYh8/8Bzu3ie/E+GpikdI
Dj5i0ihMnTidvBKEzeW8KwvAuCs8ScPmjEeZevYAN5SrFAuRz4jvgL8ovf90Dg7DgKHEh1BBAkBL
KYMRRhY8iXmWfBBxjLeAXAX0a/saqgYREBEAh+2jEunSxyDEZql/1HC6VVrCyG3zEHlWKWRnqpvr
YueFFhZ8OhflkgkMdlqSJB5RcyB1AR42aytuBD6cHblXbAydvf2LRAbOvc2byVXVOaqWU9tKva+P
lazjqVftkEgM1/v49uP89bwoGalPnnNfIrFYDi6ljTae6ROV4284zXBdJ1Rl6/+9xvg343/3P/tm
Dro5L5/VYUiw/HDlV7P6hD9zDO40P6OgSXRY3wN7kmiqm76UzgWullKzPQCWU/GuTl3hhyodMHFB
fGYZEkXmno3EjTXhDJ/RTW85Mrn10v44bQS22YngZx227kOdQlqiBH/fcD01p/pIYnTUm+9XL/UI
Ga6XHGenow7oKfg0eJZhxX1ZeCPa73cdWklgssjhMbDeL2HYYOqOhyquKF2BCeeloAUp6S2X1MPV
VFTPhOZ0GaF9Myx2p/NOmg7tjuy53QK094Y3/AaWLKZ1mjaCvnTu6sbQaaE7whrAize/PNiHm3el
CjFXe61yuU0qCjICUn0IYLTK5Sih1rTOOoJQ9eIAx2w2bmfsu7X3yuJS1kRB/HEjM9nPu9KW/tQ/
D1YC7EpV/VPgFCMEZerA7hWQApSiLGG2kl3Jk0eKmhxsbcku/9K8T4fbMnaSbjGfFFKQj3fiqyJw
JRdZtFGAAYmPVdWpkdWlEiXMxFryMMZuK37Z15MBhsMlZ+d6xKZ1TKHOlS0NwThwtsKHzgSSn/0p
sSBfbI42v+U1pLfHY2aS6iWnerDKXVO5Jd1DUNZFMKAgwm4Uxx4vEpfISH7XVBfq+m2xdCljv+VS
c011+yQsd0awNcFAcvHDrXLJzhygDXVH4pqXF0GSCLQggKVqCMSyekOu7nS5Yxkw1oFrPRBKPuee
hvi/GmROhZ3FEjDMD8JiTi9mEy8qd5kpRMe7IOrirZU8EB8aQlU5vF9ZMELTrBqTirmQFPJuNsDB
Vx4vG7QtUGp8JaQwnN0dY1q37PLzaPMpT2fAxX/srb6jmAYCXhWoG7Mn9zlHc09ZjLLPFS6kkXE3
lkMYhcBED6joZjrs/k5A6P9mpoDIad2/YuejIrllOcVN7MnbqD2YrgNIKQiG+Of3yvabNxu7VPX+
p+dsTQ8EW53j+v2XXPj1z8uIy5iKZ97hRdDkP7r0uU5rE8PU9igNSnGIiDRS0eWuMzKL8J0VH/jk
xwkdCec3Bgj9rVe1Qy+fM6CXP2EA2yUaYYcXeBTbBJJdcIV3iOZMssmlb9zGq7f+wEFCldU+adZy
4zilNNRfEMjt3lFyEJ0w8awlEznN12T44/04v9CtvlPZaoEv0bOo2rJV0aP2NiB1U4aBkn6Ngs9Z
yW81eu9pBjoynAMTBcijgkicqSIS5WYF2ICBTexRoCtUqTvNzcqOuPR96M9fY+043BBLC5bFfrb5
v+ibWq2opDVp7wPa+BoNL6V0FAXlAxkwYBvgR0Zccs43A00UiuWBnlRbdFOxQmWYmuIl0OG6Y37n
YGmhB5h937a0wdp8siDCsR36B8nPOdz4+5cKgt5cqOcAJlhLGjILhcFablpjmoyAdP4cpCuKnmgQ
gD/LmEtfF96imLjPOTWdJb2LfECBk8HPNaBas4Sk+ZvdevwIyoS5jPpBEWKlRa/ezKKisO7MDH3o
9vT04k6bqpNIYc1TH0Jcw9vLyxo5Mbw2fTKLYvVcKzUzp6QrqS+IeGe87iJ9d1rRWBb7GAQI34sE
tbbvmzlk3Q/+sfYG2JYNvFbCObh7bJYVc9zWUJNnjCbqX14iHVazDwKyL0EeWr5uhNhpSId6IhQ7
lsDmyNbWbMMOrNAXFp01u6BF0v0E2kMg/50I+zLPuKPkI0dYBeXTVix0I8YBEoefCM8fcnaSijuD
6JSoYDNqM28N0aXZsni6FnFDAS4mcxu+Yi2LeZd8k5ujrsmcUAhN7mqxAmZ7t+uOWRIl0W+Bpe8A
8WrIL7iRDzCB5luCds5TBwyhqyDZm88739tsj1TbZvb7ShXtCcEKpyOMDqan5423sibmhxX+pUTm
vrwI1+PnIVXUZel5VFqGjNNGflUoTA8A1sjX4MlANSWHMIjdMSAC8G6MnTcx8aQDeFT9y2fNt+R3
+MvPx17ZoMRRqyWrLhYoolBMHq4OB2wqkJIZEFAISMt4QZghqitTORqMs5ll9DlVXq5T3HK5gRDH
Zb2cmsSDMFb8nsYrqAmPAcENFqT7Ypm7tkpskZrjHLvpBzs0O0pHvqOEnWjkw5LR/JrbK06CkHB0
FhMh8bxB/UNi8olOisc6Rsmke+Q6M6OHtSHwLQ3Z092AOTlIRAupNm2sHppEQ9jyuJX5o/hV8azJ
7X3NZep2HwSmly8wlV8CJXQ6dByQDdOziHWcnAfcc3SXsfs1Mf9TU5WGOb999h+I7A9NzYdf5GCu
F9I32VEhseLVxJanYtyesvx3JTTNHBVvXsjcNcymxApuYWpr2mdmgutaz2OGDsltgdUy8nJLTDsK
B3HCIbDAMS3lZGWFu+iVxFyqunaZL9S7QUrL8oJwTMHGQU5gEUQ35ORd4o785pkqXhxxajEmrP+f
KwOXqGzXprLHJpoO3Zbb/RIElnA9+rXQFsFOwEa8C8ZeZoClPFNeO/t65YH0OUZGDu+Nniz6fSPI
uGViXzzQ+d9o+RdUyWQWdhCXqKIhADIco3U/w4lT6toBJgN9KvQNCzsfhjA+76LzTFdi0Q6ZgXcm
okGtquyDiwL6N4v7ROHag5FBIDvKiGurpIefCNVRb+XxuFWJ8zecLCNufqu4OrerSmXjFe/KBrnI
T9xNeNp4d7PDGuT6dc47zsTkI6hxkJ5W8BKr4M9ueLM1IZwcbF0lKddwmMnN4nwXgHc1K95IQXb3
jx03m9o7RRGGb0axT+XZ/bMHIqFmhKmHJ4aX7PEsQNh1N+ZHQe+ksbdAd7NfNi63XbjNok3Rhk1o
+CwP6v0dDLRodLHF39wwCkSlAPQcvMrrURc4NnBv6olp8x5msfU88digtMhsgp8kjKktY8+jankN
AO/eMzaOt25j+ZQ4bVFgqKtCkGljo88qVf9K54Yv9IOBPT/kG00hdP5Ku8PPlYLWRxJZsYPqMcnf
ZD8eel6DJ09wGSxmY232Cxlsm4SZsRK+Hn7U8MXgCFIRi7aEfzUM0ey455c0TRYTPGLUs/TUBtcw
MSCr+YY/E6OVoh5zV0/ocmQ/5U9wyfe1UwdaKegM0wRyp3C83RZJINtnOz0MVGrW2L+Q7P9rX2Mh
MUVtCvl2ZjHbxD/fgRv3dhEVxdvZQKd6iTwebslxiDaFsXHZ6MeDvVvcIvrHIWvA9HwPUGrR5Xg8
1kff2e9zi7yIhuesvONacieD9UVeNZh2kao8M9QZNbC4g3RyYGcVSKtL8mbA1svIHgdMZUPKjnSD
KOEzpI5MJ0LwrTa+0raf1Ht5EE3cXZGCJ3Qr6+vmQ0S5qpj7i1SFFnhM6tPZ2UMYR5EuGmMHeOAL
ZqCiITqFnPNBq8mwCGVeq/6G8Xaj70SlLyWoLyoC9ru0NDEh+I1iqben6gT+J8I7BLRJQrzIA/YZ
l/tbv2ljOd4Gj+JXdVW63Rn0PbquaaJLSHb0NcWw7iZ/zRW/DfrFj9KUbggcn4hbjMGGCBV25neq
7gKyIWgvf7HWRkcX611UVJ8rYweXfvVzb+Umbt4jTqmjTpaj/oduRFIGBp9X1XN8gMXYpu9npfrx
4QpwKNeu/KfMZul7E7BDoLctGToJK4bgYJeKPUTF42GQ/FYbaNmBj+oJg0a/kz4+8PIL5g4k5/mu
g7XY0zlNa1WIjSgrfhY1tfPleZ0bZpYXB5cgKaTz+TUz1RjxNLYeFDiWAEZ+8BVKU4ewVRKV/gNF
HQRBIT3XhD0AT5fzpreO/HMUY4GPBKS8L0HjuSibmUaL2tmUu+feMhsiJfsK4fn2qhvUd99nbQAf
knA60XMhkyarNLmRQsJJU8erZkBEiNio8ULYWzJKqD87+xhGAz1YOc5pSYD/4YxE/hgGgkGojExH
WzeqxRLpUALbMxh2wVdfdSfrCYD1Qpf3u+rTZ3zhsFgQCczkEishBB/Y3Pqr0n9Y2SwEurtOMYOe
hcfN56ZNRKtTvsRC8TX5dqThxVxfSlBS7lkHFtpAylg3lW+jTlRhWapCqWOz8akDvs0rtdOju/VV
SZ6KHU9A/gFjhX0AbNLzbnfylgGlZqdpWsxh4CcUwq4gdLzD5udJ3oQmBNtCyAgo2ZqShBPrBK93
961ks/j9PgCRxtaN/DrXQjVhW+s+IvEhA7n4gipY0vzjd6PzEtj6y95z6pvWRtPa4kX2Pqpg9vfA
fXrq0ZAvhv9MRdeIscSFt1j9kuEpzkEB/+9UM1vijwb4zZXmj8Fgci+KX+RWwQpvAusaKgjnC03F
n//kDprSt7iKJVG51NZsAQgbHLTBXzC3NxQI20PBB6r9IoKhXgCbTHq+EtqpBYtbjRCJ1WjV4vMV
tGdvPXewB9TjvNd00clZRViy1XiOfpmJN4qoGFRM+mSL9Ps4lwBg0LJ7mJCwy56bzohL83Pc4feN
C6VF3gFaLK7aTWJC/pGcCuBtlZaBx1d1VHpaBJKU8/Q4n0XJvdqZNujIg9ckAqBhUIhlmmaHvhfH
+B/9Od5fxxPFBx32Bh4NaMt8johZ+9DEcv0Xk5DfinqgHa1cnCOaA8CajxVpGs/XiOA5t3uqV1iB
q9e+o416q2lX1HVnmom0P0jMubZzojFqxGcHPh+5cfj28LzHpW4AkeBBYjKnqQzu5kmHB1IAl6Ho
565GorMbiXrrkkCBdqUNL4N+idCg79JBsFC/+xhTjFr/psrvMxx4UHmNjzE57WOCIzwkfaSe6cau
7hor8mAGi+yGiti62YuiDP2H3A6uBzLioO1I+nWDtMq2hK9LHzr0bWi/ctXVTZce40Jfuf+iduND
t/ko9QAiAxyjNQNFqV7vz6SOkr9rhMsIeg1ZJlY4hMBLfRkm2sDyaG9eSLOsbAzMokpLZAdGyNc2
/RTEGJCvn37lqWkWqej8ceQ9bba31DlPjebUWLBf0a57vPMeup0BAc4Ftn8nLML1ipxKrOs9slIs
dQeYClsCS4m0YT9poaJ1aryxeZdewnTHAOVCQeK16XQTbFqoGakAT54BIOQ+rc9xAqn2AeVp402M
dtYiPxYQ6kyw7TFOVfzZiQxBPmPbvQ5N+bdijrvit7pPP9OJ3uksN+xcQ+zNBtVeQ0xsBcNeu++4
f1S9Nf9pF5Yr1pE4/S8fFdhac4xKXbGNvYaPKCudMM7kU/q27Lm3e3OW6bAvtrIBIzC9NrQjn7LP
YpOdOWElauFe9ss4MWmCy5y7755BFns43EfLlFpRatSLWBDPWWctyyzTP8h94Ju+AbUHy4BBR1kL
Cs+hlDwlnFVqAbNpXcH6PtdC7TtZwHHxBh25xLaBVdmPZzN2viXdowWuCUZsNVtYO/stCBCvJohW
H4O1IawJjfW3p5ZIlwbYVO6j7hhUGVKVuVwsfJCSLo3nTvJneKVPEpTN5TLenAaOSQHczzBPWmMk
qJM0w79ppbl9W8SWYly+8ecfqnZ3e7U+SdFOqg1KTS/9xIKsPJZy6k8KwIlD1Aj9okrWBoHmGwtG
4uva6qz3mAgG9CF50iENI4YxZyOqxxF3PcZowiqNNKMkIG9lMDaA1vcefprf80rjh0NAQ8Bn2cZY
MN1oG/dXq/OjMoZg22MqC1a4dPCzMIDwo1gMB4JStfXkSXS72ZFdwBZv3H7XUBZ+FgrS91Wd8IpM
izXHhIhwAnQPTwZkJO3uAESq6wCQPcx3pn7Rh5ogG/14W2CJKXbr6AAdF4WLHhHvkNf8SU+YdkOQ
2vZTrrpMyXeLffwtqVqgyPPDbG5krgmMCwOX7YR9YgFyxn7EmUNd+LS5mw4JSC6Mq+87+wczX9BT
aQ3XoGKGn+979MQdHlZDXBrybG7/CKd/OaGiJOH2jreKwpJm92NY3YjwVbLEuqcmBgUwJi++teqm
eGj5t6vlDCMgGdi3iSvRoqyXuoHQzMOQiPdwjdlhDocrW48udozzFHzYLotM6iJ6td5xJcMT8dyh
3WiltFZtnrGWtKOZJ+kkf2GTs2tqBdKAXnx3IgSk0NMlwPMyIEprmso7pafaZwXp8tK4CaPUtPFh
2T0kc3HOsb8CqVDpCm7yONFBj4DlXqmWKBqYso5LX85J9AOE8mW83ycu2Qf/LAMjh9Wv8kfQx9/N
MwOVwIosP+HJfzB0Nz76yzXpN1wOyigR91UPoK6mC6FHEWUGBvzdlTjDfBUbkmXXZaFssAAOeKTN
e1P/wRjGigCLwBErvzhHPfwfpevP4XTjedBNwAbf/4XAEAD2nUrJ+PNoINAgtvs8E+zWrIo4rwCj
TWIxk03OX0eXjs4Qi2au+1sbBHWg6AJ3P379ODnN1BvqfuV8qtQ8c2h/WsmBijMWvR0oF7SMaOmj
AcSpoIBb3+POzPcLe58zY5epDWPWrnwARRUR/XXTq/X3/Nx18iFBRQ1A5Cf5TPdt29if1eVpdMIP
ySWV4le+fqet3ku76Ub/9oE/JOYtDDm3Xs1MphNpyx4q9FdHv/js6Jes4RPyF3wkgh7rPTQBnTEB
qII/02gI6K2FKACdR9ZHLxE9eNvzSECkBGliMmz4NKYo1EZVcehbtLdlKwWO8rLrjOnNpBvQs8fy
QTRnKZMd+1nn4g40JtJNyHZN6ZdYOveBi7VM6t4Hj87j641qCcEMEAL17Y5CB/uz3T7coyiXHbPS
VtHGZ/pYOVKiOq8G9f9sGtLk3EXHO+NW7Y9IUsb2S5cB34eOI1jheNG3AEGkL3PrMLGb34xEjePB
FhxwxIqJ4Aj4SX8qj92KxMW3moeSUwh1lENM7JWRC1JchXtIYOS221TCuS1KZoqJa5dWyV/la+dQ
+/qEmhxJTvRrmFQt1zQK3p1Kl1juGrmRN82gNJN9oP6Xs8kRfFKB8LKB0ZOUuoG2xboZjkdxVf/A
kTgLJCAriZDyNIubeN/R5QKiB65nIzjPi4sWroQpNiMdEX9I2pNNZinvT2fzF76km5X+6yFmKHAg
clp1ctpOYtYv3WqtjwDH7qSQJ2loCPHjH8SX+c6/ttuAsq0IdKRblPp8Fm7grvgmtpD3TRtGDg9m
RRyts7wDTKGfvk3ICl5WajdIjBIQXMiFj3z5zle2/Ppy/MBXapo4uIMoOv6x0kBwNkBPiUYU/kB9
mE0SA+V3rLt0aL61cEEzv1sQr6Qw/tDFGfqqLJreeJXSEzyiElTmwkz/XpmxyZSN6i0lTmK6+hU/
uQ4HhJErZwHuJItk83X+pGl5hjf94/tajQVGT042Bk/yBsO/Dpy80Ljj/CCWodYg/OGSaUrQNR1E
6VPxAe/KRRCC6Ok7vAc9uqdNcROXka5egL7+DE3Pg3AtI917A7FtFJktLisP5eFnNcPLcnT8UYsJ
FW+bl6NmZP5QOSO8RpjXCpHYacxiDQQjms9d/5uBnAZ23NkixwPF0iL8I4bbV5LUxNJe0vPN+B5V
jedlyS+9H7BiHz9b+rehIBB2f5zOXIc5Qeo+fLe2ysIeIyYfRNoqhL4J+uajwkQJ+OWsnOfUbo5r
ruK9mid/bPLuokGrIzPC/izhUn+lzZqSYS1k02N01L1abnTQB7w5PhFn6tjdj9gCVToZYRvbO49B
cavMfGasH5JWamwR+m0tLgo2DjuRz/+JnQEJcNlY3szQWcjPjpbgO+tkJ0FTktgql2hF3CgnhGEU
EZT+1gOQcDGYxWYay+1yfWvwUgPrxjVIttI6+19VJQRvWXjmoRT+7aUwH4y/gAdGmqjaEgDa3uy/
BxG/VgZsofL8yCRjcUeVhPrakxzs3kv6zx6ph3nvyXrGiyVE/R4APespxh+WRT77Hbq5xPutu8dh
3ESDNwIaPHzYmxPVrsqz5jaBO7EwnTFDUX2gAyrTPYo3M9mWBLSLg5ZyBVWgS0F2vjyMmbk8Ia/z
COv65Q1UnUqTpOJ4CZ9W9NQG5BRfelt3o4IbC9rAz29YxA+Cx/wiYJypRxuTqYM6J4vPPaUcujmU
l5i8QUVTJcd9bBYl/YXMU/26LXtiI5UYLFNpJVfKT0VLbL8+iur6aHTZj8Hy/NnqNWXYC9uVlPuw
1VAyCKucH23WH/nHlLendkq1hjqbMYfIb3Gq4VQVziTJvOrk8qwxzkNFYvOh6RHHXXzoO4FZWfoR
1ELjUokiM/3Cu6zDBYYtjhbf7tUOkL/EEj5ybFp+2rGo3OCEEfYxiHWK7nDaC/KziuhcvfMx4MKA
A1edONLgWD0xYWrIRM28uToLCgJNpUZUaie8a8Y+CQoHP4fbuV/K1CJmGjBn+UXRy/NeM7sLeoGA
DZi9/ZvP/1i1oPND2ju0AsyjJRSUm9TsG7ViJP28OXw8PAme385aObycYQAddDI3zsUUAh++Ufhm
VE+Vb+1Ah95uUIn/hp8W3Q1cWgNauJ2B1wcGyjwwZg7xAx7kRJW+sHcN40tTY/+VpZlFIOLpcHxF
UCbshnpxs2GN5MdPi1qGDwRJx5bjj027KkLMrhfmkcSTdChbaaQn6fSFo38wkzIm3xFXZWdLjRS9
UnBvviDJU2kpBDfzf3oF5ienHO/jPD7aTt0pXm/0UvXuktJHaOt8xXU3+3VUGCtsWG0mNPAmHOz9
z0Mq5DkIt25wlRwcOu9mhsBp16OgmyiYI+BlFi1Q/dW41VxKLoW0tPWBt8rZeHPeUHG+eLK2f4EM
loiLRd6s8CVN1SzdZnaGrFtwW6+GLjfXcRve+sAZ3dp6Aw9lAVInolujwXkOFkSTvp9qHqpM762J
60jOihcaNas7z3R/4HX98MS9E4IzYs3LxWdZWfoEgYnyab07nKvGH1UbFo8jFaH0dLveLOTARtqd
ILwfYPmEcH0OBr5gwV9fWktrkC46+THpaRK2cpOGe9sinLGj83F/2ZddqIqFzGtv6fzYFEUu5uSa
fBUb8B6u81lpqNumcirScYCveCTz5jGuk7Kx2Vi/PC7mfTGxoG1hBdoy0R8F+Bdif1YSNbxvx0ee
kZZV+DPQTsclp45kEwiI0g1NJzWtsMxSiHMwA3/KSh/NQr1VuJLwbm/BIfF8SocjpAdLwk+YZuJi
cdeZbyTs/Qndgo0A3p4fJRBzWQODoeBA5qaen19c4Ngwx5Sup7/HtMY4FYSeyTghYAIRqN/T8ZxR
fBhOxqDlYb481CZ2KZJQxq7eR0QTzzvnYt5OxwStR5tdDvQ+lJ53Lp05U8yrsR8VMN7LnCUso7e4
nsY9TNA53n1PEv5ZdHvsQ1Wn0DP04LoZM0qAmG3/cRrao0/+paxTznTOAe4RyJ++wHkEzMGtTStn
O5NNm0i5tgw/yw0ddRdEcascE8aNOLL5QvHLVmxROjLj1mKOcEmLCap1yMnFo/XZg2TIbY294E/A
l8sghBqtcqEDR8srsKY5jIXo5+dR5wMIP1EzsAc7su06UzmS3j/+W6dxltIXSo44NY0GmpNAmBAh
M8pOJOud5G/T9A5ey1e8cXgzTshPSRPsLw5XTHfzDORC6UTcmE1sHz7PMMwS5LHb3DZinWkRAhtN
C+9K19R4tlDOxtMempqK24mwGV52blpkJfUVLs0QnjzKcdRaOsc2cg5qbeByRt4tDjkHiIkSqHQn
mG24U1sSWufqLW7o0pNzb81AjbH+Ihazg7OFb6OXHfZukKQ8bGRVLMkcTClNNWcXKlRTyu7kZYxw
sWAfvvaxaDyaO82+nA/ULGSPFO0Z7/IzcGJEwRCDgH0strn8xDeG9aMR80mwwPFZmAhgDdeAhU9h
4+IZBWZiDGokloFQyh7XxtorT8hwGpPu9t0DnQKx4jyMtnCMA7bHGx09W/F7w8R0F43l00yUa8Ze
8SGOf9cZpfJSw23kuzgvDIMoZuHLR5DZgBq/ZZDY4sQlxSuY1LsEl4CJSNiNJC/cgDJiM5+uOr/v
XMHuGxa2E1aM5wk0XVCej6AHV0VYjmq7DYBEvQ9zsKQZqPOX9ibB9aofbjtJwjw1bCejTmR3wGDD
Fcjjz6O9YRl9cQ7Wfl+cpQFrqwdOwLZTfHdWWBZok7Ov95L1HLtleOPlzU3UwVusVsk0YdCGbLJF
H2JdPdV97+tm6E4ZAmR35slAvXQ+UmzrRR9yBWI6kjMxj7UWT3aaKmG0gc8scjMjfWeZqEcnp02O
gfYmG3cfMSMtMabY4rQzRkZxA5urhkydvuauthR/2saZYMhnnH/CtnbnmgWmRqRU3ZgMLtwtoDrx
7bT33lFyRDCVAwRvAdBFHdyN02wuhEGOa2AlMeKZYIvQUiehyvEE3Qd0kbuSMcELFj0htA7yZh8Z
zOJIO/BGVSPwXOSnVr5adb0Oo7Gx7hhVtCMfORQpByzgXhDXLEwfBtoh9nRYWJZHEWrKGySt4ixP
OARcbpkqhFhiIq+gaB3j3ODP/UQvKMduARd814Ssv9MQZNHoxJLN/Re5TcFgXt5DWEEUeYMjKJWV
ZyHM8Uv4ybdyJE6GQJzoGq2xN1+1JLQeyABI4pXJ3vjEtgn5iEfX2KSgg/FfelLxdaG0tw+zPsWA
wsalC7tH7kkAMsPbTfhRVf3LRU86ApatTfhY60RvBKH5FG7ARqtmvlk4mjp8RXDQvhcGvEc+2AjL
8bK95/TCzhYoFE3WECRgDVp6l+mNC44t57sd1sJKhLhsUEOUAIpmrAKMm58jiI7VV+WcS4ETRgKG
+zYO2rKmuLXttgV6T1jM5us9rppjHpnQh8BQLYK+q8FDZ7yKaUoOWsYrbyw+M4X1SrWz7r/LUPxI
I/F9Ux1KIfm/Bpc3KBpjH7VOB2muN/OZslW97bvPPk4ubPgIKXnXZCjEn8bsZmkm/im/stqoOoil
NWLfRgHezUcU/WZffR5ZfUMhb0JhDYCEi/Hrbae3Zo4dnfUDaqQabecFWlMKI0Y2TNDlEPynxpUc
loSbP2wrRi1F0YVsxsLfmQmoitUofyduHF1sEMXPvIiPlpBDS6VT4TLLa/5GfsyF9qClb0gTGLzm
fDG9iMPEZxR3NLHGDjLACaMajjC+1l4iontvNscfV/mWEh4X03BIJ06MExjSnFocR5WWoTmhr+GA
Nn3YhIFOhzQMjeKyiDLjzJUhUH3GZ7+WBTklaj7dFk9HQxKO2EddewyGCB1kiy8rNz9pV6Anwzh9
kOTb3Sv6po77fA4wqVR9IbOR42enFZj9pWIqfqJasJ8iOvm6G4KQQr5M6NJcor2IiW0aUUIUSMr/
fRL1OTKfzP0cUqHf1Aim6tScVQa5nKQiVsdvnogFHm/ANSfLjLSDtXa/FlVDmISbq4iJ0o1HqltX
337IoydyFAMQJC1SiE842w25u2Iwz+qqh1I8v4dqVodHokmbco8HMt6kuhDPtetpLFMPzP1SQXlt
6m1gDbmccjRmFKgpp/Nvjupvchki1mlyKC+6vC8+cpL3I29pNmnVX2k2rpuE3qpi7v2jZmp1MthM
4x1i387pa58wa/gPH430hmFzSpioZOup1pSlyv/7BafVUiaUntU2PXEgov5ez8tLqzoYKJUbla+1
CYFlI1Gul3RFab8s9KaHMgJ+9hEBWAmvHxwqps562lCdHVV5v0jd8c2kwEQorVGBF94Ya1XRyc0e
7X1vyhHPP4HUmurj4yM65POOUg5NvsLCSfJicDMloDkXHJLzOy2k5jFzpwTNb8kTTtM/HYPNmlq4
nf/9/wtrBohoowksZ/FZZvVCMbwAcFeOPwFGVSN+jkYy+1BciFiGjfn4wdG6iII2dxbMbxBj+27E
/T90hWXWxR0vVE93SqnixW3Nwrb0j0IlPKjZmHggDaa3oiT8ui+YB47qyzPswcaBmA1SlqOo45yW
dJOGZskv2HehqLdgxVvV18VsCVuG+eFmve6uezTVja4VIw01cLJvhmeo9vyLBzu+1t7kkEn2zT7D
xQeOlFSO42yF0MMxMJRNp/KXLV0rDPR+9P/Ob6mvRjjc5Ig3ogKweyvLbjBeQ3VGS4Dw+KFDYIyr
xbD3XDrL3V7vwpuXJidYJZ9ylCZtZpfYE12IEgMrFc0mcjXVWDa5KNezbEydH0QkxjokkmPWXIqi
HO4h7sCva9ndc1MLJDDM0nApA5aqcII2/dqPaFWr0Ty0XU8pXJ5u4oJX4Iztm+IEGAiQhiGz1+rg
pjOchnbvmp89NCKOkdS0tq1Uv5TDLrsykzHsxkQVacR10TQzfO9peZAPVxEatDfE36bYd1GVYF+z
5dJM+cQzP8VWtsdw43m7+Bs4qLutsqMG0w2SN5a8NZXRp8ysYHQM+NnxgTDtAE3n7hhsN17pUHUA
scwD0yRbfXejX+7cV1BWaIgxSqzNwoSxHzLJL85OkdRfQgp+jhXeqZIUJJADXFiShqUS3DByexeB
C81IzwFtiPC/W/7Udd8i1pyMUoPCNkspdGfEJIXmPAw5WUTR3WNJW6gr11+I/xtDJMQjMJ4+QqMZ
7S5lhph2gWRuarA+WZbithjwWIHRueT9P0mFkXOUTfvuZdGbnQuXn2pU8o6HZGJtGXIxS6i8YNJm
hR7qgyCYkiTJ/pbEvvGSXiY4lFodjx0CV3/YTriNZFCbGr2K0EkjazFCBipYwy49vp+f9mU2M8ff
NdqpBu4GbFuJgoywXIcjU32yjQCZujpvJx8QgI9MDX3SrTX0D3s2NOBgxnNAn+c3l4xoYuUaDeyl
etE87skY8IQq9viAmShCvTHAb13TtWFe0OEmXTNVoNdXbXDnLG2yKQTy6XQ/iNS/A6BnubeI7wIO
bZ/YNsjpqaqcgT8D/U17+0W8b8fdTdFsJoyG7RqfR5GfCiYujZURmDvG7dZ85dKKJjjLX9rKJyhn
3RSTOvJCFj4n+q8sLmMo7gY1CGEqFS/zEySj8wzAbz0kkhb/fCiHvb7I7Ml2Kgxn8ZxYW2x/OkKQ
SGWGIsDpbdwqwjP5kvWaMdNUlVA8xE1r1WgnkInP9uDeK3wCy9e9IaqTR8IqPiQHmg3Ry0RlU6+B
565dh2IPLciUElFLjA8OJWKV+qg5EJ/mKjoz/yGIxsrZWZDfW/Ugm0b0HYWPmRhjsSR7Tz5UVJJ0
8bDBxoxwz19z6dZUQj5vzqIzuHUWj0obh5DAxprffPxhRgC1vM4gkuE0K+GjDEhqc9wbB/ub0R7a
m9byC87U0/CPI97WRsHJrhAMCwlqQ5k00Naib0d923YSOI+exAChNxyDRUxMfUcP6MRP9oYKYZbG
uB0pZTKAn/Z/UZk9nMPm/msGlptj91/D/WbUNTHTl2N2aH5bzXqxfbY/SDImDeQdakOlQAJVNhDj
DTeXTZZymxhCO5pGlmdKo09J9Z95eK/iK7/GcMpCG4TOqdQ1ZCo8LYr/qQaYi/zGVG6PJIpXgFYy
FmdSFq2Uz7dYwwOmf/IdKrPm87uhFyGNkXK4KahZbQVtQ1DRSI1lFnTtAUAouhuGPR4dnp6FdHkS
CTRX7KzbaPFocu9iFcVLjUPGWWOYnPbsxq+qhTC+C08Z8iWrXPs8dnjjKkO5tzx+d1/VjXtq5Zli
dLI9n7mR+Snl8GtF6BEqZxrfly5+Gfm8sVES3OxObaZ2Ik9Bp/TKe6NKYW1dIUSqv9UXoWlIW7Ya
YBO1VUYQcO6y2GfxDzXvRDkHaBjfe2XhNVdepiATT7agrDZOZ1XkcBkC2Y5Eq3Jy/D6VtKwRkPt8
gy4zw4RYjEJcWFcLoyJSjNbkZAf4DXKFeebphBzbIbIARImWDJVJlOB1jCF5l+Kol0icnjZqJfY3
2S9DFC5JTew9Fo6XMFrG78yvbPr+H6VehAINrq2oIAFK9015aJ4SeXcuM8u+5g+Ya9FY0066a2gg
KNciDqSZrf81tXrSvbJfn2gcLhAMTFdsygUHkpKSSIu3Ffs8ylaeK0LXeovftYVq3nUieAzNGWW5
rmTu2YHq+AGToN1WBfT8zq4suls1be7aC+6C38d71OmiMQexSLz76Y6o6hiUEd8j/VFApoVyzqPv
tkVfumS8HeV2MTE9hB5TSYYtVXUlZnLWjVhJFD997W01916gNOB5iI/lyTk3c5B6Aiu+GaNnsKt2
hvnBE5UISvgnRECuoiz4mRMj4pmfHOi4/McJ4zCHEqA28oJXVwz1t4NUQq0R4pr1jdN4XblGADRH
irWuuel/hGFmp7piMso7f5fl5lq2A71uGEMpDso8vAWmRORI93Y4eqcbSeyoKDqdXWAqdUdCQf1M
VOnfs2fOAKBiqpg9qX5RqDQ58UA5PeBAqVDMJPvRneCjmMeqH3/N32UGrQCR4gWG5Qf9U4WSWcjh
VHoiEbnbnClcwdk18wuu/QKRd1m9H6K7utt4y75Zutyj0fwzhmnPedaoZRWqEjqc+QKsEgYiEGdE
XAIHOB2U7HeKYR0JAzdwLxQ0EPECf+G9pQ3VMXSGH8crw68KcLWCRMVk9iJ+C585Yx2zx0B0ctHn
mQiQm4PtGQZIRPvFnXq8YnymB4D53RepZTfPD0Vrz+HYDC9eVslO+qvNMthgdirmhWDwUNngy/0V
AVb5+ltoutiaFhuav+YjU0aZvfPgNMELwl9nkrcAEoBf+9IwkGAH5u6vetcyNGOWi7mpHeNXwaIo
zZQbAYNQaum8LPnvgVmY4lwC5oATyNpve/nPOUWSw3iIkCTueVUEXGB8Kebq1PYofyP5FU7CEJUw
vesnoH7CS6SWdSSAxyybp5SGgT4WbEV4j3DP10pBwh3dVfuYRsedzlmkqqG8/5jixO/6CrP1uFnH
85pTBnxNV0XBsoMcPkzYtEHE9HXvUCatgPtbzpjM6+mGQmWn+1OsuWxRSdp8PCCapc2nJ8Esw3Wm
i9XA/rlBKboL48Uoo+UJlteU9zMhj9zR40mqGcI02zRfNzqJSGf4NRakY0/hefMTeSUZ1oS+jGjF
8dNVaSePcLsZBAlncw1HEllwgUlgmX3BF0MLd5snXZxbvopbmxgwUQr/7c23ttfnDJvfspjpueTC
tQ4WLSjsw1ealb1AdlhXa7DcyjNHuo1Ba6ezNSCse1pczy1IOtbSoJTeo2+TIw8cKjPbGL8GR/CQ
ziITAMTW+TBnss+9QLX47r5o5fOBTH7nPxMNbNMlt+KFDLkKgMRaC+qRvJEzcUimRXudTBNJJ4iK
S0X++wpbBQJ1go06vWzpIqUJgfDTCY5fsVIWyT332PQ8Kz+BZiAJ05L0F7X8UXM1L2sMmq6bLz3G
Uj3xfImvDnRc+oe0SKtoaADsvpen/op59t8PrAvx/o2OaHe/EqRa/1Q4iKNIYMZQQU4Fxsl9kE77
EeP5gWBrEEZk8OvmmeOD6e9HsE2Rer5xKmKr7xqC6h2OJdDvqoCEZyqyIDwT4oEBAqJ2tDZR5WgD
wFwlc1F8kH0x8pLhnHfGWucZGsUMnYxXpyOisyYIwOccYN3vtyY7vYXauo2g0qouPEIqNUbuV1eU
2/ZUbkZXTN02kN523ULK1XpvxDkoO7eAJ88JNIBUZBm1wxKoN7xYPYZfvt7hew9BhRE7URZmBt+e
g5TDeVomyeq1Phfln3VInAc/wHvCo1eGZv2o2auPWq8n3Yt8LyVByHErBQQNWimA+MEKP5iaoZ+s
dX13I4/FNtQoM4jGr8lEMLqevp0jsiXYcWqFb8A8d/ewDF9gYivTIyv3WUqDQbwcyYbOSRdlMXrj
w2NSHCTwsYZ118lbGeyxVcGFuxAW9f2hdiJ9zYhqWd2FR2WT2aPpOUfUDYph0Oljv8iDeHCa+Xm4
0Hb+zuXGeRI0LSOROKDGelHYQhXGnv4olB3WmL3lHNtboSAq8wTFYXFqg2U/Qhe4RN4KP7pbZP7O
xz4bql3jaxKcv0T63Ct2k2T5P7n2qKDE2chMGy3C/MHQNnY6vpjmZ8kX0fgeDi9OGdkCVPZMMaDD
BIuZzSUhW/404IFEYp8ttjXZzyH+/t89aMLueUAaQjxZmpYlBupvXRL3emsL2qKau1joFKKPF4NS
p5q1q766W31MdYXVIN/9xkNk4UgyBrKr0kHsE1c6lw91m5hUnVG/EpvJUxDMuXpXEGns/UK3abF5
ZhazVdLOJFDdB8R/8zz+7fa9Q0vAjqOQDJUZKZGX7K5uLHVwt7R+7DxeAE3M2ZioZ46ySc/4uP0G
NfM08KEFnlMMRzZ+izS+NjplhGef22LDc0VvmGqLjw2OJl6wlVJM+yD+g/VrlFCGFUSoD1He2Z2h
eZGCcyvo56GWyCQMPm1XY17zPzieID12TWof1ueYJUcwwa2Juk6thyrR4IReFRnhLn8trwHDXbcH
s+dpjdwcneRTpSPhlYZTDV9pyQlosCgEiilfitmfA2wS3k2kvJJF1Pw7Hy7L9FW4bazHpu1gwqHt
8G1kWW0n3VU518rBLz0uDFyV4lYmmMVbR7k9nKNyrv3GVjzr5dFw5tHUoI1ABLPQQ0+bpoCAeZAm
HmM6PeLV5GcLWO5Msx2gB/vJ0ChaL3emqt3CqFZNgk4QEJGs8HVnla4zpgl4lQY3vMmOWT8XYj8X
5Js9ZvWCZTPmI50nvpuLNVN0SnpUaNbCvXD+nnHQ8BlWicL2qa0sPbiE7tw+pVAw0MH7K/REniBC
12V7zj3hV0o8Q9uYadxnFgQq/JKuYwrVxrsQKPiAAgn+ZmuoxTb3gV7YyuesR2grPA93EiwuHOOS
fjPn8V1wSPeuJgFmqk1KhENeWVEHaUvEgfiCZnjyAmlnZxPYIsvWTJ9btAP/Tmt5WXxqBBuumHRM
mNQuDr+KwAASLsrltyyavSyUYw0B9qgaMtwYe89tVxQ8u6wZkl3K6wefpBbgTE6/u22gOJ3wlNKO
+oVdTnOatNZOcfDwswXQt4kqc7MwVoA6sztlA8Nyh3nDjSHwAg9DblYdYke5CL9NU8M2/v507di5
U+aE/UqaquSuVJVy9SfGxfJ65z2lkF0Ol9uCP3Q+8yOiTAQkFn3LdRigdJV/5TpIR/uJSyH5EQsD
L7DGc0N5bBf19jh9P8zBtkqiv5CkxgRp2t9N755Dm6xvyegNcYOeG1MDzHfRGrrnXyqal8cIU6Dc
rH1GZy0cI531Um3t2+XHcVb4ZtyHgd/++R9N0YZIbt5NsbzkRpLxWTtjYNDkP4K27VUAqSwieUiI
t8JcgFt/fkke1amysWRj78/2nP61+4zq/Eo2RRz6zEOodb/G+9bjb5ACtmkNfPBMyLIQj+kxxMmQ
8Qfq2S0UGGmBT5epheA7YpC2SKe86bMTVCLt4UvVcR4Dizdb+5Pa8Pcmpo3FLk48KOoyN6e8DHn0
No5H3EdCReRlETNB5ArGmMiMKDoF7/db2xFtoRMO/N+p2s45HNsO4tqIxuPb3+QGCzOal5Zn8g1R
tJ0+ajGvskQLo3frla6ft4VRVL5ijyvdAqtAue41L8kdUZFb+rkFgo0+kURH/joYWCMcVvNbXJgw
jqgjIeCHOvcEHDSjqN6K69sJlkoXMVGsPqJyHGkgjO3Gy+srj5uIsV8czhpi4EX8fX1mtPfH27GS
nAu2VSDDwkNzIHmPSn8xL7i8K/OtJvJpsaIiuZJwMCL4eUbh7yQnAZB+Z61I+eJyhXX8h9TNbinM
gR+0dfZVgFfmt64YUAxPql/aTyqMVg4ykYnHNmdbFWM/2no8rqFmE1waTtGrXFZCD2wVd86iKVF3
2PNqrwIvnV7v44/yIb1Q0ron8y61uMVysplDchYF/69kbeCLnRwjehg5k0tTmD2LlSMPjiv7SsMu
kW19gEt6r9LHJTziktfrw3fCmkRnUwqnd4bBDa5IdZr/kXupwcow1LEz1yqow/vzARhICB1YdsG3
hwT6SRsuoVR0gv2RyF9C2Tuqz3uh2+ChDWRWvtd58TGKvxEFq707/xZ4NxpwVJ2DG0qNXz7wG/W/
PB2z93/zQ1NUh3m1OxzPC4qddGZq0mY1ig3zHE0ikG7ctF3J7byT7D6+xr1bng5Q09HNmsggq2CJ
QN6OZIuss2aZ8rLmVSkX4yKJoWZ9fLaFeV04sLZI/zadkTs7bccfjcWe4k6AVXveL7deOr7WWQWJ
YZbV0qvfSLx4zIdqTr9VE+iS0xbMiuYRQa2RZQiIR3LVNyX5DbCDKpLaZVrPHE+0a2J+ZE/90IVF
9HzyjdqRjw44vJuPDYc2sdFvvY2YASJBpuaIELDi4a/pzrg3bUAcWtRWkTfvLnWQVYd+5d8Gfadg
QMdPI7EBOcaeuG4l/1X1W55M0IG8PJ42lzlpz94v1E0Gfsrn0i2eJrPhsidXlFwyt06GNIDhFmPp
pl+qeBJDuc1Td7zB9svj0Wk125Svai8KHUiWFa94EJFVFJ31os6sTOxZh3ZJJguVLVCldBx7UpRy
3HGhhVb+i6QDG3m2me9vHJth5PTMgS/AANHmgRQOpqIBAXENjJkyj9eBYfdO2RI5t2zVUpd5rwuh
J5pRwLr1bBTCVLiXXwlW7LRwEugrAD3WCNJbHFlEB5ACOvpw6x0uWMrjR1i9cF8C2omurDZd+Yfg
1xYoNIdDzkGF3Oq+2zfVTyZb3lTDkdVVZ1iJDH1BJSh9d7RKTmzE0huiBdS+gS1Z5Mc0+RB7MAiy
ujuU6kQDE2YJv2gyx1SrEH6hng/IUxEsiXDS2frPIo3uq+XgNSZ8M9h5eXhVTrb11gsp3f2N71n0
fWj7Wv5Ehx8iABfunrH79JUq8Etg8vDGB3rteOPWTjXFWwQd6NFfOgZFIGNkO0HFaET0hSSOE4iz
q87h6n3A+Q5DsfZdxXeZw+dW1s7bPhVjCBVNV2eISHB0MaQBDn7ucLB3LGvIBlEKPzVEUxe6kj4F
Xhvj9aDk6jmfGW7z+qZ1AWur12QWEJt1+Buzc+/U3bZ+YBuNwlJlvBvKATfRwEBDH0ecD9GnbZJ0
4f7pxJyETUOEqxn/HfuRD9LgL7LopSEWNAgxZ8MNh/GdihPM+AHfjujtrQ/shHNmqNdpkdw5bpSv
Fqjioyc60tLf47BGB15DgTPgBYGDU4ObSSb3asuXN1rNeByidflQXfbGhlaAk+lRAEAoB/sD+Xlq
9t4/qvdAG6NIkC+WUEkKGS1f47mi/CySuu0RMldnYI0s1yemuGZ92Pab+31b44cDtwN9QPr5ozLK
PGME8nqw3rfyvt4kLSVWgk0aDBVQ2b2y/TQAem1Wg5m3FnwnvL0FjqssS76rJQf7r+gJL3t4CKaL
Ox2aZ3e+sf0Rs3vz6VSGDwFK17PJE9wxWIab+fFYBeYCN0+IST31rhmufs9AVF7ZqZD9agnWqbEy
aurbFOiLo0H0dOJjDOjIVBaRiRV6cemVRRF7YMxM0rP1jh9gR+cOHNEH9iDpS1xRU2iLiVWTShu9
KNCfQNre/dUkueYyCKyJLjVh44yFD4Jqvg0rVTHfaL52p/ia/fNQvNgr4phG9O6eMOlNyHjzcTFZ
LcgKCsVEC7VWaMnvdRPpU7A/rfpSEQkh21sCXYLVh/uJ7qRyrHyas4Rw+GH0YDUpFrphmUDxnMGu
F557tevaB5vl6LW5PMwI6Q/yH/Tim4QSRzHQqxwwYdcUsblWbHfcRVc8UU8+JFUI+sP6mB2et14u
xbdIUohk5YPyAAl5AUFqbPbXZMT4/4OsmRMssbxvTnnvnZvJxhdhI7M8R56IvxTO9o5PXNytzkRU
QDq8J8yKu8jjMNwarlEDhSge8pXaeAsqjL4mT0A/klB0I71rplb7DzmybDWYmEcM7PBqI3d2KiOi
vgbszKYmxUYXH1sfwFPB8HgRB2gZL0iIVxXKn/TRASMXncbhyvdL7CABESpPIHmS2Rh13g2teQUS
K0ZBTboG1y5Uu45Z0s5mioX6eOx8881Tls7YH8p4LovVqI20Oq0WkRm7+q5kTh0JNMFZkYozXuQ4
sL1UU/c4kdLs6l4v/gCyPjXPGXTRnOp+MxCnv74vdM+x1N8UpxJbKNkYBauqXU0qkeF28ymvhEu5
+6/6KkkLknzMVKthkDhZFLoOKpro2BVWE1xG8UiK6b9wxBKksYWGRnUU9aI3Tg81NHSc06NC1uyV
iqE3oYJFoe0ACnPt3uhaqPKnehjrD/iJca8GOs5vA3P6r0h99Bf0h1Cf4gDXuEQzEs6azcwd6yB3
FNuX8AAH80wjpJcDmgLDAAT4omKgnK3ki9/XhYSOsbGe0txARDQ8oeu3m55h63urZet7Pa1w9dU9
0pcBEEg4zOoy3Tkhc2r71ohfajqD/VrPpPSVDAtTEIz7G04JmkKCVVIYFVtFdBDr7EXldqPXGWZZ
AhXTgw5fBHHzc6obTCkBAIpr9INVKL9K5UOad2O7gTwXsPKL4vsTSoejSXm9wcrqMImi54vClVsI
166u0RkQ2OV1qv0FZrd+VuhteNfZTs207uzD5d22XSnJ6uzn772/kme3vgDgZHgKf3zECY0jmD3R
4ktbzIKB4i9zZQQI+ox3aAyJf7eVYNNUNMMOCOvNXRaIxO3MZF2bFwfyE0sDinkjAtEZVTOstH5F
hI2nTNzyQj9pvuysVEIkuBY/WSUkEQxoSHllfkY1NtNeKWW99ZcK+UDxOns5nJyg1PVAXetCgmC3
8PSCeBTANZn2Ttn+byEz2dt7cMViWOE08QzUzjumO0NMYp4wWjmaquNsfuGWZX1wZ+sMpM3fn2jH
YZAQrB+NPAvWOtkFc4+IerBcheOXVIWknTUBNEf8YQ8Y2lFBizrNFbLiFc/MzJiY5cY2Ts49mL7K
Gf8Y1IqsnT4CpjVNE0NJji7GZdnnYpbAXx6vMnxL/t3WAZqLuNg2pAJ2fSi2qCt+PwcPuzfRj/pf
oBLBv92ufwl2V+oreXUMrPHiFa06wheM3ErT+mpKtO3mlejl4mEzMF21jbNOX0TySa236yCLdc41
K9leICsYjrG+wFZwvQAy2RSxQ1zXu+pIkKj47x+Sp0576ChR0TLrKce7Qa2PKJlBKKGpqgVE1+J4
I+S4ScU1YHNUUDp/RKn6c13XqDa0m9J+xGBLoaJvSpSv99llaYdX2Y2xtg0VCab+O2HxcQdm/D0p
ZePB0sBFVJ6Vd3+ZyruVs3kBj9DvPNdF68/zEBtXfqGG+NmappEOCpPIV3515SrlXCPFtnz0M8rf
rDw/4By2csvgZzj2+PsFLB12LpMdTNYZcpePi+/7gQT8HzrFTj1i//3TLnTjnwVGRYSn17juYQ8P
5xjQHXxfnxH6FdHQtu9HLbKcF27fS0hkABDAbsPG3pRs2/Ji6jcudrm7nunGyp6trL9B83mDWPix
FS1wz907SJdyWXpGK8HATM/pdHDs+xu1SriylcqDw23kbWGxlCqAOI7RataoK3clKDhqLBd9nDZ0
Eu6EJ//1lhRMCylx0sFRydx2kVQu1uPNrLvHEQOpaOOPDR1fsYsPCMYvsmRl1c1HxhLPo2btKAfE
J+9z0zqDqYR3pdDCNncZyvEFgwGsgHCBc/vc+l4ibDfTUOAIRQNPE+uEZd4Utrxv+rDZD8kNaZvA
4Ppgq9kVQONTrmSuOJlMb7mN5YzX9SSFW0XuTfe1B0K/Pd1R3WlXh6n8kK02VnaOQPfs36/CgACw
19Zx4RouBU/zM6DAQtZhWLJcUu2Tzn/TDUdskB5ZSJnlTh8Gs/bkg/YQNOnLvXT4pWP3SVxrHdOH
LDE2elusQOW85makarAZbI3M3UJvgBFWF/OMKfZdyf9ELu9764CiXqZR2PDRJev3SXbCgUfXDa+c
+DhjZ5PeqC2HnZxLi0zsbrt7kVbeUKq+PdSW4XXiwPscT77J9kwmsXghqO5RzMZrNZdGbXuIiNuA
qG6R4X8ulY4tfZjCvZTJw3y/fGtYksxpakObE3Glgvmh9T8Ir0D/qZvrn1exWsCnP02FTfSWWdOb
jw99diWhdJZ+7Pq5tCJxTrPWnGbcDQqkyb4XsWNPygxK3Uekg85cjEDV17pQYoGowCLbgJMMYErh
uVbXHy/9RfQZ7P91RYZCIXLctmakWrYYD6bU7Wh2yWRCpEbAa9FAimwWMpc+9pvSQAEckQuCbN9F
mN9w7nYopoG9g0WtaS8uGJXBU92fSnLs2mVi6ouGDy0teT0mJwakEivNcOGU5MgwhGhgkyPENlQU
Eh/sX6mdhD0db+IkVwn35vFn2a1wxgm5ssEi5N+2hPXtXYe5iT6T84oOcmavgGSQle4y9dukhqty
Xg9luyhoNtHUfoewT54VyS5nAej55TjlzjvVIGBWTI9Iyq+1kgeqDH4BPinpBB1iuAgS+3pyefem
Nw3vVNopFrv74QGs8+ulhWCIAotH/GekAWTtWx0Jr8MwEfXCRfvWFT5M9dDaD1GOkJipaFY1iE8E
UBuihl5tU+3dZMg/Q7YDYRPycPzVvMk66Z9xb+XvmF5MSy8OXo4j9kgE2zIZVd+6k11M+a7M/3O+
FqFE4WDqBRvUolw/IMnCm2rYShuBCeyv1SEdVz4fwPa6GusosTWHFt86v64DHqf5mS/KjEmGl8J+
Uk9Yo/80UE0FX9Z/gCsvK3tCbWlY6RY4cXnTEVGMWWTaexjsRJXL48iYrV7uqeAncozVOr80w65a
A2dgTVh2j+ZL5k9e4/iISHy4o2UY55OxD8TRe32g25m0qWG45hfLCftP4O3c3pQjqHHF62OdjCzH
aGKwC7H4msPFtMwiXQrbLQkrWsiE0c5nMQEZiaE01+U+ocI3hjHaPXyoM0pI/R/LIx4S0Y3m0MvU
hjN+q2YYjDHw0jHOwWpgQJItY/cCjt6WWsX5lILboPl5c7crel8I72CB3VSW8lZb6pP0/5NnwXv2
1qFDOD8QVN5K8Vp+RLE8J3U5eRg6tX/niX/0GZKyUher4EemI9T4sk9IKutH30DIxxrRl28I5lSK
46+cd2dLqGf17220cv3QH6Df0Bp4NUUY+pfonAy8WTW36U1IrzUfZKoLJLWWrhkL2anzMInsCZXa
hKzr2xX0FrqbB7xySpCuuXzx4GJ8KuiYxQxZQzfmKpSfRZiNgFO4ZXORv8XMHokwNusYhqUdUy5v
IP5C8Vz12PMm84I+onr1D9ds47xB2Y0cCY2nHVhoTLzQZ6Fiw0Wju9Lg7FGSCxq0QSUsjgT+8IgN
T+wCcMN2OHw/8payM3h17CMoElKbkv507/ezD/x6E5bocyK2xrWRchpU5JgNFsbc9L1HBbBnGhMb
4SNK97xjlPRvTkR5VrR+gZiER6wOAGdcauzpWKwFr2mtq8U48dnILA7gIvAPux9NZJSSPfYAf0ON
q5AM8dClOJGaOhPrt6sfc5SJOgLZB2ggVxIEztFIw+mhNRk4W70yEtpu6ic4rqSEVVJm3+nGx5X5
fdHzd5RifcxRE9qgMlh4Q5V1yJ6s9H8tm8/ursFvM/dOSyFNNsBB++yJQ2lseGtIo7De8MAU6mZb
zRH6RZ6JOFh8GOAsI5GiNBEkKeT+N2eTSa0UtyXttNrRGtKvloxHm5b6WByXE1lPB7C6wjI+JW9Y
1CAN8DTWO+LwyFyRo2a7hyY3Ji0VkKrr1/5Hw1cMrsCygxdVXEqDLQ3e6gulJuy51mvqfMOBviF5
MewmIJx0sWom4W7kmsW43E3jRgOX3kD7fD9Uml6PgKVy1GrRJb0v9Atf+78W8nT0inoX7naxqJZn
FJt9sOhls2m5Yoga2lSYjALZkoPJchiX+LY0196Qy7Qu8u8vucJbaZodoAz0bky/LjoGJ2/u1Tfy
vTuYPkpoYuOlZPQUuSyTA2KvtcrqOwjucgZtR+jjjM58CFZInzYRM1q10X2IUT9Ev4QMvvd1qBNH
kFhzyzrj0wfOjdileLHTXj5IioywAsVYrD2abYVIoIaa9x850grQAa8n75C7ktPC5yScCapPlvkh
My096riW3W11BdfXqC7WW55ViZ0rUXQOc06mIe4xqSFRazgitnKZ2qx6o0QMzzg4kWistnQ/DUbv
X8D7XMu7z8jY8JZ/VvxjOvkgQwEF6uCAZEh5KK3VqLcVGRpy2y0yPQ4biWxrt/w2BjKCUrERTfFw
jEuRfgkQIqdktc1ux1eqIKx8suM/ncsiR7VDHmEQgz7FlmuhwQApsF+3YHaZkNLz8awnDV0aCxoh
C3V7xZgK9oyGrBS5vPrinJbmzTLubIhZLpZq8+7cbjXn1hIUAQ5sdVpB/fYeLp4Hpr9oK+KiYpIi
UlTrmw7a4RWcoc1YFbeQSMmNGO7LYzs13L+LhcCcjij4O4ziZB4MIBXOZSTQBAMZWswFR4C0cFHW
AaqOrt5qNowOZHpdSEMmt+yT0ciY52TIIWsP6fpUdmK6Xz1SUo8RbxEXO4yLJNaZsN56uBH+mxVn
iigS8J0th7OTuuOHgUfj3oHmPynk6IUSwwQJ8NFKQ1A1UiKbF1FtZjNm3vc3MgSjcwdiJeMwTqlJ
FFko59H+JRUunSAoUfidM3kQtxhloSXn9qk/7YWlBCGfniVDWwQ3+odS7aaExgWqHXVH3Xy5horl
rmq5/iHagj1/GB0Sr0V/zsSwPpq8eh+W4MbJxHmN8mJ36+rC6MS2SZqT/YlnuH2vLPz2r0a479L1
UW0SZty2KCj4F8w0fU/XSf/cBhsIs02+4M9LFQPInz2bNHP3x/vY++IV9VSGi26C45kEz9OC4wJf
fKJubyUezjgPuNYDs05uuEVgvseN+QOE1T7zkYP2L/p2D7Qr4Wi+4d4XYJFhfu4SklK2mFEnmTN+
VQRXmpIRMnYdr5PKhAhZQOodKH9ravu3uDgd//MlbA8Io+3rgSOp0H8mcYlSpciHVbPYL4ZYF8yN
poaYorn/GFXuCHbAd1jcC415BAtgc3RqXrLkMWIrKucygYBjoL8VFIkW/h8k23AfjESgeHOkZ0GU
sKaVv2ShwWoEOaH8Sl9KBMxbvNrgOdgR4c83swGupzdk+Oj8tFv6hTf+YQ29x29LPnf/4LnJgwbn
j5ETtqoy+zkECdZVsf5KczYEO08JERNMhJulJmVtCcQQFZqOgEjM/Ai+nA48x/XLsmBH3bEhJ2GB
zU+guva0W6km8quFpM1p4l1ZZ3cJie+WQMWRN4UZISEBAAkaHHLHfJ3Du9kjNbl0PJZormCKZv7s
c9uH3aLS/vNzT35lPYaI0GWE8qPQ/irJB0+FNxyEPeZ/pC7bM1koZpPJZmDV09vAGKIlRHAIzFds
NuM0ceXzJ17gP2Eq+n6DcgL0kPcjm4klA4lIAAO1XHWtMGIt5NT+q99GiddrWoQ8SLBhsHCUNle9
TDCMfr5xbCNGmncfoOTcGzhVjf5MTqv9EdORMc/mgzjvixUYK+uvCGhuZbkgW4Sj8uZ97cr09BeQ
T9sJyWCwsOd5gzYEyeRmHCC3/iDkwLhcgNpskjUIKgBC8OiWN82UgRAEpAOCc5p0rWJQOaAwOt/v
DmvMNv8pvTRccxUviIclAU9es6XML1ErDli8DMKp3KggKHVtaYxy51hJuoUc33BtN+AO5FDY71tq
ZpDrAt/7BaLt7SkjO56BhSwh0sP/NbdYEX7VFW5y8n64RuHmQVcmCAlbZPKx2BNtKUmm9UnWKlBa
XZYsay3l48+0N33JCRftXBGO63kb9Kyi+fIgk6+BO1KBxQYYSYvMwj/YJAYFSe7+PpyW5K20oc1w
ijRm6KOuLg8hPMaqiokbJtXQOl64f44XmTIYSRvumKJLFD2I2k1taC+OxPRiH2aMO5izHHYk/4Gv
Sn1825WpsDocEedH9jw8foFNDRaIfylmOTziEmDzz+Zczwk7X2HUxODm4s8FC2wJOVzoQki38+4G
TZ7ixFLgsQtKeXhnAkbGjg63bd80SsK/nPYN3lPMi9EB1h90YZz+eHn2jDjU+dP+bC1aVkp47utU
PxACWBma7Wf9qysX7kssG8vj1yRh2AJvEmEwonG6k7CIrrXW9Nyh1LHbZW+IPXOq6NGdhvhyQIQ2
y5DQmqOdNX5JDwsxiFthAxfcZpBjZINb72Upx2uoB8qfpLfmrDDBXDy+hteHtsLgENMtm8dzqXjr
tR9GLmymo0nnwj7HqMYKw42PM62Oq/U5ueaALLBYi6eeUjdkjEsKxwwwrnRYqBfHwhuS2cz6M7Y7
lok55tBW9Ugw6q/mSNtb+i0qjv74YBzDhok/LRVAQScWRreLmgO9BcvhUzRwhLjMfwWg6owxcdiA
eR9FH/1btRq0WCglz5GDhpyjGecJ/PoxsQa+cnCjRRmzDxM3rwG/+vn95SJmGhSbWm9flOCdare+
HBN7qdRlwm8GahRadi58y7+z/PYaimFydlh6v25dHniMUttClj2Axxw7J29it9mLyYN4T2pzqGnm
x6uITreOmBZjzaeTLXnsPJrDDT8fPo6v+RjK8D/vmdW5w7WdKIKX89AF+HSJQSIkMuv7bW0t9vSE
efC5uRKMSPcpaIuJV1Q3tDYuI81/2vHIJrenZMN7ZqcJibV8KiwYxMpwo3BB9oZT7+bzWe8Gfda6
IH+uYA7ANR0n+QHHE6uHOTIaP8M9vj/Q9bJ8PSNnXaPQzMWwg9/IhiQXDklb0vobe4TZ7fxWkJGO
2rNjSLU+dPx1a8uu24d1VQzXJNJM6TmoDd3oBKbwj27WcXXQZT+z5UOEQgMD6QFqQ92rrAlyHS7h
d8o5RC/9kv4ki+ck1Xy2LtKcfb2FYhRUJf8SHVTFpVWS0KOoO3QP49o9TWzOfNkUk7xqeYdKWEn6
jW9L5D997xQtRx8BrguoKvaruYVbUekgdCXoaCEgCAmJvpX6Z2Xet1zBZzqEh1ZVOv7WLABel+52
aCBgVJptTM7w/NsKy1AhWcQM2IUp6HCjke4bLBXMU4JX21+X7rntUT+tr3kxKH/m/h2Lfazhigyw
ipswnaNboTJvnsBS8frBAezNvSEM7P10kMR0J3ApyU/8f236l1UkqawgjoKRCojz6GNbaaxEcPcM
Rl9CleGQHIaRsje6nEgFDyiFhMnxeSuwNPLScwZIRsvjT7znDFguCo0U5bAegrARfzx7Be+4+mgZ
6JbwnVB0wexXd+olpyyHkwVMnJo35Yx9N0mlMMOb7mRpQ34UDmwKZr5X0yCQtUaheaQsXxxhYq+0
SZuoZrFAytPIQlEAy4Eoxz/oiJTtugAyfrxb4e6VcmlNs5NA4TEKIWrdTHlVkdcxz9iNSSRd5r9Z
AHJ/XkFASGjbHYgz2boZ0NdWSSaDfBqAfp2AdAqFtXr8/O7tcf/m9/8+lp4lYB304Zfz2EDvsgJF
0TT0BM1kCfxdl7gldQh3z/ISI5Q1GebCWA7WGKhqHdHVfeCRLrT8L7wY8FKiBOVAZPWXVkmSU49U
/H0mDVk6KJm1/IEpMGOz+l+E0hteaDcL2BcCrfSznmQ784CD6mtDsQ44dbWAlmYLfumCdhUs+GTT
1/NnW5aXj+ZF65U9dDcsRTHXEH3JnY0TaTMDqoGZVj/4I0t+ysnl0xCnq6wHtYRFJmnZqDRaDfoV
yT20no0TS/73beDAj1rCuUFEbEKBFLZAX9s/ynuwE3x9mTKN0YzXQGbwcnj+Ofo367nYMDC05wPY
FUWNLYwi4J/DFZKC35ofJmja0h/fovrkH9LaHHY00cxazTocxe5ywbA0x+TmZjSJBw4A+1lPYjyb
dXt5FavU8/mFS8CANwaeAUFZ476HJx8PlzbKpwg+oy6VTmeTQGNiWptzG6TqGLaZ1Pa7hWAaHN6Q
dW6eBF74+0kaUbLRrqhaXPMg5VSrwiWf2ST30DZEjHQgtiv0vvRyeRuaa7QDn6L76g2dBe3VjP/k
wNVcqt8e9WG1FDyrTBIl+shB+Go/+uSwwtZ72WnPiBqW+PoO8wzBnEoO81O2aByLLQI+DrdyAMqj
FODGZ2aoyPJb6n2+Ewon+zLfS5NB6LVFfkYVCr5NS9WAtLcSWAwKINLzYhxXFgjUzaLbm5h8J2Bb
Wy2jwztmEQzJceaPNvg2FKfEmPl0+UDpRG6R5Yx09vxDDBnyNG/D+1ahYjSsIinfgbNGdpAeRGMS
CN8M7s18Cu6sz8bxxE3m/c2c7ynr5KMdVWhfyzgoXjIuyd6pHbKDFB2g70nnIZDayxfXY7bajTLP
lwvn0Y1jKevop1x2UamnKm9UFbwbbP+QsVQRYGWTHNw2NAWWuIxX4ovwCquQOjxOx1+yhybaIY09
p1p2dv1N//TWstAwCph63aziTdUGYXh1iDaRBaZdZecpaLpu2bA9/j7zFMiJ5GCUQKHhcVl5zDmV
v5nU06t4nXBlr0csEod0oq8mPP2lN+uNOWQwd8gAqqY1J0R5yh7Vi0aeDzvQ/FddbaCC8ZAzZYOS
dl5dQx+R/2Uqknc36tsGt6zLWZNK3+BSNnefMrkHz5NWPdGqVqOxrds11g/IxM21yzMzOdk20aDy
oX+p6ls0QgAlLyabqVio5vxJO3j0wVdnvZiMnNKJkCFLz21XSju5SHguiD1j2KBwMtMEPO7ZJmzx
fTdKSnfjNKe6s/hv+PxRCkuuSr6UzV9yJxMDOq1QqSsL9oQ/jPHpBwm26ngRPvZtrLcdzDWHB2wz
W3ZQnSeQr99aOtcFVF1u1PwUZTz//zIpW5NFjJOO9b6Ig7/4h5r4zDI9LnSnJuDvw//NChbSIrBQ
XdEwwPHP7ZoTDnxSzMGE3n8TcSzBPxwl+GMlRegrgz1rVMbWBJjfcSh9I7G5iXjIL9lKt6ZhcZ6u
uOzfbk2mBdHOF3Z0tTm0gh6jH8HGrHIxO3HVLFETZXiaUuCoDa10/azOvmHkhs+Vre5JTqKG6c9V
bkF1pfT4Nk7idrCq4Yhx6wTXUmy7jDgk6cF1dzp6FwW0NIpwRXpWMuquTQ7gqp1+Y/IgZKhqrThm
zvYBacevv3jtHnLm0iMhegkGfHlluojTpRiIOVZKnEK/PK2M5pKoOjMaV7C/tD2vZOITvHTeOkOy
qXuA0WzNJbmZb/LeX6FRY73LHLSiqgUQQKnsO/CBDjAnmdlwXeNbHuV0e7xETJK4WPDObI9adHFY
hOe8GFdxmPNzsM/qs3ei7e7zPBmARJtTfl1u4yiSQ/zodoOI4Fwt/32G9dN0sLok+TImJPBo7tQX
yZ7zC/u9f03JyFU7MCcwHplaOHoe2XN9VmVy4jtO+jDpu7Zk/TADKX+OtkUB8gy1gn7udd1a1ZOl
xDtYOpVwGekTvCCnNwRIFMv3j/z2Ls2vSefzCYlPZQh2vELzwct6XatZicKqh2k5q6MRxPkyky82
fdBsJDf/uC8Z/fyD+ee1MJ+vsZ6DRReZN7A1+UQXRp0YgFPckMVpXO3N5BJ61YhDi3osfHW4w62K
kphEOti0hNzJ2JYzOW6S0EzdarXMzO+BeCnJtrfSMu+GgDryGIwghGj3Tb0hJ7VrPw0qC9jduj91
z+6fc6G1qMSakCS3zGbcG7SGOe0GzUS22JFKwzQB+L9XLim5Q6zmC0SdUIRdaXEFrrBGIvORtCC8
5vL2C8PSp8gaEftRP0xuBigCm/0YpMIwqHMyTOHg+j3qwxtQg//pQGf3zLh625AWBLRihdQqlGZs
llx4PNY9Zyv4HVlXA+OGOMj47m0GmJAD0SvNf5SDpyKgJz2I1CJChqlXppQHaUOjrz2+tvOXn9Ok
azw7dXQWcfiLhJOEOgtVsLZF5oglecaQvizJZ8ytXPNRMxigW15GGvpQOXMgM4gAfu7BMnX5MWN5
5guUk3mvSNTyssAqvTTW+8tlgjIAVJmGz5FGgN5IcckZVN6XIDhL+dW/AqiLGfhGjD4k5Tf9aUuk
Uwi7AUa/g6n6ph14ZLUVvKh8/7b2mBuu/Mqz5SOhKx67SN0CbXsK6ny9Dllql3+x+GHOCDeHy5ad
E/ml97CYaqMK/CPU7AbshhCf4AHjrzB0MYlXpkp3s+qcj5YSp2UJQK/Lb0BsVr6kXPaWHdFWtpKL
2+XewE43eoraHngy8AYgghHROxg6J5OwkmXlgYFNXy/Vo9dKZ78WcV2ElH+hX5I+2sNRDITNgjrP
r2c/+K4O+oP3krbPFM6A/ckc/X4ha9e68wOyFij/iqEDfeBskIX6WUbVcT0DyI9gOogLsie5DoKK
uRO8By9tj7MFF0S/6fUiJaoHDmyL8Y+SKILOpkAxPNmJfd+JYrcZYuZaS/73xzdhSgdg2RE2HW7C
DsDshAquWAR1sVGMHDxKTYMrm/7z8WhW0UZiXuMZBsYcYfsReumrX0QAuJ1ASj4XE7lm2r+cTAiM
u87fNsE3SkQ1mHsfsb1moOfKxdP5UzE4uBMO91Wc2OisD3G5kPflX9yjYX2uBH4wj1M1sePOKTAy
C4CgWl9837Xh39kz+PkVGE6TTBN2ZUc6P02K3NLPmWL1Bev1ePV0a/iv82aejfz3BpTB+FNquyVC
F0twBMofHmSwQg4zR5cC3uMa/i6yU3sp31cf6epq1Orlph49cU7oLQ9fsyLH+r0vqjTOpLKbtGP0
nrJ9NngOkvR8Lr01dP1ore6V3e6zsi83oLlsYGHBXXkM2xEdyxPbjq2XDPOjl/2m7dXIujnLu+9b
V0jUiygcIcDLZ/uSXvexOz/e60fJoGITwri6EmSFlm0KUN0evqmUI8QXoiBoFDPNCd71rzDNIYW/
tIwNygYA1pQmlMbootdEcLN4CbtQIsbNq5jZdBavYJt2eZ6qOHDP5/ve9M4lntrYdN2yd2bd82O0
CF7m+maaxiqadKLmY8KIvYV9XuorETMa3e/tc2lexUQozI8A4kmtvnbVyNxaiOUdZzt387VWd/jS
/HMLLeJ+A3HETIgBHwMhXhtpoalGhJMQtWy5BlTVXXnxG0n097EDtEg8z8ZK1AghAkSFiOyTo6x1
QDXFuR4DkR3cRR0pYaVkd2Y/tn3zrHPk+64lVPZlLULz9tPr1LYVseZRLNSLhNidRZrmmktrev5v
aZJubpc29CLhHKBPzyr0TvlcEHPuyQPP5/nHLn3uq/rF5v2Bv4iyZMZDmyq9Eez6NijnxTmKS3t/
Hfwm/P0frexRKPsrsn/b4RubHAuhxJbjoxAgE7VvGqqMlMOTUy5mVizQeKYWbcDN3eDmrp5eUzM8
uRnMfasslp+3T98tDLSveavIY1bUdt2h/JoJOH9hsmMcnS1GpJmIQ39LZ0H2aBY29UEXWGPTGA7/
rPyniENMLtlIQUpeLimJbqLqkgLbnU2x+UhrPf1zmZr4cR74HuIBCYTitDnWtKnTloDQCf5Cyw5r
q+n6GMGWtunFrmJ+2WRodO8vC+XBwERmlTDXVn0iy21KfHugqsarWpIGL3jGBocDKSbLqde7oJUP
FojtAAoM2aGe51kGud+B543KWZdXaN2f2VoKOs+fH2ft4VLKLs+bh4yPZciIWvtiNWI+xAZ84hAV
FeuYzL0Nd+CB84afg/hAARfLLsizlRl4ZeYDU3E2b129LKSIg3vJVOJN9d2CkaIQibcD5CpLj9gj
sFkcOHIMt1FXrPlbd4MwdMksmBtSXeTHCOr026AOTdPb/rjK9BZ85i72+HE6PvYLbZZAFzj+cQqK
WkISOyyLALc5tLZwB5XxZvUnqKq+olNdpkxRzW40Zl1bht9sr/9B0BOYFpj/8yytp1DXUPcpeMKD
4CFbFiMVdgrLTZPPmgBTCb4vnp3Mez+7Euug2hshYYStBR4KBktZ0pDY8xD1y2ojHhk+siNo+CtZ
WtfH5/tO4PC5q1uy8r417q1UmArKp5SvgXdaFqHmJovyZz87AeKEieNfW7vdKPuwUMyYK2fdQWJH
gJjSnSSQpUjU7BZUMAGC9DsSFjz9oSsnRWZEDqhBgL5dOP8egxegpy6VWlSLC46JdMEmaRLCjorp
7MXNVQlvxQs/rCUbaX4Mpb70bni0xBefpI89vSPjb2mXXa197CvVSJRIKyqQnuhfYZmuzZUaLz5j
Y2LNiIGoUBavkCRzjTlnTGPak55adSzluLW0aljos3u3Is81W++jEsFmgJq5aevx/rc2u4qQtuHG
0rW6kiwauARYi/SDM+andboVUkWhJGkg4swl8g+S2gGPvIdjjFrlxxz06pJ/DPuBH0rz2KYpkgK0
FbZChHM4PLvYZquGomKsDmp2GXUGGTwVH3P86yP3IVY0BscuUH5JI1cWaiM6NfKuMz8atxnTsR5R
R5jRQlB3rAm3HDRAgdEk8vbJc3kyuSRmGc+uSSpzvMFaTcaK6+CcQYbQbJxvnimRBgEhnLQxm48w
AtDpbT/sWcWpRYoJ5uMM8H8hBneftdAVvkziEW+x2XHwi6/wHBUGPjASOR95wvque1AVDR+KbwvV
HJEbFA2gscx5mSPlyuahy3kQt0bEm+nH73MCuuquP4z06G1n9huPC3cnon47F7U01kgKDWGJvInu
eOmReSjvLPPaMKfebfpiXy+T0uA0ZnNojZxHZlkgVUFCWkWHShl0ORXZxSNK1uKQUGYc+9NKSoV1
4hgWt9BD2l9FO6fa86VEcGpc095NQPIsilXH6g1ie2y7QHbra9IEeW1khAwHX9r5AHHwAyo4EKcc
RBmD/lIWVh+WPLVh527Cp2K8PmZzIz6TNoVZu9j6EOwFS8r+t3C8eshXOx4auqCyLItgvD9ATR9o
P6Zjzgg/2U6WNUXy+8fgjx9v9NNAZYGAhAlMA+R8tDS/CTEXPXJGSt2SQWlqzyp4UyzyqYakCBQ1
NkyfM9i1zFLpfz9btyCnUcHcveNiqouMNeQpn9+1NWk0pFROq6Cp3kkKR0ry5wYYL3b7dOZct9jX
prsjC55qQ5M4wXF8OAop+8WVSxwfj+verdocfEniKvPAMELq0fWXI87x+5PzZsIPaEwfRe/s+Jq/
mtaJd49Bx46OKIqaBXH54l8nqF/E9y8W8WgUloFzXRmDN/T8tw90n/qXBTYazV1YLz1IzjdsFLMA
4Zn5f8FOTZI8sVFIq3SRpUFhQCuh4mVSl0FdpHzU0KWrSPNuAE8RNmSUX2hPH/5cdZfyPZFC+7qe
RLrUUQ9Hgu7dUOqAkcaWauKhY5Z3cul/PQAAysZssc734r81fd7+8IRjwmmbpLmj6btzyLq2y1IT
4S7Q5tYtq2RDRNbm2Lok08azhLhg8pN40dTRR6u5e0nogaTWB6r/mvcS6qs4Viw5RhL+cMFGgAQo
FfgsWMonCGeNG37rPg3YWpKEseRG2wYjWP4Pw9P5fqeUzmSolqPqiabGwYw799SNu/+CVx+lt7Jr
Of5Z7qNSMqa9ZFEjQrVyXn9BBka3JnnrgKkJZvD/c7LdSMhu5mPIKm9ThX+71lLQUJ6dgMuJ22xK
XXbfaZ0hsXy5rQNhHcyBF7ixpKWfYFJ9qAyJeesOfDj8Ng21qfrP3Yc9x7zPlDuWR7fg0gQjzvh1
D1o62RZmqIl7g1PuMx8a+9Vg5xUX7QbVLUJZMCvIiwK3Uwuumoh+wNGClF137jKcJmOyDt70/TYq
59VPeWxAPzpyt7dOctt+MH2bEgcRDRtaxpTy7XeEij8NSxa0XIey9o8G+RXEN55jOG+OyXIuw8Ge
XZgN56JhwBXyDZDgcBoUgOT/AMRWkEj4JG/VduyHBwXB4pBlp2cagVw3WupNz2/Gt+boyoy2N5Ot
rlrlgst6JPldg8t663emaoXQtWy7FbMgbLjgk1A1KmMTbbzM7B4r1GXv8l/8iPcnNRBXzU8wFztO
TKHpkSkMARozHjwUmpD2YFagkFHtBc2KfysZcO/+0JR0doGIz0rUbA2ezj5tjflln7PWzI2p3EwP
FIzoT/FdQu1AvVz+v25G+T6qRMOxMg30OniaMn4tc+fIwqGGq/RaJXnoVJMyaVMzfozhQPJUHNJD
V/6VnN5Epq5Gbecv7HpiaoG/6sbG8q0mlM94RrkCcC4EhUhfFVQRc+ApYGQ5zCCZEuxWfvHzA5w4
ERQuIBTku9MVunYwzCUXdqWGQkG9B3UJcsO+s9iE3e+EKpTXfOvRIeZ5g4qZ/ZE/WBGRTJWQOhFs
Y/xjbDRpqbjV61BZ9C1KXA6bBAfza7t3Trf2BMeU2+bkM7DpWGbR3pUBC7H5EAiuCiE1FyUMLgRs
eGCR7mimWA32C3lYvmjTrIg3RrIPExzPAbghUS/pA/zM4b9ChoR5P2M7Zcj+QYPdkIVTvw45JMvX
jZPQEVlZKAZMa753rfjFTZPGnNWfxMw7NmhPuJh98ILkYKAsEsW4tiBZeS9XSb7n+gmqnGmnhhnE
mNrt2k+LHz7gu9m96tVzdPN+5vksC0qjMZA1PT+Iq4bOfIM4NER9Shk4Smyx50jGpRcxvccF6Lp+
7PxlR3PYkB5FdgurFV5S1KOTekUHl+UPUgOrgPVXCaYXmyB0AGC6abPkOKepin12rhMA3Kw33pYV
/klVsY1Ti2+PwacIGK5ApVpcLIl7HvUvVYPc5QU2i1DRfBJsR/3t0GDcSu8/dizcAHh79BTWqOzH
pEaC65McvlHctlltsq17Ef4fXI1g4NQoaWF2Bzv7sGbYjChNIssDsv7/c3hvu6tL2CYxHo525UjO
7P1fLagIiKQ35TH+bkfebyuFiPWZqKTT6Cgb5h9F7c2SV6H4YI3RtRmCYrEMfM6xfSSoR4/+pmQ3
0sFrVmoqaDYPo3fegdzH2C8y+Gna3YCg3OcYMXvTT23a+oSqsKpNTybDVWiMQrTuXh1hBYMK3uRW
34Dd3zQfIlqRoDA50op8W6QAfp6ykC+vFpBWyxJIy1Q+55sEf+92PHC13I4Ri3EpCj8DDKEN2/S1
ZYRy1vmEnYUsoIN7cShhYilfuE5JfCpuX5By6oQCKLLNt5OgYZR2kYsU9Pd4QvR9Ivy8/4Pg3OzO
iCONV0vqz7nRfHIKEW2EysuPBx6eVTkcFaajpiSruyd56qbqp+u0m/HQp0a2p+U/pCFtvnGATJ0U
59Ta5we6Nx1v2D8wfvOMMqS23yjl5LzVSNhzaKzyOxWdJ1DmesouXKNLxz8/EFtAUpicEB6r9fX9
HEJUpxEmduK8MnN0MjNbC9aFyQLRbYTQqUFnXMqLUvDrw6uj9I9obBG8z9YbHPnQPvJJNeDHJgzZ
i+KWEl41gDWBn2Abq8x16SVR6vlzGc8goAY7EjrmU1WrMWEhdpHalnAiL3EJQIvc52AKgK7o+N//
SYf/cUaA375qR/LgDs8B6LquxysWlR5/OSBC8HBxye6NOtbylqNUw48CIBmKi+hSzhIG+RDFzfJ9
DEQllLW9vpjjlFSWmRerk5ucYpGgzKe++vidz8p5BbV8LSRPUQdiACbWCxH+KLSeq0cm11y3QZ5U
ZfwIZe7qjyDoNI18QsX/Kw0tXvjn0kU2V1e1X5Evia3YUj1Yg6KDTnmb+hRKCfSBg11c0s3hS3M6
AiHgh4k2yi9rUFRYbcM7kAJ8DzeH7+mEx9vuv1dyN2Qx8rDDhaDHM3tBCReBC/Whpf+KzbDTBrKc
eUjRrozBdPxNK+zZk4eG3sCX0id4yqHRhkFu1Sw80fCpJy0ED27lQ/tVSdFzIZoiFYf2fike/vh/
CbZxFA0C/1cL+KkVDY89YNLMV45DjQVM6QX/eLBT8zb0XYGYqqLOTm2T6atjbuHP6VMKmZMBJqgK
19KkimBuUU4UWvYeaVsrF1y37E9BKLXNaHg/Odx74P9ZiVG+1le7PTJhGPKPN86wk69utKFUX2wK
Zk5NM81wn7BdkL+MjWWuSt+k9liacvl6HkLfylOoMz6s68yj6B35zQEBC3FIbbNO8qVvwGcg/NkL
PaE7NtRrY5UpaLGFq9dGZqUMuG3/Og982Dq6pdrgPgglBXRId4DoFUcqQa5268ewuKLNxFnLZ6pr
+UG5JxZsKas23x88m+UOCTuTQboaflVYdjX8xosdEj2ffogG138Rgwd2kIQDtZHvDodzFagvntrm
0Ib7blpECXnl1m8GXuIl6LcLcw+wcn27pU9zeS2h3gAhYknpo2qnQtbusLPr0h742yqch/oP6R39
qlih4m7Tj5IHVQajyD94a4uwGsVf6qLKq0MN7rXwkOu3qGKjFBJYbg9dOfJ59kuREqx1Wx41RLEz
NSa1qaFJHr1QoaPLBoimYbZ+LLtiWayRNo2Xb0hiNUEgW8jWdTfjgpJ+QmXvW5FG7dSb9C/WlbwO
XrJNFXAFaSaWtpXFV7qm1rXr5I6LchDt0bVMtqToqhW92YC+QCgxCe6Yx4ZP57DC3PjtORXSnTC+
KNxFEayzXpnRxI0YNjObLpuxa69n+r0HDQg1SFnqYYffbFe/zkaZnHOTclyd/en8rFLds36Y0ghl
Ggfl/64TtSYibeQOAcw8ICr0YuJIBzljaOu2CqMnYUvPDPZ0DkzI/1pz4nhL0qk5DdLnO7nkXRBy
zjRPoUG2N5E5Am7y7aAlZ0EHU2Nu529LZq5xhQUXUSdU8JknaAFynAOZQsANCctwHqPEfPqMreQv
U5eSBcktv5RXtazRpaY+fPT6WdGP60KBTDo/nelrv465XpY6c7LISoqBqpYOmuqHzLFoi1PAeA+B
NTbHVGoWTQ5d/OfZCUdAmvUIRGV9gU3+tvwo4nKQDFKfKczQFnXKZDQFeI5crq0mUdLEJ6fu4N3b
jkRN+MdLRUqf7PdACLjbqUevnuiLrvMWjc7kg84zg66GG1Lt6n20iLrzc8191W6NRwDXGGrNitHC
wGMcNEdHFTEolZzTr0RaRZOTGUnAe5IQlWe1maq2j7crW9DIMCi4sS+lkJ3d+lwKoOJDLnHunGGz
V93WcY2iz49pZ8ni1vvDrSwZrq/2rsdd9sMxZBbeX2HytJ8Ibw70DhaFgmwPNgCND5habN5XdPLD
w3w4xb9sWnibSytMwp2/ANftINQMnV58rkBAP7WEiHs/iPhm7wPrWOQhFcDpeAOF4ZrMJM3rqmHc
+YUA0m+Dc+myoF5zeBndqYRUDltzpsdaSB391SB9Fkuzwcwg3r0U0W7M9rjiLz8HsJUZguM18U1s
OK5Ix996Z57J1lk+iQchdVs0B6RQWDfBfczCPIumYkazpEZb0GKMGrdWbaUoZ8EGKxpwZayRn6gn
swXyetAIvUfDuv4gfdjsVO/8LOswkF7ltgRfZScJzxqxtecFhchC5mtdCm26zNQZRLY3SUY20z25
Dn7b2Uxd0XwYfgYUyXAHCGw2rF23Ji5EwhvggdYfWvmaqHTwbE/SVsDO9JKysU1OLBZMifuKWNiM
xMnAi+QQ+E/iaffNk8MnX0ljy0rl5inQ6JgRqozvfki7v6nagWoLRkJGhl+AUudPsjSsmrz1BCuc
+ultyikyOywbC8LGqqPrOOsS+iaGZIPgL92Yz0WHEqXubILDbycnsD2jtwExZy0SMZCnw9xo/9zc
tfVexWLb5ICuyFwriyY8iaWSaq5n6eQ1sB0UGdoQpKZOHHZzrQ0+v3p9wR7OP83VU48dXA7Hy8rV
utqMdX2oS++ZuDoZIMt2jFhk7HR2VWYWdhnI+ShJLEGxNVgRWXdO6RwNigJVDQozCyYOWH+7/Rx3
uwKUSrfF3r0+NPte3HPUrz0wkchGGv282t6wJmQ6eGKxXYc13AMlZxCP/bteUDPnv+EaLH4KA0t1
wojWAN6ZVVpf9fo+cV+331Gw9u3r5uG7hwQeCRWr1unRP2Bx+9IsUEQoxaLARNgq9G/8jwcWDljg
8n1Zy7Ye7QTUeGthOtxeWhRgxvCQIohOOvU6qEeXUGeTy02P2jX0Iq/oQYJTbaNGHaSTdlN+muxS
Ph3GFV52BsRRYH88E0vYQHhxg278VtDbIIkKTR/X3aijDBTwQ4/LSwn2XmCrsmPE2FsEWr6qk/TF
BYP1DuK7vwIapqQhmaKjRwG1Oyj2NLcXR1mYQ7SQTyroH7vOEyC2UNI+yf9XPJcAbAVN6+bbJ8Ui
TFJ3bfsGUqshHSeLzW0AzMDtINnlt0idLdQbAggNjQZ3iWGEnlbbKRxelqvgz1k8iGZmmukH8i+V
3qGln3R1J41emEYKj5DGcEdVhx0htHKEhqWlPlfyePQrkdpfXDUrahlSs/L7JYCT4dtk6EekbfSK
pLGJ591jRqtzHkOR7Q3iR2apcO+oYn0m2oKhoJ/v/zlrBYZmXe28F9895TPqaC3DtJqYzpOJYjcd
jPS/E3VRMwROwrXXd5y4Us1azBd/KD1FXDnu7O2oW4e1bU9PLUw2H5rPbVBHpyaHd1pKsXVENY52
UDaO2z+SOXL3rAAGeN6sVBem4q9X81RezfsjG0a4XkNECkjSnIQmqscdbo2wJUjwK5Hotu7K1psA
WWfRJ5N3vTZMzGlbDsd/74kbwO+4Xc/Jp4ZSIb9AQpIWu6aM73WK28eUGUHyqgjM7YJ8R+Eh4IHz
VAkObwS+Z0QQMSDQB64ID+Gjyf6SxewjDPsSPZhVin77+epLsvcA+g6kD5bLbS9IFDwYohFJKNXE
IWYKg1o/VFGPi7InVik5vhHOmL/7b0hWTZSMky4cyoylE16LpH7XQMfDf6tjJlXXI93Z/zpxHg27
kZPWi3lhnbv0FSLbDhFDDbDmvC2Ya5EUH2lotKnxOSiYXC5NhwBGzX/TDEQVxMGks8TjDYidbcE+
T4zHoMWZzDW6/t64Z0Ixbgpoj0DYksTdAHt6BxkXMR63u5odo63VnUBVQeBjtvAXr9y4sTQUIFhp
5yc/im6bUBYj3drvD6EQhTEs9T5wPVmLs0RjsPukCJlvJ3j8JcE8cJUGCR+t6w963ZV5evhYaST7
DhMU/UbBG8h+urIjAT8MAO1othfwQLOo544NW+lpbBC5fsGBPDzi79SD+l80sq5hXokCHh+Yc5EU
yB6hlu/9C4xJe1hLZ0njGeJsiCK/rQzPblDOS/cJvws09JQHlGR+qiQ6Z/3SPJo6eII5PLD0A7Fb
c1M1qWGRiqjWDJy1B2bmxcvHYBGVh8U7Zh/RBpSGKswNb1dkCNz67B86IRFox+vFeFEcJVxdyJx4
+atJdkc29oCK4BhLmDE6lxO3CsYTlstr0BXpP4B17c33NjVcU8AOVWfKWy0K+cGnbnYF84yGExXJ
FwjWghtYPEEnZrAMGsio5VfSjC9JPoRpU6wlDOERz9KbPJYYbvFQfIsUlqGDZP4KUM7H3f2bmZys
UB6XDNvA7eEysAB7cZArLjVTJwRxcuV2kFcIo4yp1m+p3UBLvw1FqkgcvDFBfReN8vDW50RvxS7n
/1QmBcqN++blS833eKX7aMmOxcYyQp9JVZsuZzJ7ungrlN4ZKYBNuBNh6YRnPyk+E41u+/qcCQsF
DxmjrjgpJFv4yQE5zx3vfunaHhMF9DjSESxWc3MjiKjSlG7kMNVlBIBfoowOd/H4raspVFiTyQ1J
jha5RzxE5DgC8Bm7a9V/xkGP7FR8cidUSZTe6zxViqjlvaj4hNwgvbcEGeOc6nr46Rr9/eCLfVBW
eLvAXTA5YumTRLYbmntRZl016rGSq3Vo1QK/HE5KL/Udi+FoWrdSAdZJK2Fgfa+OocQB2Qb/W2Gr
RLhHLU3FUc+vuduB0na7jkRdYFydty83cOMG9kJ5PtxBhHhsnuoA+4dLWV7drFUCQbjkq4/fs8vm
EHAOKldLDBy0AP7/iJhi7LsZ0Vo2+xSd1vgHoukXj0ZQTksblIKbtTLuYiQ+Zy3KgWCW4l9eEofB
3Mhk7FLaPglwAaJ5X1x3koGH7KUKe+TZ6ubnM/lugeF7O0EKlEZNlFTm/DZcPQ0a2TPFYdsM2ppT
ufRAdrIQJ7H1LoOV+OdNQYT8mRMzUPsAudeP1fiDq7XMO1RDyf0/WY3Cl37svVemrF5dpLH0bNE6
MNkqPGpENnP8yiwEqgVvex1/ozgPZICKPFK5aY666YFLPtWYdEThxZZQu2B0CSeCuHNMsN3fSJ2V
Qc7N/bF+ZvczIwIWpqnyUPAWolcoalbNH9f1iTpOBtoKhS+C10/aTdPiXKwb70wogP4xGA+vZPHD
qS8thm7a2bMRSloFDeZAMhNO8tiB+SaOroPUYXQbVXMYjP27fG4ExBGtgKrhOkjxK14gauJOsvAy
K+C8tGEZSE/OsCXtrz5c/LKO393dXUUq/aK0ybbJeYhHCn7v02ZQA7ghw6D7T0gw2uQQLM1HD+Xn
HrUygGLsU2xWAJ9GeWy6LaqscC7+xOzSxpBPx+hMIRyMrSIoVpMmELLd3rff192uzFpMTE+1vUos
GBjRFWAaNQOoLxXgIaai8LSOCv3h2oCGYfNMLl3A5CPhaWMAUHPGu8MHST6jOdO1R9A+N6+RSzQ5
IlU1g6fqi07qNjITT7+Wyavrn3gwDR5M7+J3V4AZ8Vgele7lHFDkpKCTLpndLSo/g33fSnk/Rb6j
ImKIA1ImO/+FBHGN1mm1pN8fvj/lAAgcyRWc70uB3FdsCnbG75/dXzQGt2XmcEOfAOCoIagWuFt0
MTlyzXiDJ7ef7lwG/OG5mYUc1itwFJ5h/HKhT/1kPxuGHgFYW8cEN+PBLS1Nwwyfpp8m3sfDF9zY
XmgYAL/ICMiFyKU3Vm59hwboU3G1KPI8BecJ+P4zriLIGWLQUhRf6ZdfKkkQ+dKYVfwS4+8xn4Jl
zyXAWKrVkXYnYT77nnBAszUxYbdhqw5ECIMy0RFJ/WAuf6+J2H2DzZQVs8JqS3yIvmt8BK+7kT4/
ta022eWJLg6Tu5aOV5ZdROvN+lSgOgalpg2sfD0q7tgjyDWPS2m3dbSXWiX92ZZXrcqwiP/5jiGR
AECrbKLmPc2s89lWJ5pXNfj6rqVZjzmjpNUZ2Y3LDCL18lajll6O11ubT/5bSocOqdsvJH7VNquA
xte9MBKLLqrSw6RBXSlK8VqcvYJphhZTkTdxyv+QphyVYXy9hzQSgo4dfWcIg8EqvOlFPnbCSrO5
ILoVkUTf3AJxcBqtZ2ZscEoYw1LxzKmBZxhFCJtm2vvBrTzS6FVCVq0qPVtVRX0isVyL6RHrgfco
fXb91JROqKA/LYR4fJIct+RWeDvd4e4uNmB2yB0kfQzWMw6640KZBwQfqrXY9YnRd+ewx0JCdaUE
C3e+091ZJnr8VDqIqratuLnELoVVW0H05sAuJsSh2WzQyxzGm+CN1RL8FtrCm88lSVz7aFNml4bY
w5OuI44yCmxvtmrXAxmErJ/25dPAds7iGiendJI3ObioxTyPYGQj149vMawpaJgVn8YmiwXZrTOA
RqELTIymulOgWtU2Bye8wkOfc1iET1zZwuPsxFiXVhQ0ic03fvXfg2g69RftGTvN5wtvEelb+oz7
BjbvGGJCLA0mBCIcErse3yuH6uWnFPbJt1ccV/dnqGa7CNJHyoaaqLeZPLRPzVL2rULjqMfw3kYd
Wv9V5Y9a3g3iq4njOkpdMLwc/cto6zu+SEOwCZM6WnotUAuVeoVkL0gV/MtYjDNYOilnKU8UU8FV
X290IXNDTbxq4SmCVpgSrSJ7UyhaZ4F0QSTKC3GckpLRB4fYDK4LdacYLXb5APH90Z97+A7Ex2qJ
A3xlx7tLfDSeXpGWr+GkdCwHGjN+W5UwtksbKGaA08qYoqdACid42kBFqZ6vCZbnUS7One4MGUCx
j6gQMSr930ArbeK2eun7bRZwYhGxO0REqU0FYoE80Cm05A5EHN2NmZF3gNAO+tn70QunQCSPZeAW
NuMzUSGfMns/iNsrRUMX8EYSC/NVZGqhgdlMH6xSgel6J1jeyeckrJnIcvM/ie1Mzu96RoXEhcWO
Tf5cpvzatPypk2f/ro1r+8jk0iEN+3yGfsUyi6wLT9G9iykfpyyjChWgN1xZuvmwhleXZqaQNOVN
+iNau66dNDeHiBEYEW3Jz+hHipoiZ2fZbW18KBQMwDWNBafBLXyJCXvoQxJdbXJ7fYWzHiFs+g/C
jpeOPo2akHLsN27Ogru6Mu/XL+KmOGbIgt/XUVjyhRwHbiLf6wOYVAQos5cXYj0iFSWM3NsOQtoP
CpEtALBXI7w25B7YBzzgJuV4yzpaqoFNFvPohLoq2UN8k3EtlQsh7X+pvaDV86lx8n8QFe8VP4rz
KwHieCKkaeVybTLt3qsjIBpndr90Rhva0z+U08ckDIs6qQ5vNw5NyucmkMyzirAngGA0BDqoJNwO
8ypcQ5wyejr2pWpJ2tDnBTLZq1q7QC32qhc1m1U9KFG0I4c+f536c9q6ruN6MFNHtFroyfCsJicb
3rpkejqXg3lGhq30YdJQ5CwDCXHYuIo//d/23usTYElnefWfY29l5xckK2jLI61XbIG/5kD2xvtu
c4QvO3WQv4ZPoFofV46DhrzpjssaENL+LyFhEvtpm1AtdMT+XO2v/gt37hFOAfFCialFHRwbrvB2
sFiHqRT/lSNfcSIC7+i7A5y7C9tJk+OtFKlg0mIGgXI2oTOmOINSWEkGfGZluAR3c1IH+Ex275Dn
yA7ts01A+A4hIJZ3BHOqYGu8QiW0DKOsj9TBvx4Lu9vbKrYw5h6xxDus+ryEA0LMDiIoJoTxfXjZ
GqP6M/JRnfsRenAVL9QK5moLnc5Hoa6sjwnVwxsKfXSked967Fiq78d/eOvNlHRxBzwL9NJD8vV6
D9zPCTd9Y4OyvLK+KDdbKlVx+gqOOMjAX+KYWF+fuYflHa566NfLBAWT3dffzVUzX4JPbHtIlDK/
IK4woI+ZJP2Po5KPJMbSy4lO0z9doGg1pOiyquIJqA49KXEHWGgAR/Y/3ocRy7jutGoAiu/dmxBH
/3xJLSGVBLGZp9/7Jb3mZnLPasbw8aBuqadHNEHeyRCyM9kdpg1GbpK6874fSuiCor8EJ68PwAsZ
Y/KW30pL4JGL8pKvD28LdopKn36bndqVFkK+qNuMgghJLGbKcMGJWn4/Z11ZkG0X9dq4pmIzqlb9
K8zpfUg9YlZ2RuAaW1ilBpYzX4dKAkaVhERH+8644XJgfIbWO0MUnr7uEah+ayEVvOV3tt3ST7GC
OFdmDPuWb/qYyVk8ZrUlKeOfamzwwcodctRQtWj0sXSoA/rgrHaaUlKonHPpDtUk6uwttV7HQIfN
cY7ndtkqXAF2l+SLWAhmt+5goWc/QiL3qQBC6ZFKsO17dfQQ3anP4DODD+qWHw3VWiUD+l7XxnPr
SJnAZGsts7aa8IKO+xwcEnlap1+ghSgDY0OOVWVO98FOOK3nqqIU9XKZr9SbQplJRbM5w+6ksmth
zjYMEZaLMGIyiBhG1nlqcGlbdMcC7AjHyGxU9CXbOiUbw1x34sHaFpu/7Q23QWyoZa4yrQzHxKc6
+Qo5JKRnqN7Hif+pP3wBNalgZSGevNf9KGUSxlBtt7Yca6CZ31x3gIUpOnTsGpgbuGGasN/M+glz
D9qtA0VmdwAWWivnFBKLmO+R/UJqjCPGnUfrlTRj7YNEIrVnDEdC+Z7c0B06UQUUuIkobFw/him6
ecZPqSD4WRveK15jZfEcaeOGr4dVvZaa+Xmx14nITEgmal7y46YbBsxgV+e+3irh0oDg1msL73U7
XYcerakl9fWQVG7XzcEQ0NwgwWjF10icbwi1T1xqOxnPTcwiD69HGHM20klpvRml5XLe8dh0R3at
9t4ugh9OaQ7INSOcaGpedD/pp8FUz8KWO0sXFUpKs3b4zx02X/NXhIjgdKqHfZsKcDfyg+6ACXWS
XqKBjVh3effI3ypJy1uVz52TyPxdm/7Ly7ySFA5vDjtS1Xugc2AjD9TEySeZ4Jyl6TIZwI4v+DfV
d129eL+qpQnD0rLKfueALMHSZZBhsOWLpHjk95k6WzHqtTDH8KzSEQguhDsDX1D+1j3UixzZy3lS
dyvo9NlLLn6ldJWNqNARdnK+g4t+IMEc9ysfWdfThXNdwjB/BusL7GTkzbya6ArqlkcRTiIKautp
K0qxpYWFIsxsiZsFABaY9yN1Ux1lnw56Qe9GgZXc/NPNW6XWCEcNCdAbNfRaEghNSUhxegcL55uV
56NVxAzbl6VD51fGtGc1EkdSJ+xY4iJfIakBTOaMCzAHO9/OaqC/URjeoy4CkwuOYHVQcRzJXE0D
rhz3DFOlr4f6dkwrFatCHu0neagwOXQSX8h1fh9lK5kXG2Y+5mKHj9ZyhjqcwKZd5GBZs9em3SER
4XM8h+0nQXOVawA6v+VtvCh7z4GkLsGrIZOM8x0ck85b2BI8BDJ7jKkUz3qBh8wpHzgPUK6005Q1
rqPhjWpZwYCOTDa5I9eEq3l0aBYrA4+nbAhkV2ZKt/7V+eTf5fVum8DO7Ap9+Mfi6J1SFnMLu4vV
UU3PoxP39uHPJEV/czvDjAKRdDpIiVYnYvOxNfz8HR8w6lW73dQdmsLtQAdreLNBUyWjUwlxFof9
0xBDkNuidmqqEFdAzMWKMlCojJ8m8dU5VjuO0Kl3uNieuXSvKS2PCMJd0z8fXKQeQ3MbcN59bEHP
gU+ugDJLguRTgo+Rklx923Prmnsh76XZKDC10ONHdVZQnvjDtFmMYxw2W3Uct0ZNAD6IMGlsCsQ9
BQoNIRyOdUINit26QO3YZQ3x9BTFf/TZR7Rm7invSsOOprcSeriXg+pTb7Pk4ZgpPgcVsMnoDmU0
JmGorUezIV0nkKv7fu0vD7leZSyfCwUb307yb6aT+AkB3trDSMclHs9ool93HjkZJYBYg4NczFEw
aGwgXQ4Jz3Sx86UGaQg0fIe4TxcMrmw/p5UCpO8PC43T4izIG2qnwhUbE3pgpiMxf2a+Bid6c+2j
Bw4Q3ZBwXrHGo87cFrEsEdrTaXuwHO19SMgcEBUWmLOLLvJrS36WDz/2nxw7UvrtHhHvCFNiJZTM
/YZdNkVd5CqaTNbYoefSbNxrb55th1dibBkozD2KBiF+UqWYZHRcnA7fI5oGOb3Q8zlRCHLaNTSz
1I5H/h34iJccZhL3Hh5cPVAg7JtmFisL0cRhydvdEbqYNi0wlJUL0LGU5KC+4uoVCQDLM6xBMNs1
qAb62ixI9rqHwSfn4stmtKjs8pUXeRwfFXpRl9MW/mY9CwvZhw6ty2ZO3hnpO99vEZK5+bNQg7j2
hawSknj+YANv3L8zct6gGtr+cZPFQeSUGCDT111lX4/9feNG85pAiA0XQenuzndkVOto8q2vZkxZ
to0XqRXvwIVcCHe8ngOjSARDE1nA4tqfnp9m7vCOrwteL9FlEo0SHBQ9elxlgs0djeZdtJUg79+b
rjLWmYMU8OQrTO3KnFlR9SznTd4zJN14nrRcCVRWxWfomde54zdRdgFEApET8dHfPekEGiy8ZZbj
EMhgyAwYcJ2XTAEssFAHYLIMRF7jcTvSXzkQnjWZPy41D7L7BnB4iEMESAo6DGJ780I7B5wwNiKn
fADpdMvAvSS0ErzEyjSIRmTLrwn8P51MrzVHkHcTZLC1ERJoSdXp91gr8A5Xe4LLZfKQFVsPehR5
IDrlHG4CipL2CAcDOwR6oBfCRSOT4AD+9oknYq1r6GEBwjEIRI0wxvQH2HPqgqjT/latwwMfmvCo
PKQYryW7dlqhZvbOKxnQ9XOKzkJHvc+Uzu6z7jz7KM3UL8XjqdRB4jLEgXe5LByzIiO4IOhLmHSt
5GZIP+2JeRUlXYbL6fciFC6MpPbrgZtD+HALs9g7z4Y9DfMlTbPnDYxXuVLfrwXyAdYS4BSCSwl4
hP5CWLeouhDtizNIF2e9EaIu9MLe+Z4ZvcjOWW9vEHaRss9PjZW8Nrgck6BFzYL0OcLCBLbOI8vq
345o+kbLabuph8mAGl6mrvghNF4xyjSRRT5XfCE1IWVJovzMeb2YgjW0bAC8roIUf0+BcUtma6Ii
2E5x0Ymkg8K6O+EHEIQExeGuYdVKjzfDjs5spgbZEksLpm1EF6GAL1FjSKeTx8HaQ/Lsezr+p848
T+RoQwuwX4EI8CF37iKvc1wQ/DRJxnkC5cg10SqdjkUUHTV830OQT/+rjaYlvZfTBeoLGSTEvOvk
k2xgdLM7LpgYpE8t7iDBCru5V5ZukWLMknByxHfQVtmHwtCzucSlIfJfZmi3NG/rM9WSmyFFDFBs
nNOqn86p0+tiPdswUC7nLfAI2A4/zKYw8YhBB3CCRY69uYW1JZ7aeluBKXooc0RySL2fv2VusUO7
ooXzJpTgqglz0TlHBj5UBKd9dtPBWCCl5b3i3NgMcfmtJKTMXvnVp6Q6NCO4e0uuGXbhCUU1755h
2Lcm1cc7fpKU1+EBNYmby/fedW2XVOWmdz8CL7bK9ItnmlpsHT6qhVDVivcZ1lNDEahZQenVeAtH
a14RNcFiclAsJSJwzfn+qanNxyFOIwV1WZj1veOf0CcbxaiqwHTx4NB8+EJE2ur99L2KZOy24v8P
WvvFSyYiErf/rsj6Pq3M63aDPGFiox2M0A4noUGF5wXPUI63oVqhqs2XRcxn1Gb/wu4pPCQoz2L6
AinZ1JAeZRm+L+DW66NbpaNo7DjLqnkSiEDKN315lpEOa3EpAnW6PSBWmFHX3EVbjoMZU0RLdZfV
bTEpG0L7MvBs1uVG6RysU91thtgdD/qOZoCgtS7oJrpH5CrscI4JbokX3AiscC5sM7uVdioEpMVa
7oPVPggz/pQIzW3fnSwifydTXv6EWRboYhWiBgBpkAvwSQCbFPQy9WAI4Pz5R6qmotf/tD9/mJCk
dwD4QkyQWcR7HdZgdkagz7RDJ2xI1+McAfe+MYw5WBmRpvQKT4j5Ls+ffF+GmXdrscl41InZ3nOp
rj+fEokUDQ8yGL7eJDHM6NM6gfFHmfLFasJ66xaU3HY3JEEYsDlS0lYO9oROVW23bfCuYOkkGP5e
LHoHFFdW3yyVD3iU/LxwhuwPnqvWEj8XfVYn0cspQvzpC3eHf1Fd3tObNSpZlHH5cFx3VEsUxgH8
T85reeIVmsPcLM0YJncqucusFRktYKSGURG4XOXiVKpZaUBelgTT76wiSCYtranhveft4+SBBskM
vJ/oTzPNkRsaqDtMTXxav/1pOjWWoIv5Y0LYnNpvE+9KJ/2wO04c8co8tc/U1q5OcOU/G93GjR7K
0bRODnBd5eYT6WnYoUPwUM+EjbXfAm5FkNBaA4TpoJTZAKAtFU3HQzn96XVlSBQ0fMCl9OVhfGZh
QQSfd35RbCtHQxk30FfMnW3fuel+7FJU7RRe9H9Oka0PQjrdLulQpivgJDVW512sjeTMLeibmxZA
RdhjiBryn52SwUrRXU/WOu2BdbNFzMrKCvpxr8PziIrZodkrZauA0qaYuPySLLqhQjL6ysjtASrr
G/wSeRk/jz+A3GoRn0s+Y4ePLBEqsMEAx0vCpQlkB61Grgre7xXuqEvbf0CMTewJREy+t0CdKDRH
CSKfXxZJvIXQDYWyYfbQcAl3hkuTk+mIDzb7r0HUMtE+r2SKSRexZmHv4SQIrr1mgkxJNSX6cFH8
VHuWGUPINDQ06lGzepjkFDquUfLsoSYZd73N83/1JOMZML8mpV+SU/Xhqqp9LfsmOY1oUDF87iBz
ejoQI+S5fQ/BpvHrvY7rilmDw+o3XEz01cQJHHuGy+2uRar5nLKcC2WGkXSa24ZwAl+rziokmVnS
iuLZjM2fvWonlT4BmvK02TPGKYRQJ0gSg0clo4r9VfbAO5l3mlchSVaAYoBud9sO/XHWXjWUdkuz
Z0HWJk5NNFpg9j+E1g/2qOWdOm8xNSLCbBOLmdbMTtoAGafk1124hr800o6u5G453y6rIXVoyMD9
RKc3z2y54Q8XRcfTocSi7THII/UC5jfHYNI2pnPkFtWkz3YlaFqNWPA1hUx5qlbCuMjAextFWo07
OwLyd+W79r+26U4kwxcsCh8IeHLyeegLoBiHBsJJ7XCfv+CQBjukEbDGthh7Wh1mbRnnWs4R1IG1
HLuX0e+9Mpq5nsPgj1dHWQJCi+zg4oeV87Udro2xdL0r5zw7CTX5mhlmKKy3i78gCZopbwLoaMvv
o1XzXsmy5qoYwJzUQ0GvZB8zKY2bOTPe0uy/OW0eBQQ13AN+nrz2aPcqRQroKn8Sd982cuRf/jm8
Ajcd8O+5uagleWXfkeD7K7tfQDDmWXmMuPjwtYN8edQS9OHnL7K0bGajcVQlDE6PHpvCD5Injdd2
6X+DrDMOWDjsIgatbJek12FE4m1xgeRHIbNf8V0WuiFBM+Nk/EqrHwEPx+OmIovO/yN0T1GKDiLT
Qtk9UB6RfjWNESFAKAImUVYzXTLpn/MvbfR4Ot45cf+IPxUFYp6UHuN6rBeHL5TmvzxEnbQV5r/A
z1BDhHG9gPPupgvTehKkCZvE97eAkBkTgRvkWNqgC9557bNUFhzXyZjSkEESFNWclcgab1+aCK8Y
F+JKi2uK8n51uB4Mio8dx0u5ZM602faF3zfexb8C9c0FJpTcjFGlApbIWPJDPkGICaQNFB2Ruuqv
dyPjfIXiG2PLJ593vMohuVJCU4R9CBZnQAgTYmICh0NFFAYInr5lFQ9wbXVk2HRTAX+d1a7Aapum
wJEj5tOKr89nphJZ59G6hg+EvjmNkvJjCHPKYCJWK2PCn2TRWO7mlxy+uMNI3O4DOJm5bt/POTDD
YiNQPgPZj/mBpG/jjSFq0OhhT8OjuG8mOD9wGZ+Z5iEEsQ2evF1ql4GoT7aP2/K46ZLqFPmTj9Rr
nuiiyUMior/T8yVO3fXB2NlO3A5RMcZZLRBEAc6myxa+nNAnV2JHLQQtCFvPFVS4l6wFxoVVtZG8
AJOH5tX4HSfX12nJz3G7GF5tvtDEp5m9CF9l0XG3ydGIwWPPSTnIAcJVEn5aQ3bhgoerZx2nzvXg
gJTrAVppzbk8XRaFePXH2GG1LykytY9zq09EA5CQJOjmoITvP62Rh0I/PJC8EIM9u/EysVS8psDn
OV7Z/Xxtr5OqSNhVFnP9Du3tZVgw70dOff6HUGy3pVSxiQ69gsAppApGn07SyjHevDwUU1FzgRXa
qDpyDLTPeYZDlX6zgMiqeK/334e7cFNRSBatO/uQ329MUh6jt0mCc+c+1G8xzdnVDa7zbJvy2EON
kun/EnqozeZ7LPQb16sKbcfFyficsfM/jxHMTxJ+kwH3V8BpY+jd+zxtyLez9+z7CltHE/jbSfGf
VmTYTysyI2lq01b0tmykAZumBz2/oSwtQ0xgFAeMnop4sWiUzXtm51C8/YRlpaxq2uN3i6C3XQPY
qUYuLJH2M2B5Ih9opE0aYBpChOvagEJDEl8OqGTv3GjnoHyT65Rcowj/H9eP/UhceOOuJ/JHldS6
5nHwA8K6J6CrPSg7YzVcpyyTrbGOwVAj7MPC1y65zxkpk2R4q8DlhgnPK3Q1ZBJLG7tb/hFEHgcT
4MaJHH8YeCVhQLQGQ3qbSyrVDT2ZKqoLrpXvnTUjOVrbydfSTFN7R807HvNC8556zPHFQjMqmr7R
tOVz4ielxKZCMvJ35lqkuZQG4OsrMDGcG6NQCAcQRwo9zOAuSSMa5y5Smze0kJaAl97RY7AESQ+7
RZnL6gpex4ULsks5/Km8qN/PKbA1JDDAsYLlIT9RsF4kUV2yjBIfGVYYIbuKSs0Y6DH3PbGt5rAo
kYLn5oVKbq8IkTitxGat+t4kWDr17dJwbHJc1Xooar/+bnK2vgW4kLfUroZdWxRq0UNMcf88KGOV
aXYGnbBW9P+776qnYOk+3FYHFbP02ybqQOwaqJBLiylEx8nBh+VIGuAFRKGN949UbI10slMb4lFZ
pcl3APlCWFn0VvJH+cei4LklY2RRSp9ARQMt44ej14d5r5zqqiEVqAIWEG6fdG8/aJyolOlrjB/1
af7kcuG7r0qBgunJXa9pyOqUHK5kK1hGLpbEYgjF4Jl9zziz4NsGEU3JFbPPY/lml7+BNtBtt8nR
dCsHsG/Ez1WxHH1xgUxtbHg0sqlRw5BeOckcaZ2ukJg0HeoBlYXJdQKdzFFapZu2Rmnv843r4/5V
S+r8HB3KH+GSNlnSj/0D1ln+/h6Low0MJIB38hhkNAo+Zcm1J1TC0UEeUDtQWCzX/WhSdZY4P3Km
VTbPFDg20zoBcqNSFGk/k6D2UqgBTQZFMDXRQJUzVRxnC7vkNGEY1PtuMF+4vv3nFNtUG1rIfPsp
nLymHJXaqUAsCVAv4CHPH9SRhzrDC7XOmXjEQFFvlj3hz4r0lmN8pqUf15jEtHHHHPxhcLZRIRis
4SP9DnwLbzZUXFJjqAQh6ehTKD8HORlmpT1pCI3vslwP7H6abA9ZokK85ndUfXYqcVD33oemg2qF
T2XZEZF8PT+nWsHul1lxLZX44IFXqPMERbMNcz0TcDSJalv6IQjJwonqkqOLeRX9G2oVtlTbMebV
es/dKY1NCmmsXs3iuTKDLcoTSnDmoXNrBjVxWB/GYfKIPqrIiR+bSVP+h31sKs2nX9e9OOZZpWrZ
5ZHrz55t5a0JBKVo07UrdtHW9tlUS33CmiICd3tLsF6Iapt6j/2LhJTstl0uHX7/G9clCLDDalNP
0zcsLNccyxNEW/74S8QkZapilWe2u/swzMMisisYjWRaGKY0OTbIQd4D6Gi6q4hbRTW/5Bp26kkd
PsEkMdXm3jsj7xWCB1mC4GphOnCzDrxHPScLAItMPdGFUFeljO/GgYz+9Apzn+8HV6D1C0DuySqa
GWo1x9a0Lk/ONo7wxXM8ScIAdFdyg7EG7H9SNN7zj3xHwxplbU/IumVnlNFe/Q48xeEkILQ+GrB0
PDLb8LbZFwjs6EjWBxDD/nArqYQ8FQPsRH6GLNxr1j9lP8Kmej/UvOUPHgIkCK2cvNMV+v6mdb0Q
os/CgOTUJOE9aoaftSCL5TRIkGVUEBJgoRR+qdsbLl/O4tpEqtuI1OrhjYLn57QRP7cHlj0n5Xv3
oVtnWWlGu3vNOM7S4Gr/ARw/PJOkETRzLnnh1lvw0EPLUmYkkRZ8qXfw9k990CDoDgn0oInKGcyh
46+FJ/6yo88/nJngtqJ8ig60tLK71mtrT3bIAveVlMIP/K3prCcqMCm9FYlQdvXFtuN1uCqX1kxJ
2swj5KQjRzbCHtgLKP0cWXTiNAUJ0nCIOR4LVs6A2s/DLKbDVkxX5puoNHKJVlmZ3SpE9ShcMeoc
MXcLPXOpBW3BCKxxxJtKrjg3pduM6wWLtuG13A2W+HOOOT7IJvOU6arC/i3NZW0JoJdMmLCD3xVv
P9da19CwvrTeuJVwGHW3YLCYCf4tW3vtTAzUWC0Sh6wvo6DOHiNWQGAKefQ9X9Kf7bLx9vWroSeB
DnGHm06dQOHIaiFKW21l/UKegt726sY1kzZ8eOIOND7P9m5ytPYKmIRp9nvEYS96vONrT4RDL6lk
8zXU/bXLk5PGRe2K69UXPF2n6Gy3DN79dq87rVxqPflhgb9vF/QckBK8Yc9ibzSQtMTfIA6CPYoK
S18QQS9Jf3D4XLFB5kF2JQm9VGW1UDh2g+FAfAYhDe7UbMt2DWgZjNbvzI6DMp9DwL2VtOzu3YMs
egsp5K2Ul3Ht+myj1hXpti0rkhTRqsOUHg+XwIy7ud+GxRGE8nE6K3LsSBS+TF1VR3xk1DWqpYkX
/1e9eImBFWo3LBWqcYG48tKKQ2BdZlSBcvKVxw92hcPMMaZmxjgoUsVK1gUably2wwr4XcF5WJat
MVDPcM1gpbdKA3mELxvKOzlyxaOplqbMmZ5cnJH5lka/PcT8yUIlBhEHCbtijjWRp/b8f2cNU0uf
N0Lr/xmUlz3Y1+MsxmGGMR+j7LwIu49LjwY3Qsp46cG7rHM2IXHt1SGxpcVqJYVhG8PPEC0WZuVj
Few78otwt6/7ykpF+z8KuKn9ltms2WBmKeXXSGA66vPpIjDijdEo5RaK+x8PD52sXlW8avzRNf5q
uT51fotLwtNY736oaHmGkFM34wwErlHMNk1QGYBeR6ONw3mw6SRUqexNBQVhKoI30xV7nj5u/Wvr
MYh5HNWgNcYrPGzVSzZ2uQw+wEyHCdH8eYgtojeMmW+EpqyURSCHQ85e6z/KeTo+2E4zmbghhAdv
0j6vgdvPlKKLhzlXmxy/ksmWQMYqA+4rfAsYwln747xZGzdugupBs3ix6eFZa89VOanTP/Iv0PDh
G69wn2pzrwUuwgUjtiJ61Uo1d9Rjta2Um81WLQqIRk/xaLD8TuJYXC7JZntnT+0cns9Q3lRzOYaO
4N2HZaCwZIPp0Dty1BTKUdGGkiLpzqbtxPNyqq3mRIfrT5IuA7QjRTfhaCRn+9ebUTJNDS/6Xm87
MyI9UG8tcKC7fZnq/QxzF8zbkMNnX9XEMtFg0vTcLRp49OgXnH6lh7XJ4HYdjy/0WlbRScsvbAGm
7hzRKWldlPW4t0S8U0pb3hFIKAI8YE0LUGk9RNG+KbO7I40UwiyjFBl/fehQ43OHrrvl+FLP26sU
+mYsP01WfJVNgRP9n+6nAU7jblZcpZoWCcVpr/BLTHmGVYsemEDnxfLp20Yr+BLvMs2Idb178fhV
Kw35DRYuaweNrWlMIIaBODuz6/QjtVNZRiZN1+LvWawC5uKy3m+AfScygUScQXg0sjwV0hQRLLFX
rCOnyRj5YI5NohmVTsfkwO/EKVBLSFWflXyCYeWv6IYrWeVTtTKE4XbhkIXbuLrcDY6cQ9eEQllM
7LYjqsn4Ty9Rnjw58Wrw8DHtrXPgXZVLHebNfgTiL6P2pc3M1DhvP02hj2DUAieVStvfI0vw+y1B
PW/vDwd5Mw7s2AUvnfqAsUh+AVQtmU/s1fF9g6KhFolB3t5/0MUQ9LEF2uX9E9b+zinLquLLiy0O
VIEAqATILNa1TePz2pd3A6WrAp8thsPIluuLnZeVAbbguc7HPbz7XP5WpM9O4EET3sH94jDs5o/C
gMWs4Y7+iEMw0ppTlAH0sTxDhiBTAAna90vo198FeXxt68ln+VzqW6bCl0yPAqtJvNL5d7Bqy6pq
aqehUDD9VZbHsj17+pxxRayaEVuxlrw0PxOopMQmmnkYxEDBy/yxBQVbolGPtLyEBFusnzJqsAt8
3GKK/QNlcb6G/VPm5ztPM/CVkgzGg0vI4a8Ni2Zz9PjOxdhNhci1peH6n03q56Cjpx9BPN/gttmh
mPMm1YUELI+MBuvxjMA1GVcAei7QxuMp3uADr6TA3zyd3YZGbPh7nM6yo7xURsUpi+WyJetv+WYJ
lIcJF9UL7ZQ8cvWvgsI6wEJEdbtvqMQPfpu4kN6RY0t6Lr5vnSerGULbBRBi9G3ud46mOsLI1pNA
u7Jj21Lq14RoEHsURmnQSEvzFVI6I3UF/YeKCzYLgC4o6J9aCEeBgtDB9hS/cBvSZZ6J+s29Jqsk
2udcxyjsAj+IUlQ1Jh2pM9ogncsoz8PXcXufD8emyrdjFSGX2LW5rx1NUll9Jj2Jv9KFoTWf4OfM
RAwFR2lM+zBk+j0PCPlY2Pf9sizW2OFRdM+8CO5mN3UGqnam+4fksCRp3Mg4Lm+Z/tXDvxuOZPzz
QVyOCtFRr9a7vawyT1jJkfLeff8jAjh8eFSUeuez2MRI0VEZnUTbqJBtx+lkSDIk41EKfDmVgLoa
ZFpZY8sZpsKAlILbbx6OjjE1iDfpRlBcWFAl7e0GcSPAmqcGHkfHZ3VM71X/ZDB/QGIIcd4lag4W
0zRaiqz7/SiCN4hP59212aTd2kgH1LbraRiDj3VpV3jn1ilDZFf3sPfcYwvjSch2djOHZIznESCf
y5RDTK6d8NWzZHObiC7bDP5xD2MYPUKp59IwpBX2WhrCC8oPP6wS/mKlcjiJBGDrpUKRrh1mFIR9
H6EagAo1gUvdlrzVOAtDsZgDMWLwuD84RmHtOCdBKSU2zponLQEvrL66C83ZbMgfyhe0CFa788zW
mhKymoL6y3FD54n8npCFjylgudjciZD/a1Js/Oh8roDPZ8TasAMAD67haKtbwkBPiFxukiladaTk
pZJYOkg87+VYysomw5j2Rhc15SBUA0MMqitVjaZShD7cV1PitxzrAb7mo+aqORKBho8YFSM2uZ/b
Y3xyAMildvtkigkeIYuL5G7u70nct1MArcGb2AEOtlowZafHvDhp0yxvXnrrMfT0Tj2sFwZRlzHM
+HA584SnsZ7m09IVfL4Daw0+popa0v8bLk5Iu9EbN4vjklKtCBl5MTiPMCPfO/+cI0Icf2VGOiK3
+b1NCC6mkiZ09guNoZsqIzJFOcgKqlOzTHmVXe6C4Fr5H9gYbERM1Ut2N02WYthTUrW2AzIu5BLX
LkGMlojU/0wiFccHHHj8FtLU3dvn3mRoOpuiHWUhzlR/fL2JBFKRfSKDmcwhVh42HyuWDPu80D5s
BI30iMgg8E+c/RMEjipoEqHlL/umUKWLvEBMMKKF0rLIHe9ssboJ99zoVjjeBW6vUW+5UIXupub+
uJ1NCOQEbe/3dq8xrcsRz4188oDJDHiQ7iYFXgXpHs/z37AO0X0ODXGNQteUbJWndq/S0cgELhAI
AtoD0NdLW7mr7MqPtDKrGg68COlkPKccJQHlBwahgThwzgmgh1zoFrH1k/LR6BOv2qWo1oRF1klZ
HI/FhIAEZvnTVVdK+fhbXMVP6/RHYmWLaJvAG/HkVgOsS71SF2S/UwwzUvKSjTVRZE+GU1LYapaq
Ge2i68crNDyOTn59j0yMkgH7l/FuiLwc4Ir+wMzFSy4/EYrJElWEsnJf7EhMkH58ei23IxtUT/6t
pSLrirmEEBPNzW4FSLBKOw532WY2wwj0hmPGp2HtM0/g2Oj/ee5PzvweY/eQHfpkvR9/eTMiwF1+
qqZHdUYQiLvJsjnpVuJFo34OqyFRv8Ub04EKc0Aif6lH7A4j65BRfrN9jv2LjQVEP83KRa6p4YNo
aH5CdRYTg6XqESIZLynAGfZsWKoaMiipOyAAgZ4ye9cQc02vlpRoFl3ogOsJ2/FZ9G8ShghgAn7h
ELlBWN6KnD2ICg8k5gQk1SN8LDCiYyHhj6AnNOZD57dpUswcFOIWxXo9HbpYWJb4JEtMkAEZ89lI
sdgxB0dSWYEdznJ5H1pUS51rztZTh/U9qTpmg1nHykAqWSNwK1MRXYPlh2rFOSvtjUcmfkhIX0WM
c4blBEs1A6phSHfqBXWmEjkWCVpFmOCjMhankCG9Np7BUMvn8ZuEiTCt48k6vMoeWHJ42XtG9vhb
qv9JICh+W+Q5UyJidY2a67V9GEYtQIxz5jo2k1OpnGE43ywwN2/d3KdB/d4iWm7xzQ2bEwTGsR3G
6JJRcL0MXebIvSJvG8MaVBXzdIrXf8PEmintYe7SPadIuE6ylnpAID76GG9Lo5CNtlrdkuOtr0k+
NyM8B3lmcesjAXeBiFvZkffH1m9CbuQKmQHLTLKqbL+CKWcM69kqrRn9LE/lNcMSsqF12SBUn0XM
pNHQB46Q/8z+hy4vedx75QwUocoU7PluP7YKFHu4YXnqd8VwQ89ygJVy4hN9I5+JzQ5Bxpv6TmJu
QIGrhlx1L2aZR4lfLigPnUWWGFbeVrsfuaa61eVJZ06qDIQNLtiysPuJkI5GmY7FqMEXiOlVVJy3
BB468n75BtcMFpVEeCdlRexFVK4Pmd2RgdbgTKBgd6NHJb8qQ8uwsoLi+IQenNyOYsgElsdX8Lmn
91/y/NVDvhMCd9hxVzlwlnrigTsLvCcAhYWJIAv9pQpKctw92UKwDCv6GhlmkwyZO0HQHlioOaLT
1MCHQYnqk9xpCaQLHqgH+qnwq2hCm5D2EElqbhk32NpOPVN33RUAjpgmCSJI1aokEW+8VV2xU0h6
aSjitY94MxmkPpukDDJUnc7PNANuHH5fDxYxDDNMHriLYwkFeHUFQ3je+uoSsFhyL9tUr//1yd84
Rm/I5aPhEO80awRYxMlolC5FjMfa3GEoMgZLdNQzw8ovrtb5AVWQhNSoqdeMt+OMIDhWe7t+DKJV
S06FiMDeQfEkldFkGU9BxvxL6BAzMdrFk/trbRUOPnMy73pcb8wPzcJJkrxosCgLp1QzOqbc4cpx
5etq0RocA/J/L6rTie9cfk8kUB57DNnd/mPuAMis8F/fOraJRLWQmAgJj/MO69c1wS93Jk3ty5Qh
sDjfVqMs0NdUD1CLPPsDgWJWMAn9nkublM7QUyYrs93R1CFPTlXujhHoBrBprogF8wtFK9xy42Iz
PDfcViF0puE176KfncoltV/ybWHaH0VPKhia5lj7PyuKXIBZU/5I71el49wvrEW4Cqi7f7nrRRd3
fedassVAmWbgHsKoYPBM9p2CwK8JDUCyfMlRTRtLVYNZMj63KmErjop0NNC+eftZMn1u3taUequF
CmPUx1Qj9nGVEigsGDWq1XEdixhApwidmwWXhlK/4klLSPtyBgohPCkuz41Asu7JPHYzm63Z4y8+
arxy3+o+U3SyhCRQjYfDLhE2UJ7EfPEt21NtFb7GYN7lQh33iAef2taL/M/g2789G09TtrERHmFA
rqP1Pqa5EurvBsOlo56liYL0cGeeB+5cjnXm5mtLf/pr8D5fCQLhLMKZ6kuFuOSPXGggTaBvfvKS
F+fST4z1XJ/vlrd7Yce7e4ar1cQpOlFsWBHtg1KgecAnyXljFd5bKBC7c4owIVL4g+TZr7X7xl3m
qoqxiyvCMbNm3/6I2hiEO1z4BWVC1LyeLdoW+sFHgXl5RrobmxCJoMTNWMfVoL62kAtVR9S/it0X
D91EtVXnIXadrGkprS00AP3qTTBiNATr22layTPrRe7/5PbtBq1ilI6GEx3afEOo816FqfoHoZsZ
3YuJFVIjA12ui59nQCJU8+EwhMvHX2Be8wPxIapR/oxVuRLJmctBZVNUSbcpw3CpzTP5PqxaRSCj
F587RJgueQKQGz7F1q0uKf1uGXZduztCzKJaJRoO/VW+EjoOyJjTHsK/+ULmfqCgseu1FfslhHft
S3C35qQ1cILqbgwtpKxMExuo3FLUFIqyU1KgnmphimEZV3BoRaIbOXf8PytTuT66OCPZGeaoi1qw
pCpEDshO6db8zglOW9lsqBWfZWiAifAVWTNe00N+o5O18MYRx3HXnuaeXsPv1Kp0Yx5osvWNV0UZ
2SqMC49MqNQoTvrk/iAvVZKlH5OtwwX4gzQwfRDIAtcJKcTysRUbrlKrh8O/WvVb80XWN1LahMU8
U0r7996giosgx/ZvjoHP9Chiw9YLxydU0inQqwqJIEMEAmnxBphGMW53qaeHlcTNYopBAB26kJYq
Gq0bREGp1sUelAsDpl7jZpegmcPQYveIUFYIAcRI/gWldqslnCgWqpxbQdO15EcNA0WQz8V/iE+5
DXtfBFnQP0aSpkXIKapJTDiZFwzxkiLKgx21E9KTzohYSHs4DicFSs6XC5QRazC1vv22e3EK1gJ9
QfzcKG6bvMOIzBfHyS9K9QQx7oPnXukXaZc+u3jn1t9NH8vGxESBxIcZX9gavDpogFC35pUUFuuR
XXapkWCWZL/VYshXILs3gIgZnY3/h/X2PS7AFX2wNefRGpKZlWPqVbfnBOxJEXdfsDuVhNlodY/N
dDnvSWobHcR6cVdqet3rrVHhuSVwcz/inNE4pthKDpqDthY/4lrqKCx/s1nEn9cwaKlDCr2zwqhS
s6nhgi+JdTB013r30VgLzyw0osPsYJgB0Rxfh/AvqKDeJZXqt0Z8W8Togc2Guu/Czm1GNC0xYMZk
1I8CG2rM6glYLzXnkbpnFdZpydPodL7dlGXYp+LuBi6TGJJxwZOeTKmpIi8FwawMAPsRxgrqX+By
GDL6RAL8zaq5xYAjjpErVeeAnPFM3bR+ZOoAijFvFCyZwnEiHV/nbP7cwS1Bf7wclOjWMAH/zdS1
0oUFQKEfXjnUV+2mW7DGgJSNz5RHMsc0AijwpDNqzRXVa7w7bCPGDU9rKrXp/dK+c/vzZLDUZPiH
T2VmSPgeagT/fM9brgWoGjRYtT/1VK5J3La4AaT25mkqQLeaYtav/KnjhP6YajdpRXcVq+OdEpA0
y3pZqvygKAcn1NPhGaUrC26p9DLo9QFfe2TPnbh3KViPlaWo+6gqOl6wIZ+7rTNFCdy6QrzVfx8Q
h1lQPUE2pmv/uTu9oWQT2FB2tRUHLGuAMvt9N4ZtOr0b3SJTb9Dqe3QUR2aHAIHxWB4qVTMSR1Tp
2niq6msu9Vvn8vONq2yuO1fZZvxIdNtj62QWJKheiGbab1EqbfMGZ5aPm+4EdrPImn1khR3IUzlO
XHFVrmucOLjceJV055XblIp3br8OXR9ggSMnji5b2q/g82wzgJEQnENGoSdRk54M6nesMgzfXrte
0AZehyhn3KcQPpwqkUC5ntKBKLM63a8P2kclED2wkAioIw/rOhrCJn2B3NXAMEQbnmj50GVt/lTa
OiHAkcohN0iy4Y8MN60W8zSFEHG52CP7y3a/trQj8JRnCPCIC1b3MYQX4eLEOgUvWG1YQubYJIMI
4f5FpDF4WdF21SwN711r4XcZJwkUqMyDgcQG/edtA9Wos2b7YGF9TdDmu6kPnsXCCLH3RQ9nQUfA
TYCmYomEfWDdXaMMjWVbLenQI0rjKUzuAiF3Oy9C4Ubejo4VkcQTzo5AGWlENJltby3x3Tv9zy3h
WCSaZh382FiMrXjllRS1EPChuBT3oLwZ/9LMLl6MjdR87LbIPubl5oc44mjMlecTiarACy83Y7dY
C7shQjsh/A9txdVTvJRS3zX5IBlSTuPmQ4N1+MKG2UgQMkJCI0CtkR8scJkPmge/SOn3rKHyMxOB
q8QGTDxaq8BdM3FqRrQ9+SuZzecGjX3wmHgzMgfmQU9fEvQzLBfZ82gbGHzZROIJePSZbAOFzzfQ
cvIcSDNqa8c3XHEpOGO+42YrCIwr5kJcRTuNJNBxYyhovSHt4Ye5X9TGZGVaKuktnUfhy9xcgjEF
wOpHzy+dCExT++9s5ngt0dtQPDXbcsZ3BQvjaR9RY/3XYAaG914vbgZTEARzurlrD34mMvHmj68Q
ktLrWScyetyVSYOaoNICapPpf2WWoM8Cf3NVNuuRO0emckVUYKTB+g58LCLCFEgerGLZrigkWWok
2pk40ChHoXz8CStRXRQxZBcCjPu/Sc5RxHafDHGMLkVtXka18WhS1uE3L6QoziF7Afc1/xArEAnF
ARdW6P9jgRZNzr7XuylrjBIBCiIIiqudz35hWCxhusXrTBC3LF6ydE6ftX15X1+N6emo/6V4FPQE
km71SBfI6lAbbdYEB3Ptssx2bRpeVCIMbroIKCDVPLk/NKq7cH3hg7sIAuV9sRash6eB7R0dEeHe
L/EXQ+AxdAp7hEsH3uwFxnYIJO7Lt6GrHTLn3APk6jWFsTK1ZRZdXzVeWEMa4mP3o3Nvl1CN+/xL
nx8+/44LHAfK9xg/sf8Szo5QMjRGet/9mdDcpBA3yrovk4mH+d45P8itti4+/9fzQZIpgt3utgDo
FVHcbH3bSeU52fQ5yctxmqKZZuGbxONhTPgFjso1Lkd7B16XJSIsYIwzbbR4Ps6SpOXkxFU3vDWP
z3jkPDZtCOcjosyRH0oCMZIfetFepMad4ocU8QQ+j5yXKkK72UpREdIjWUij4tZTmfV2Rdo/4/cd
YYHGPVZSnwAmqV8OS77fzwoA/1q7zyF27UinY6rrO3aqk+IyCxHs+R82fwKPfN+xgkxDCDodrhB5
WLlkxIfgiZBmx3a0DPba4o7sw8Pl22r/euqFQihlReSg8paR8rzb600vH1LFPGIXXOD8YXvGPiRk
WYtmjS+qWicKsnVjRcgGSJ5g0RtsCK6OtnvgZoMDG8RLtNuE+jCCPEi2zrNSC1oIk+jFrHxuSaa6
Lv46nalJL7q7f9raKaQ4GRCab4ZpinJXMBaygwumKyaDbu0b5ndcWDl/xwmfq82y/ehBN90/CA7Y
imXMduxBQCDFjbEJWu1hbq7p/pbltmUx+h+iPa8Rn58ciSMSaS3I2DIHIBkpS2u0gmVBj4NRMuu4
b+BaY6+MMtdMAclTQ0U+C6vyRB5ktk+65GS1d4KHPY9jwUoEg7xLjrjxAd8FJl0DWATk5/+YC/FX
yqPVj2vGE/HDjWtVKLh63+MG9Xf0T6UMWcGudutak/GkOQv1xR3zzSziliLeO+L5j/XhKdb0d3hb
MwTiV5FxjY2P9q3wJktQPYqSY67Bn8UjaTzZ6HlQU/V76nQpF2Qd850eLkkTGX1CvRNC6tL9Kz7t
HJFaWAqA2Q1kC9ZTkRnUV+PgZkiCWEerFD5DvGpwHZj8+4Sv7tDD5tzbk0l00ArUWm3frTCSMcDf
CIdCGoNyOqOakB9EahukPDe0ItMSiqkr0N+thaOCVG84VV5TFNsORI5BUFJzuLBGaquy6gGkeRdQ
BP5HotyL0a3KxDaX1SMWhtWqEmsHYSiC+DHLncIPMr7DNewj9EJu/TN1QVi1kMt/OQi64Ux8eFyk
Elsb2jOdwCLgxlc8hsblczglzuxjaDDWimF6dZYTXFyba92K4HRc3YhprC2YjsTUsx3BrIwrbqHl
RQKK0/XaGb1AlxyNn/+Ku/CizLqozHGvLB5wMn/hvOvpQhckKuhXtBqfT7vsAjYlOVbCkzMFn/wF
wfRp7EUsrYAH/0O/GO3GmUggawvwI9aJ5fHCHGg5MPKjOc3ByV35WL8O0XEA/b3V3koXBmWX4grr
PAEkvR4HYhP0YQHkZ+9QSQHXpCy2lyQT2vohPmDIqxIBN4R6UCp6r1CwLQKglkw8LGE7dXA6TMEw
5DrnKnDvA2UCse34fH1NHYhm5bSWXBvi6HstO4qUuUxGJs2sDqubviyqoZlmKmC5bIxfJPmJTSkc
QfJJ6SvjdJblP7XGsZ8KsSMLKfbYPla3P3Ix4UUbIbv1mEQGfxGpR8U7wRw7sDU7XU0PIk06GhSN
eM1A1ALXi6sVahRNOT7/gBSTwAR+78rJ91YOB3DzT+bOVk9agwFi0aTSCruvida8yQxlEvuYeN99
aS4GHucBPyJjhlntYsJy9ovlid3WKdYOtSZxLhkX/g/Rfyr17TUBsQCf3HDxsiOqFW/yNg0LtP1k
IBzRF66nISQDKqnQ4TTBx4Susf6SQcjc8j4UnnUuHjmo9BwiK4ZQzW2PgpPb3bdpn+d0YLlphVXi
ZbryCuV46GUPe5pgTAI8beBPtj3N3KQ/agDtCYPV0bBiZ4fhanLKXQnaelFcIdPHlTVTmc/gnN1N
RMPD4ffywhgcBWE3iTc2atax8RQBl0bU3P7WEcQGrCPKTfFZmZmHm4KcOhEYPlxrXO4YKWA2Zvpp
ESM+FxdcpOFOnzoziWSwmKewiH/CfNwJoKUT/60dmIEJmUvPYfimS81UTQTDs0T2+melLtS1jOD6
b+lc5u/LyCye6yF4mG6Cb5ssQNAz3uYwiJe32agAt+f1e/vR3QTB92wxv8jjjLovV7F7eKQ6ZEbB
2cC7Ex04/dcHz8xAhGAcF9pOB0wtZIenP34pa05c1+j7lY8uUF6N29GJOCVkW5d2yitx9r+b6gX6
vGE/ELxbSazg4konnkyXcplfvyGR45I/BOKbzdd6/xWcqpaQU+2ScZ+A1BJ38j0aIKDjBzQwA762
pcpxGW2bmV2gIn4fOIeCvXmI2nClCVMdjwqylU0l8gzbeTpaByo+KiIf6uqrMdfKl18Id9g2mq/j
k3lq8IpkFjkIkFt6fr+qipibkMArzCAmq/0JAW5uMMZWGMHDrM83TC7VKIMod8gbXyPZBIErJczR
JLAeMqW9XYnH7+At3bJwNw9V3hLyuOp2KW7MnxVwA0niPiV8+wF3Z1nRv+gZV20JeaFgFafiJWtJ
Ry59aU9uNCTGR23mLhK4YzF5WH0fX8RcWGQB1qkaS19rfNp94MKjFTcNP3GzK9xpYv/ROCovMV3C
JoL6yXcH7BxO7tGp8shC8KLP9FfAIk8HTXXMkx7CUvfz7cjKke9xY+oN9Fr3l9YxjInlI/0qvj1j
ZF5FeM+Y4mgJ2X5lUMaR2Wd3whTer6araBsA6P/KjLUgcr9dhoSN77Vs15gMCveSiccxJOp6vp4o
J0o5Y+LqOzjh6myiEPGtRimzZSfUOcTsmtat84KkVpnTLEtXgIfRazgH6waKWvXhkL+VxzkENyGZ
FC+4YicCcEMRa2sig4fUX2openRHBpspoU0UvYROZig5GP7wh2YKdJJuWhN34fxm8gvpp+efnJd7
RntTz5Ox3qjYQR54eRqfLTYySDPo8s9zpAJnL4xdnQHjILfmw+2+MMwHWUnwdS4Tto32QonMUXGu
OwdV/TFt15lufSvCDplk9Vp4JclEuvX57Ivn02KOznxV1kVh5/Nh/Y2JgJyzmOJBbRYBjysMwaLj
KYRMVF8NdWtS0uLVxrF26h3Ckvxi2MT/+TivpfZsegjIdhcljZG+mh0rvWkhQSeppv0RRVneFS5S
viBsNUfVZtf23LXLMwK/nx0byqGuXGpBOJO5V/Mkq13pDssj/xWHTS2VgU9EkNysHgi5Q8Q1ci+V
KiVV3ob8OCKsNQoYDzdGrhqxAuGmXADpFd7Uii8hmiZqLKdx81i5Dj2PCmO50bjILJRoUXL8hcNe
cjJGVMkhm0O6jGwrXxvrBXk6tJuix+WZaJ6BZCAwnVlF1oIdGLRp8dLOipyM72U/rOlgJ4VNl6eI
z5qcPi4FBdlufZDa0QVxFITwzIjxIxzkqykqK7RpKWRZ3c1xDyvq8nWIHPiT4kYeao8s8JjZJyGk
GOhCQnRIY+HQYZCtOBGLgzfIPzv5MtPpQTHBoZkpfMg69r7NSB2sOc4GNhg7wpCC8cGc9mYi/T73
W7hMLNvydeoXjc0ywsnkr497ryYf6QfRQYZEZK77nP8WwqGVcyWYS9VFpaR5PcbVpJTdmsK/MlZ6
lMIp00G5YCPhREa2CmKLVlTxqlMko+ShxKBzpPCIXi/MTikYejhJqQB+MFVqF01/K/jDQ7xMEki2
G288nMbsgPiBDE91eU8TqBzjvhQYF829RLMbKA9wIa4IvL2pak4FjPv/M+gDU8oy0EQPShSlg+6e
/hMUjUkVB3wUT/mrlGcFntmc9y72j1BbEMCdqvntXewMykkJ51fesXOYdjjWxDxbyRijnsJu7Mib
+XQMYcLh/xPN1aKBjei6zym+Qdy5qUBwRl8KqsxTMPD0P4ktezudJA4ygdYrz7I4yD06vnT2u1T3
XQ/euSaqNGJ8RBALbFB6uWQGhKbNOz/tTCG1k23f+enh7V9le3ItW7QXNeahV05QNYDNUNSdjOro
b+Ova43xbRgRNK9yHKYUBJBZNnOx9+Sv6fuBU8lDzJVaSBiWaeMBdC8Eyolz5j4TA21sVSct5td4
istr9TPOmQW6Ly00MauhZkcKnARAVuLAwquT6TMp6Yil71kSnZ3UyYEEHVIN2jFtevg22oiULFhz
IaRKdrmi9c0UPZJXiAlWEjaNiEsepziURkgcJm/o2cPRWLuxzdD9LdqgH76AigE4diFDzgZgPjWR
Eqiz68TbvDHYkGZq46O1xV1UxItdu1jRfv2rI2lSvUBnNmtP2QxzWLGpLsqNWyK8FBbfPnIP2TzY
U9/OExyfs8sLXxWD4lMxda20yFnS8VaKWDfBXWqAQ2fb18KkriUq08FL0Cxdbk9/pt3xCECO4liy
6mKR2tz9UvHjGVvCgTDa3fDmTHJQeX/PcFVh6arQozIjiUoBXashH2GD5xzVGvBqOYdaanwYk7Sw
eYQnjsw6ySsWPSnIzT1o3IZjGWbZaZ1tipacwFytf6KvARdAEq7XeFYXbmoZJ3kIe83R44jK8eAU
2wLXniEMqniqcIc5iCbmBy0DXJ/fB94u1b04es0moj2yohzoTFWZGwy8kH17Nog/yEXST5gjNymW
DJzuSPbgjPnB89rlugSmyIBDDKamRdplFV1UKNQneKRNkaEULt6CjgkrDyRr5hA4p2VNsOzXx750
al2YvcDpAOKwtDbY8u2Ez4GBiZqCcx9a2gO+jNLhVxnIrmpE44DTLpmGDcPthHVIoSYpHDQCwOLB
yWSjPikR2WPjpXe2rmYYYPE5SpHUCsAg/yn7NvgGqOLUdrchcAzF+VZ8OKIKqLp9zsTHwZrrn1L0
WAugIox26OG+b1zlroNweFK+I+aOvSmNgh4xcBKcMVSGJziNie+dlNTRcOhgN2ikY8JGEfNlCJr2
Plud4LRbonmus4T+RJdVLsdcl+WOK3WXPymfu9wFrLMpxXUyShtpsze1VKvUREZIPAvDlFzhBqFC
H3Chs0BF8tx6BGSzHxEEYZ1B9ZGFhTVzhBPf03moXBhsd8pbT6WyX/0Q/hjJeWdcZpFBQX8TkmTl
m4H/aK07UgNWBg7d0TsJWJTLQ8sWWk/P1gU/o9uz+1wXnxnTHHTT2kHVNG3+/71qLY1L8/Srvu3K
C1wWOfl+WhQQA9jHH7K1CJLUbxXHhSefBzpNY0AEAbRuDPhNpdUR9mH46ZN8FktxaM+O68gWsPfX
Rc0vnmemyCcXEDvUmLwibEeGMBY0kqZlTAhHcGhhrJFJMvHk1izsl4c2RXxDdjQQhvkiwfyY+YsQ
ibHO+nhM+OWPLH4ou2dBMqYfqmBb+84gUdLQhDXGQPvrMdf2aAbw3ewKItZlnMexu7RDmahZRUdM
H0Rcp82wdY+LgbtJtyV6bJd3FaDDfxvznUUQza//W1itCV49EHOdSY+yG9IxduoaYqVWbHWg1sF7
jGjtbIT22rBc+l5yCKYauio8TUNK1NpySdXKDSxiRamybz1FAPN9Hrv4aUaDtNTkRsTlVk+/JtLw
jrFiahjdLndD4Z3s1lwFGprpITWylcPptqlNOVSGgbqLEX/Npg6y+EVaFHCizm1WXAku8H0oMRwL
hn736kINuKu4kya7PH0GpCm26E8AFjPlRxZlRlIHIP5TX6Tpe0RprOY8Kg2TkBvs72tQ4q/ut95O
geZ1W+BGJQLV/brK5/TWIkiKnx99c3NcOV3YTY8peghiMmgUYMjbCmZz/9SnIgAN1LGY/mwlgJZ4
LTiNpFIfBi532zaF89j8m/KlkFj24cqyPrVYQ5GUGGRZEl2Gn/HpyyKnF7EnnVaNzaCM1S6xlrWM
1aDovZVcR0XSKMgKrs296ZIzr16o7M/tuiFz5ePNLs7G8943rCx4YHvdmpDUIboFzUob7JVqkp4l
YVEzLoFK0eg94AlNaHM0fa1+RyVyl8LJauTKi84nlb5fsSVyW4+619j9UoXQ+HciC0UB4EJtiVbQ
OrQRFlcfmyEronoaSgN+7rIr5w1ut55KGObM0Vp3aNb0+TDcz71Qqy2ye+hOCMpu5XKCIfy+RydS
daYFClmUNH04w2aJPIe9xMHpdnopXeechXM8NzhVMXUAinJYjTfS4yoZphAIZhVvwcwIPiLDLo7Y
KSONsgCNMCqs5kA59ggVNUFbmonzweHyKGhMLcAiyswLlhpT1vO+4rhTcjzy1TZX+2VFy83fsad4
iQl674JAa0/s76CH+Sadwc+NdcVjrznHzKcJzlACCK0/AO8iee99rZ6qCX5+caC4+M521l0xSc79
a569NyLJH2d0N0Oj2cKyGjs8XgBiNNfQlKDvjlRwkBdcsbFaXK4c6nvwPsTzBVP699DLhL860vXs
NJiBcqq468DAunBh3wcmcFHYegbOL79pbI9tywcF+jMC9pXggneuJSrz9mDX4gSyJ7gW0jgy+UkZ
HldUPZYgaRoc1LGD/rDFO8nAaTRhsgne8W5VOmXq5Wolmxrvg7TIBPQ3THCH1H8x8D6QePO2/RA5
YPwIQToZbS87pbcb3+z/uPoFTdvvO1Ri/LQtwFj6WQyHHhjZytZ+ekvWbplgy14i0GIJK/2rPNyf
TvrDp9KqRbT3vxDyb7VALEmZ20JVMjlqrKOdmqLqOlVEzGztMbmiNcrA17iCRE0hKM/6W/THjcot
KMZ3h0l6jsgIzbRX8D+maIvOP4hDtvQsMJm7EcdIix82YXElP+OrIa609/71YNvXVenkDm54gMs7
KYMFOuwKGcW6wm9fW1kIXTzT7t0DK+AV26s5hkMeXE7Sq2F21X19KbWuhdYqFRUrqFJEd3iLC8+P
2010/Xlq9c1isArWij9Khd0SHhQXLwg2k5/XiQavyAupoWK4mKQmV/CoivV1IyqAkvjK1tyRLSYN
EeEaZd+NeA/y4E8RXxPM/nLCHDhg5cObrcpFV71QTUb7fx9CaWkARWTGZ39TbmnCIkDQbX0k3fbY
ojsBUQwPYK6edxmiqbRG6nKpcWEJUS9wwd9Adp9AoUzuO+xuU+C4VhNCk8ZJvyptRgrEECJucxQL
pR5thxZcSSIQwCad8rCHXd56nAc08EgqXJ6Xg9Um7gBXepQgcXIGFgZAxMC4f/14OXG8d1umWlB0
OMRdeIjq7B+JyuQpWGM+PUSWXo3R64KPZXYKnwj9nPBJvNCYQGgsQD/k18mZnIr4oY6zs495wGAw
MvWvGQ39s4Kad58Re72WNnfgcU8aJZj1mm0gsK1n7DppV1gnW9SMhPAWAPI721TsICB56JvJSuNp
KrRWrsIB1VKUWVpMSBZybzuRTi0oKZOyo+RjBNs8uKQww4G4/fDpU1fLeH/H81DFaW7XbWkdeUI9
T8R+NFSyy7sz7wx8trxwn5Dl6cqYmpo6RYkPJb+94Whm52+CvcyBPBWNfXZOi/zIbnTsm7rfB3Qu
V2Oz54TCFoqjPxvCWNnX62rgXgtLx6TfI12WOI19g4OP4xAvuD/yQzRPCN/HiIj46oUo/A2Prp02
dCnjY8ijw78YdEx7cEWG6rjscI9dvQHX4OO4pWRfC41OyjbyX7N1hknmgOIlYzO1AITWjh8ISCIW
POfJpVaY/LOglqsnU53BNvSZi7r6lQH++YNr98W5yZVYwucLLoSwuy/yUoFZ6mzhhyvmsjrmnu9B
Qxb/68+BCmADzL/IT9/CRmmEXUz2pSnFKd/eAN7yO+PtUNjrARMim8rMHQnqFLBe0qQJxZ3j6TbL
oiSFNHSUGhSBhJsBeqnPkguzgu9luJvdttM0CUARkxv3yvVc6o1fzO8ZtX3CxxNSr5lGqckNInLy
BBzYxk/3Znxzip5DAFofyw7mkgHAq1AMR/TIsGC4SCAnQptot1jpfoyYBctU5kM2RdHfdPMylox5
fBZSoNR8jqknwB4qDvb5nj+OaeUcimRlRrRsOBpyxpFTqdX+p+v8HfjMPYsrqrpeoOdzrovGubnR
Sn6dWqlw0zNdFH+Qk5D5946W7Z9WaLY4/WU+ZK9Ep/IZQcV+O1yAoGr+KGKrslE54uDS2Etfodqb
7jhO1jjKNOfr2mVZpIajNsCq1JJyyBDM1iSebiWXQqzoik5xAqq3+ezh2+/mVK/xLvM+SwISMZEO
Q90LfEDxBeLhq7td8f7MMkUbN39BByUrkErYjAqCMy7xWV90PstKkG8uFeMeGLRh61QCybK2vzCX
CNbJJBc6n7CrYacyUCtZI2RbrmspPCKanqfHmfnqPVZffgFGSiV8x5NU7NR1p7p4mDYo9Z5rOkEj
z0gZlwtyZHSZ6UpYFocncsee3ImsL3tXzAdBjpEBmSCD8VrZ80ACh0Bnt1813sT/fOxCk2HW4Yr1
1WQEHeoiiVnYmW2HgOSahm9NqTDGCJZOMQw7WNy0q0nmbEbzwjiszoXtWf2S5RqC8+cWpamIEPS9
BC/6yZA2eCXERVdIQFdClkGNYJvEQYbKflZ9T9UwcalHNoXD0YerSCcXp7jyIdiGh2tFGblUBTqg
e3tcrZ7e+KmWdKgM+/OwtZzDGL8Kp6lVP+aAePg41QRTgwhFTanWlsuNP6uPkCNWcsqcE4DfWQFD
oy29Uy1slqPhXvBBajKPy3Dae0HuN3PlBoasKCNLZ+9j7cVwfNzzgtk2BzwzbMXzpOnn0qPuxyJE
47fz0OCs2K92j6kKyceln+PT3ZhkYpgnGB3O8UzcUzULc1XkCeUM9yDg1MoPaTapWRLWJNYsL0yh
tMxzq5yYppEDfGb/w8J+DMq7p4pntm/oi9wx+21VTuuEGOe9uwEorj2yKYlju6nwASnBAt5yZOJr
Zwpqe5gFpce9DJYtxfDuLBfsvlUtKy9n16P5T7CkHu7EDzWt85cWRqn8ZSufjCf76WTKHbFtWsSm
EPuQqzVKm5oJffkKcMyG3I5nAraMVpqlZ8WX+eZpB6U7L50wj5VOAhLlo/XRyjBrrRuJFlOuB6Ha
7S9lpeRX73I7JH99a0XViJgCnsZjg/9MxzppHDiEoKZN2qppa81lvWQtMLuEu0jeaF2pIodL8ueW
7LQJAAVm7xr0e3EC03rU6cfs8XaXrBY5BxZziGi7SDD5PF+WLdSSd+/R617V2HUr+KG8kZOhjgFA
IG9p9spD5dpL+6Pcmh/3Q7u63XZeDjwcQYQW5Y1ad6TqnhrLrRfE7E+TXAmvUjMC44apIqpGQlCh
kqhZbSKA3ZBoGkgLnWmnW1m6hng5VryCMdK9qF92eAOzo8elPVp+wH3QDTFWarJBWFbgzDBSbLMK
YKSLw/V+YfY0QZK9xFnCJnHPodqzU2Ij86bnesU5B2rSV5/YCZuCFjyxyTCNPYynvIrnBZuYt3H7
Xwh5fwDl8uxI4DIABZthkyEFMiysLrGqD4MS4pMb7Z+txdGEz07YyHDH97OXtzRqt+yif5XNz5xN
QUT+aMhab7kHuIwuRUWJ3O5K+l9PqN/NSvoVaxb9V2gEW4eVgnrnEVA/fGj7uazZKZoUrtVAPUOr
EFlL+0CX4h0Gdo41urld+WACptSqtOHTvZjjD1rP167LlB01XIB6vNdXHhWpYBc2TfT6BUdmEZwd
PaAA1RO5lmzVNLrPiC144v+d6T29ghq8yxaB3x1uVRLUVGEhqO7oxTGYHe0pGTkkwrnWUrTMuBzX
jmgBUVenTI37xNSSkISFO6i5vsGWEvSPfJ9zYQIaO5gS4T6kJFf3kidpxe052Sf7hz7rc2XgZ2ZT
091rBtrAAhCuM0PheoIpRhg8Q+YUB6448rBCaWg5ChA4PHvGpfNXK/ZyyPL+Wp2Qs30KKd/r3sUY
KyyuXpSHssAXfrFmTHRByffag+Sq1xzwe7MaddgyojDyGieMh1B0MrN29SGCnvjSArwGI785RpeW
wm0gv8MA2yF/ZW/J6+hHaYTltdGJmQ579UZXMNO5en1z2uG5qfgtBaFMS0+Bt1CJOA/2ckYN1B/i
AG858bNZCmzgxPq9f31+mDjQP1nkUpRvkVB2QQzcLmTlJEYDQVn/DuOUAwBbLqg6B75Aj60ulsyQ
2/qQj5oKLaaIF0lmXFHmfSabPRORh9QBAiLV5gwunX7+ZPGyxM9mmmH+UyprEYvWsoGvx8acdxPm
YxyTZiFDhsHSS445/XA4xjr3vv22vS0uZmSc1ytjYE3uh502+5El7kq2gdbIDFYnLacqSL+Hme2A
8aEXLMCD4B0fvbypIogNu82Xp5EQkx+dEKxy7RCVfRkOLs16gBSvvYFCA00Ie6fq0G8/t6d+zEAu
y5LKo+nbvpy/LWAJdK1vvdvxpjXQQXau0Splf1ersCwTxTmtcMEIVhlt/5JIkCVukYLJZ2M2HPxi
cC8bnZobb71NLP8RsjFwU7+qTWMjrymgD4CWVEkEYFsNSv3RsOBUpS2Lsah7CqttZmXfa2wxe0VA
KM2odwYirxkFkXJbZm6rNW+ti2SyiBNMOYAIRyF2ve/UjCZGKROAiGGgmqOgXOS+NNbuC0vEKPiz
EvCZ4zfoPRWpSdPfUbF2sWMqEPFPC7qedUzJ9whsaRps5+eKvdaZP3iV7SgzrEzANXy040t9MCkB
B7qK38/OT+GTr/rcJyya4VNwlQ3aOKI1D6wIlUBgO/RRj7+dmK8QqdXvq14MCUOZwj+p7+S4Rzvq
S4hNefWzYfpunAoQBU6Jlwo+cR8NQZ6vGtxBG4V93ClvuE99pcDBb+ujmVxKjagI4/4aXH+Ts815
2HtAIrujXcylpqs97CJeMu1XJ8V/nD2piC/cR/y2WBuujHaVefIGO9O2VaJ4AFFl0itLV/8C5xZl
6M4kMyT1vZCFu0ghx5FbOUY+L5/hPUcdPxNiWcEZwFX6dKBtEfyCdwj4x4Hmh/wuDlZapDCQu4Rs
S0qfYpu63Bld970zC4tYnrKpI/lQ+DOXQVu9047tr48qegg0+P1sQ0BHWfgeaGcJBJxdvP6ZusK2
N9oRNvkQdGHQaFG65oLOrvC7PvoUzJ3qwcS4XlNnPhyU8WkTUYmvxW57bt9QSFggaGwyC5lc4SMG
lhWMPjjNI3wuJmBgItJOiOHvu9tjTBTOrJO6cGZYlBco8b67aPK3Gm9i5eD8Q1qTF1jcBn7xgwzI
w3x9G/SvNhB6fnx48548iSZmYUAWtKUODESB8AmvjG+mytY7Ol7U0giFiJgb5KYVxss+u/sfyqoZ
K4jJlss4qfkQjEc5Vj1gx52QvkrC3xI/fgF1tEUeo7g7jUkmCXo9xc5xbrgxYR8FDJCazFohiQhs
Huv/X/mR5F0OlzxrfC5nbA3ZSuXbTEgf14WfrCLxeocSnOdm2N1KvWf7Y0n1rnR5ine09zRRuyy5
m4+YtkOAGPdrDoMEUyq+FsPD7eQ5yuu0pk2M8137qJM5ISjLqB2GXVpFTVbhuEjNyx53GfF4ruul
zOjoYU9p+MOf5w5kuK4fcoBBTTtnYJcIka/A3zdkJ+aBTIzwS8uTy4TszABhy8Ckd6+rQLSiOts6
dptNhS30U6PPPw9nrJHafEl1vMR41aThmy4/PjY32x5n6QY1Djns9ZrqhGwJ97Ps/2b4kHlCWjlP
61HthdR/OgFlEDF3plv9bZ31lSpG72hpm51ObLG2DWkcicpock6kypXRp89ABGtqug4H9Y2lTTzi
m0f7Tt6Fy9c4Hka9sXeUKxNz7/IVyxe4ChQjigdpahqS5jQ7U5/VrQCxdYz5FPQSTexmEujL/e+W
Bd60uYKh2/FDnqsaJOcaZAgfU4gzq1+jC8oXgtvwqUgXd/RLpPZT7qI8+lb9dhhzX/65GwuJJkTx
QnQp+y9/nnZbdMrTOdEwmVpIJv2jp76adB/wcBSq0VuCqf/2TyGBYIZWDsjib4+eV8GaWfC7RO0J
kW3NZBR/8sWDF4pRD1Jj6IyMN4apWMHOQD9v++LqOrOCL5eGh4ndWndefqRsr3bQEn/F8gcfQBH3
+DnBLmWhNKVKVdPLxfBQ+HtBuqEHlgcrATXlRbuauzsFA+2bw9ZBOxJ1+XXXtuiSUzXV6tP2FSU9
ksesXmI47GySNMUpy0ZX8k3bA3dyRyw5gacsjmg+pYBGBD07DMqx6Hph5DGk8CXVjUb0gQjh5ps0
pnxtAHULoDvzsu8xufN7Wr4qdBY1r0zOdQZnbzu+2I3GjJlS0dB8I4Waoqbc4XqSRSQox//dDDe7
TH9SqswvyFimSu8tIq0XInBrrm6bJRferXAzEoM2ygYynryWpizT4QImqI+JyDsVkuYaBIaIkmpe
3dJjFXVOUAZttNXrvpHyzMaDiJCq9EYgwdIX/Mk48Bj1r876PqVNGtDjXRDC7ej2Gpb59etdt4fq
DNU67nXewy7hYxy/70OenDJiZ+qFWUO1Gx0ZilKsQprkFQO/sZeKE9xmqjUlU8OB37cXXKTDApEm
iukxSm+5v4oBVhi+5Z7Oc06aWZNegEiRjSq8w4JzfIpxyQ6J32qzyct6qBSJmVjl9yz5tbrSgn5F
Vq6NeHV6j3jSKrRnN2csB8gOPW4sZLDbXjc6MWAxucBTVM8L0NwgCAT2ftstjz7Inr7k3LRdIytc
dUpYj76JsPqyvqYWFYk5ylPmsYWeWktxn/+cA6FpYoM1CD3LchxREnqwV6oZTkyD1k+J3WH/40rq
UF6KWHnWitT/w2BG7CcSDm0PF9p2g/L5rwIqE6SmfubWxXn7gVXrnUjCS9009q9qOS7AD00lPo7k
WYJXLBGeb0SbTiSFvud1Pli7YC5m58jUTtRTtPIbCIsPz7U/p9vXZciatnB5vLF4cbTMOecarumd
bqqssDg9XP9rHXqP4mDCbNQuDv3qUxuE3nNBjVmWsN2n3sFK8WoQLg1CTAxhx+zBdwnHPDYXSEdZ
CIzv5GZhDVCskaANp4623br8coSXETEfsJoRxtOTRlrXs6FsG2q2Olaosjte+ZXSGvFpjMMOqOUJ
zL4Thk398kzXRxYFzTXMHorLUodd3milGXHYx97vJTJXSYjPscoaJY8vdJ2CKp4r3f+z3D6M2OcJ
zeGKb2P83YGVh+TcDO1YusPTTMutzd6bBbBBB1PYMZVeo6l5XbaGEkSkqZlS2JCal5oN1DzfyiB9
YRQyVh06cR6k5wHGTuTlkuMtKhqJR9LYr86BaT5oo2Rp3UyO13E+VkdiMtA6ytG6PnMcKITa0O75
rPdnTYzvCYWwd0jYMKSsc69m2OeqIAYwIXZZ71cIDGaOCufxEpKPXqsicnrLlJHQJtYLNCPdpdEw
1X4fRT7qqalPG5bPYmlugHxGxbVvGGMK/RDk5Iq0WJmE7MgSfLToWx8noRuk0nRPH5IY1vYBPeEz
wGWURo3m/w61gvWXUSjPBCPac1nbzWDwNqqKxXoNf9CuIFQ1YhKec+NXOx+Qd3CHhvzZ2hqVNlzS
fA0v/Jl6I3C68+PeWHEIjExbRS9hZ5lAMveV4Nps/gorrPPxT0DjI5aPznYlvv8FbiSfnzY/Lf9T
4S/HEZe/7l+phWv+S3XGiWOzKtJ9BfnNnEZ4wSSRMyadRXVGTFBBot08cos8ln21Q2txPeBeBy+I
Be6MeV1ZbUd/64KqzOAT0vJutFbiGqBB6GMW8+QZdkjr5hahx352jAGYT+/utOXJheQspd6sFJMK
t1yxf0j04OrB9Yg2fqxbGKWXC+n4ATuf9MTsTO9DG4o4uF0yzKX6Ve2IvBVg+NhAgQh+GRuSduas
x6ovOtEVfr/kOfxnYnz7/N21xodCo7feZO32jE6Aj9yBAPZYtCgvYhyzeVYK2zj+wEy94YA5X6oX
FBEYI/x5zs8nnLBlXkiEY6Nq/W4r+BAmGCQU4pEFVQ7ZMPuZDipT6JRc/WNVBGW2pjGiJFSgxwwI
Y5TQgV8BBoU/5znIh2iIjUjcT3Wl53Z1mjdswHrZeHjOG5v6h0rMVSyn6lKclygMhl8MCyv84ld3
nSR6eVyZsM5KxX8w5Q67wFqApEb5+ktr+NFdATYtMU/N88ZJm1iRDWou8HMsPm+ecMCGwaJBS7gj
KmJuHfFvxmQvcwD//7MQ4A2DZj4CfqxY8rR0Q4th0lQhzs1/J7suLBTedfCKB/IiZHZGstZ8olP/
Oo4BQ2FztqlLpLxQp5+i0RQg4Gb7+l9c5CUNjV4rFFhpOpWnU0ESFmRh7md+RHYIBQ9W2vbvGZLG
ffFJAbuWm9Bi4t5bcvtyHmKSt0V10DLwT+t4+pB9yfaNl4FWRhvXdr41lVJLFOSzPsqQpoXRPghT
4DuBBSmgy70RY1vUMw920zOPWLZUp23ualW6SvsdFLcrDoUDnctPBHIbLxSpq/DuItba9MnzLY0t
N5rCnnFtbMT0nr0xaoLCjxnO36YPs8bggHSLnpyUv8cNDq6ItjeiDMQsZmltRi0etyVBsrIxZRKG
TswGODrwU6gPGxnXHG9ALjq1y3KEXPO3kuPd4TYe2zXLDJ2kQpzXBBFvdLdMBMIep5zci02eKoNK
k0d2q2CyAdFDGCQbr/RVNhXaIpddnSmB+WVuM9/L75WN6DN01Lsvv5EFXWOthj/A3PLwAIyrYGWE
snm+M+a/nqox9wAe6aw6Fza5GUhlq1jlOvBPhPdMGliCibf4Gko2shprUZMLXhrZKAMhT+NhU5+C
w2/UdUQYl4TxMjDqCIq4pPh/QmjJ+4+2dR7oT5+njyNOgH4US7fKvXLAu5mfwkg09KyVW+XC9M4T
Yhf8uGpovyDb41w0TvLTOKEBNnHISjvKs23VoPjY7Now/kapfZ489qB+pRMVEBeSAhYzNZjBF4WU
bTNSbhuy2gXuQO4MSIm66kfUCSMDlvR/xEl7RAhTUlbwAB6dael+TyM7NIbWir8/l3R9yd1ZophC
VTkACeejsqJjNcN19bzzO5nuCs1tVCDhe4hAGBpetO0fmgTNayPV5Oe1b7823BpHe/yrdvYTAoqo
OyLLb6PBpmPUxnRdfG/kXrja3f91gItGsmJ2Fk94hUUjsbYIxQJqUmzcBjOEXIx8R25eYUe06UGA
tjwGEhA6d/f8dFw9GaZx9CHBTgeVDaCULNUA+L+Ah+QF0XrlsPWsMXDzUDOGuX27KtT79mfWixvt
92Tj1qOykyZO5AWIzBKAWH2abeHfjeKjhTlfAag5yER4FJCOViFJy0sZ5FCOd7M0Zm7coA8KEppo
I+wYonqB1K0YAF65P9ns1Yp7kz8c1MC9Wtt+0dYxtDLJvER7ccXzj//yv4VvRyKBFePaVFSbjYIN
dT7U7JOmX+ZyUp0OWylYaK0NDKI3Rq20POk0wpvWmwBe0OYC4/juu6pJLCo15zzMfstLJInWDtFd
I74woU0SWwcBV8buYUj/WZsfwGhW3w0ZzRpb0JOf8DsU1eG+6aeUK7DyQhamvg6EWODc8b2fboJo
8skfVIcIedaE2LMdvXw+QANpZ4j194FssZ+ylN/G7wx9q5UFoxYzoR+HCPpCp1swwgRZxF8RlrSW
+O3sa3zUWM30fNuTJQowuYw0uW7zoav4w6Y9GPKVGoYYt9GwoQEadxeCQxCHUgl9VU3xjhN4UIVP
GW9qYZ1vw0sJwC+e9L3Y1aWkyoPNOKw22HGlMMIAkkFjSN68u4juBkJchQqji3t5IP3uZnzQCuF9
nXoUbMl2wALdMOFhyJSzzvJXFEH5siQOAAeI6mXBOYvgw/Mqa4BBN7LBrQxStksDOiW9ePqbTiIw
mLIa3NEK8hMQE2R7afHl1jdvki+k2OsMTMFWNB/4yqosVCUfyvq7yHzuKpFYB3MV8ZeHfQpmxmtd
Eo8I+TWP8qOiobx0S9pXXM7JRSn91buaHsvWqh/hOx9LMpnytJFU3UzF8DWngqQy8ObrP3CLkyhB
fhUYsVw6PuhdM+8cv7CCWiD9r8MNAJ9WcVhJtfyCdA5AH/40MNmlkESzwUp7SEuVuh22DAdzhYDd
45M6PovBFOzHGdm55qQca7IsZCNvY0Gax3jGhWQ31A+0Gbf2NJBiERwlO+WK1j1lNwGOz9YJHhxA
7yyZK/5bdQxlLhgpE9lCBIAWJjre6tPnCV0YCfeJhlhKU13bjCV2xyWLIulB7tQfvVjSwTiL/3xe
CQVM0tRnQSLfvyqsZXuK60pdWtccZ4a4LfRso9chrB0u+nyzZaYuvL/hz9RceLrWdjmDKFrtNF94
8GSwLEynRhfUiwm0kMJTTidjf1JWxSl8bwu4gMgzS2a/LfVjKqcdynIFLhrcg0zIY5GZnerzss3g
GCLU0bM7KAlFApezYt3aPFU74t+70NTGJR+4pr2N91QhJgi8JiR+pBMC4gm212nQrNQhUbFX5Nya
TkeDV+6vAt+0N0HQljhWQTZVNE98H1d8m18UyOPYQBxFTj7E6HAarFdNXtv6lNJ0qP9bAo74q+cw
rc1zxdYsY5FYEDr5DXoDfCnclovD3vnsRlhjBUFi3287V+wD3pNaq4y14bSFC55oKagsSUOPR8e/
YyXWg6nL7iBBUYj28xuSrcZvevW30+Cm3sI+bvJCN2bf4sAzhbmB4wjM8GdTKrh5f1dIJs8dFkaq
hg0+BWiiEJZMdYTWKYqoYN2VLtulBjf9GlawnvNrAmtWThy1gAdsoYjQpUkC2Vr4s48lLkWOaUcy
6T4fiVitFO75yD67kd37fjSYFTLntCL5M+uJujGbU5JMJzyQV+wIkJ0CXmGiX556gp8pT58XAkY2
ftICiyy6Kz8yKA2RfaxFTiVqLFNNmRlvlz+cJb1SbSvI76ZRNMZBsmTos8CXPSuq4//BC0/eA34O
8EmUULX1p0XL893HLcruQ7wK/GJ6yYMQav+H8AJVFTXXPZ4fifrWVx5DdXDdQTDYrKD7az6OJnUJ
FiNNBozuLwzaRmNKia+33bYv/dwILXKV3DAnmAgGYom8eFGOK/Qx57MDFzEKCaSeBE2YRKPC2pq9
3Su1m4844lqZo1fO2inC/Oc5VZc2TJjDMmUT6GgM39SBNzWxufNt7uuUWFk4gMuwhCjealU71SYP
MJmWnbBHYSuZhjwemVaCQ3qQi39kyZlTZQ75CI0TX5ELmmlUiR1VS12wqgLcx+GBexCONwTy8qtf
676LGNJN2uNqFXQpPXM2HDd5ZBmGgxXmBfkY90KZ8VMqdohrTdQjqWCO+qPjFN3ihZI21O/V1Him
gcuZi34eocDekaLeBAOo7EHvJjDeOm92N54WKboTtx6tPyadkOvKo9IuTCrrMLQoa2E5DNEavVAX
9CPCnBBG+LWImf9dD8n0fSITf2V/onpyWfXeKX/TY3EQkZXTa7LjOv8mOn9YAyOnHSN8bG0MMJyd
YVssytQdIsHImra37WEVJhKfvSxlhgNS1X+8uLPn+OyFYmWviWxUKKBFPBv/XNs/P/yecABWZz3V
VqMys1Xp67v3vt63uyPrHCjJaUuAAgz3QpRK3RocumW2g/QCC3QJU7kiVpSiJdojeMzYg5xuopDf
XhVD8CXHGCwMfWvnP1z+JT3uN+GZBSQkmHMJFGTbiNmHak6m9IYqJokyMFjC1EIVCjvqZ7gZbaMM
Qt8aRQWY+JgMKBJfdxZuj50YhCF67DpTzmWjmDmP5SdJKqXgLVXugJ7U9dRbCRmJtRcOZnukw4HG
QC8SQVbUMmYAc4kkbCof+rIOB64ttjgSpmQPRXv29D17w2UQif2hOCmD6Il8Bvpvb8Qi54c1+cM6
sC/cuI1/4WZuylzNIIFH3ELVJhD81sj68vIToEA1IKP6FD9KeGzWAS2cqAJRPQVX3tIrwC0pcHXZ
an9dEz/C+lcvVqy4iMRVZ4qwuHsNhq7wBjuU96vbn1H+9d8+/S6agE9QpYbQVxabu+cLP9pgApOb
SR2IOLE0Ev21eX6mDOUtm2b25mgObklgBGw4JhONUpPzNBvCSW7W5vH1deUzsXhAlANqeaf12j4f
rVL2O5gPToe436ostAi4yvVE3h1ImYFlhSpQSwsdtl+D4EQ995Jx1s4uUqOHtiwvhCJYL8uoO5D/
D6hK53nawcKIXPPUHrfKDWmJIz990bqqdSnvHxmbs69hU0m8iXVY59dFBaWpT+TiHHSMxuBktRNO
mlU6+zBcUgMvkU0JrgMbBCDuZDHzUcz2jEklUWmKMv/eR/IpRF3HjzysYyChSk45Yh/cuAzyQINl
KXRMf69hRYh3bU61BRDJMJx88miRwj7rTrrgCpiHOiGS1U+htLSzMFBXBF1VNUwJ9jtlWDtsfCsO
sWD8xk9nHbKAcZfWwBmya78kuC1hflWSfid/yiQVBzd0+LzqLws4QqMc4uyx6v+LIjlWfBPjkby9
I2MhcXJV9VVUBugLcTyDKI6y9BmshNEt/AQf5UcyAQcINqkROdcBfcUTXVMhFA5GsRJBTdHf7rmT
c1uAeszkVBVrk/LaZ3NUwELf88fI4wTXRsJBXUq5Gt2fgv03hevP7rcRZpL0k1WlIX7RiwVdjWS/
jjnxgxjY6Iuh1KC+/E+SPA3QX+dLi09ZeWl2CoE2DorJs+9TLe1Fo5HrFMUXpa3KNZuyAe+ovhzq
hHyBkUNhvm5pvaoyMxwAzMQHNjPIvupIfLOC5efPpymqMgkmdyX0oX0BcxwpF0Mw5AqdXfbnEJGv
AtkdUGvtEDzacg7TeecUpfg9Qlwce+iWu4+j13GclV/R3niYMSdLotDu6FVOexRinn5SsrHS1Axy
24Y8p0tIxQSMxL71nrV8KSRjPi6V+d42r0uL7zEraY8eZ/LKGYyw6w7ylrY0sYKORdIkJygXDWe6
KzaMqRvcBkbSTmaENZAoeVD9fEg+vsorPrduGzCiqMZJ0LIuwU/z7c9OETt35ITDicks71mXwxW2
ZZ0eCL/x6ogTtvuGzCdFLru2wEaWTgddxv5M0mtsLK4WWxin0Juxx7nHx5XY2dVSL/hBijbKrix1
sWfUq6r0tqubgPfFoGihTEXXocYDR9ebHBS/s9NXW+tsVc50/1iD4dTFJNDSE9c4kxJNiyOkTGa+
Anadf1QbnO0uRofCN1efgMpQBH0gyAcExKNlNhi/JVJ88vqXjqpchhPtSFY28T+soQ5WwCsHHNTR
l2Qw+g+/PVesFrnZMXo9NGaPW6zVcTXXMs5ggMRUwm1QZWa9z5aY6SZ0ozrZ09XQljb/lcApq/2e
y+QoUj9cqbEW9L/tdZRpLR8w2FZEnCI1idDp3SQOe1PoKRF60HUEswkTB7yHmXWJ5pVrAM/p+zbe
ffN2EqAW1XFBwWglK0PMeOjMVlg9n+M/F9NxRyg2TUH8OnB5mXZzhL4PaScLEosTd3kfPu55oYoU
xUXYBTSs9S/Xe2K6S1xdWFhaHJR7Y1Uqybl4edUgPsvXrCnBkO2B+kkFZnLPl1elqFKe+ZfBk4qn
jLM5yPmfYA/ZMEdioEhGkzopNH+lDXvLETyKXG+gbl4EVliTx7K73FukSJ0JM7bwHoQCngrfh8Gu
ErsJ9NRyekTRgxg788n3xRrAcc9c3f41I8vbOvFx/HQpjTEihl9UufmnEoInc8btD0+Vw+gdthUI
uJDGSX0zWWRMsTcLmF+VgFbvIKThxVSmZAfKGcC75+8Uj+RLFBNGkq1fdAExYEQTiZMJAfaKeN5L
eSGCt+lES3otKxwjVQsOJsDHZc5R949E4JwJd5CK+HuJnTrnBolhNPjW6FmQ8Dx8rDefa7Ki8ker
+o1aWtNmrjJvc8f9uLGXqUvryudyzXy7QtHKuQ5VlEOeZUF8kNkTdhFNdHtRgGlTJuKegdNHsDQZ
muvXG0/6iN/gK1qxfc8ld2Kv5aX39a5bUDZaVC3Tm+9mEPIFKj3hJHpTq3uu0n3AZJIkM628u31w
N/nfwwJl6vWgAvoiWfYIgALbZIQKuEuuP3q/VZty/8aBr0We/a0EWQwG0wvsY/fVJDqdQNZRyWRd
I2CKsFz2DkVaTbjxV4WmMnXq2ELMUbYoia1eIBlNRLE4+qsM7AkEyhbFhfPORocNhdfpk3L5ZoK/
QQH8VlaN9OXrFmYLfoMPZeU+XlAE9eUUzsCy7aZPJMWJbwUyBdHFxIV3bvRXubxuvPZfk1PySA27
NZS7ou0Jy+80+5n52N6YTZnJnOXlkfLdp22S/VHR8U+IGYtWJn6Dn9iDlYMEOwxG7w7mnv524tuv
haIEWewYZwEGOodfYisZ9GOIVTHuQyrtUjjJanLRca/CtREtaBNsyR+SPeNKhgn4dPvoD0owiH/+
tkXn4ST10IqkGysmoMsZN/ixSyULdJOB/IOL7i7xVS0uzkKEuIoE4V/d97gPG3qnzBniiK3eI2rP
uB3zjiEpl6ByDLrqGyOR2tGEsfJlbsOzKGBMUknyd5ZCNUj/Ofz84thqm9oWtCBnzHL4LvgvcF2m
yG4CyTC8Z+9+/qlO5yvILLNf4Qx3SppOCfFC4TGMnox5EI8RBWendpNTGUks1D8fsUmjYisAd6r7
o8cfhECgFFAPR6hsQtjs5P7CYrMpIK8fLyxH7OabJLV1jXChG2c+LdJhGnCqYVV/J4IbBRVJDHAt
0IjL95ZB0ytXMDJ8V3m65M6kTv2Y36oF9Urf/hoDYWoGNUoq4BQXCBtjizZu0mWLLXnK+gcF+IXW
TjQj/ILh0JGzkbPM3IL06uT40aIxQWRgIenajW9OQSxDimEJfAbgfnsxi7SWqJiObeu12cTVNr6O
NyGRk06ai9qccjNJVZK7/noSss41IgKWmLny8ry9YNIl6Sn29caQmj8/dVN5CdzAnznekn4dQc/Y
utbJMatvfDrcYtC6iUeZUK5qFoJ5A79K02XIa3FMbWSztUDH/x4bwpeOoFYUokYANobuqCeQD+/g
pCmqFwlbDSfjUows0Dy2P5gdgaHHuhUDLV9DWIbd4+j3lcr5UpwvsD2zawVp6tB2LEnimfGG0g/O
WPACrikYo3WAWig4MsN6+9g9mAJXIvUkusyZMPLm2cvwWWeGGIUVEqyf5PMeoaBj0JETlsELY/1S
rRMtZ9WwOCDQhihiiJrtd8O4InETonCkqi4MyQ9lytvoeGDlZz4Q84wIv0sjAGGcVMvz3/m2DKv5
g/M5sRm1yeLgnFTSSYOwKBnHHqLwkfj282UhKyGqVjCfdik78/JaLuhgOUIrbeZpiNHJ8Rt/F3df
m/cbD/vKX9242J4EDk3RCgaqiXp0azVJ6ePukRhy/lTybPmU7YQyNcLDLW4y9bsjqj1ZWZUHfpLl
5RjgORu56ZEKYbj6T3jBhr6k2oj5SspdujNnoK99dIpCH5wna/7dIf4/AvXxdqeBVenfUy2/+tL6
ns0GS4vqfTMumnPELyZ+yHGy4ybB3hWBbSOLnqHNpWAPrJ2N0uYiozpnSCiksGgo7kXO62xckMhx
9fL4mvDZ0AgZu8icllcKKSnq34EZ3BSxPwOEf52lIo4c1GgMNUIWASRBhZEkQPDpl5ZXw7+SKUsj
iXojeHdzdW5uTqIixNs7g/653oUg09IuQ4yEZxk3cO5+Cmtd/5pGnElKrpi+gLVnWY0MgPXZjeGp
2czdv6BXeXJFwInIXr9tpr67d63SidCVaQqrEq+jsoIHULIn5aYUnRUXClWx02CuXXOfKdZMgHT5
ymu1TnurBgvO7UXv41nTzG+mUV55h++eu+xniKxUqJgKY3BSDQhJbUR6hgt8CI82K28ae9Qys9a8
a+NEI/5ugsRYIA6ZL7rZ1PppyDCZI9XsnJBBe5PFqhJ+00u5zenqBBrfkUAARo9HkjgQUmmz+ruI
s98XYQcMCU2cIQjjmsT8r0AD0M4cjSk8+OFXTdd5yl2VW/HJ3OAGIDBArPSQ08XVamZqs8P+dbWy
MLOhNEpMDoXDlC/JWhBQ9o0Mjekx8Mv/Y/zKsTxXYrQTwOnsx3gMhikNn93o3ismFc/rHRvYAz2P
V3+SzUnd96ZS+6avrHRnRwE7rX0qvQXVRoEE4zvv9mthke0I7xehrSrn3bdi5WG8ao2puLkKNLXg
EkGgtBu25Ek8XMKhQb2yT5OiGvSwK7ah0EF23dNitjXkbnPPMlJyPbZKiDjXdtqk1jMo6Ea2rKBD
fvcZFZ6ThCa5ZiuBNAGhO0PSib0mA9dW0vOiX+tSNZrTHw5fphyDpe8rP//Xy49a8wXJgvdXwack
T+HD/OdlzBcZoLdm0AgiXuVHWivqsRsd3CXI3KWfxYZSh9+TrC2PMtZ1HzNurSjdk4JbCQ/b+7Sh
a2uXqZuiFknJjoafPO3oan3R8ZmYorlkGi7/yms62MAjBEwjmuo+OeT1LHcj7z8gl/EyI2IPlCRn
pnCCSejlgf+lP48RfBGaH/dEJWxK6RVdnGpeL0wODaiNcC5PvBBT6e5pYRB7inimCtXR1fa9l0tB
T4LcFExzrKU41uLDOcI5RSIeQWpEhpRrWCnSo/nag90LNIb7tN3GOAIgbp6VRaJtTOvRGTi5wrGO
W7ZMYfkkJQ8e3g9Xb0FpwNUtHQpyUEJg3Db2G//BHTdL56ejpK0M4kJECwmhUheBu24DPHoD/shS
SOhu7a0E06E2wAaIC21xJpM1mLV4nFtA3+QkK8N1vyLllumshcyXxdpAd+/wRaPg4CbP0EhwdCxn
W846TVFiq/4tAENyeOgrouRaHrJDk2B4cmmxhA5miEthq8TEEVD0kgUcUrT05YN3Ky/fbGejEs/T
1A/48PtdeZa2EdLUJS6zspM174fRqksLEd/gOVVZwnabfzOOirdtD2Ob5cBnPnPR8012e4bpdu7f
h4SCNYQ09eHUuxIkP8tL5WpjHtwlA/oMTyFaQMFPfdF5ycfK/6dLBKieHCuDu+75JvLfisJrliNo
9OOQaXpipdATuzdBcBkj0BUPOXjIjcpPL2XjYUxMxjGlLinsiWtkQgHNsWRUzf8QnDMoQd2pakfz
rhyVKd/iRPMJzFtTDUX52Wcv8xRe1MA1B8mF67QfNobdbQRzkC56/YpafDXWlH1bd1XHt16rsW9R
B8bzg5sprZsdNPYgo+ft4Vfut+OQvvW0TwExNIFke0ZTSdNfxFgIw/y4rMygE+bfzePtpdlaW3Yd
PSFVsAZLgbO1uBBLR4ZvEaEp7YoJb3EglPjX/bhpSyWpPoH3RDWsnC27xKWng48HgfXWcV0Jjx1n
lHEv64u9NFM/Dp68ySfBslIfz1e2aKb5mGueFEnwW4jLTecBoytCLK6GVnBBCRKZsC/8XzBN8s2T
JPsqne4yp8m6Wcw9lNlap0qfU58RjsmrFPXJlf2k1ZrDoFreXrOZGL/10YUDCGiKwrI9IO4Vq4BV
DIFslWVEWzaxAqWOLnDaHSNLuUg+KoBVWyLUiO3E8YBIcF8llGPsVqmnDeXJmyeNi9I+ODj6m0EK
7L1jJtYZpe7gbi1lXdIGCUoEcnxk+Dv8w0bN0UiUe28SEM+lxW+8RGL6cmQ5leOMmYIRyVg8v4r9
9B8bvR7OJ+EFMIRGZZzlBb2KwUMxzmHJnGoa47/HTsEzC4qyEORC+HRqzAB6Ork0ZllyJWgcMSW9
xN/4VS9zu81UYUjnjwcrR1r2r8r9LVQ9ztkCVT7YH2X9XKJkNwbSeQaPbpY6J9DyxAMZ3EzltJEc
hXFn7LBieJ0VcjiPDVy+xfB6I+6EptcVvkPRJNB3O4A2p1GKk4mxu/kOcyFL0OQ7dfInvETbUAi8
c3u3eJGHPRgs/pEbKAOoRuKx86Bt0lXce6vnIlxRMjIv4xLS2j510AcDdF3GAtozkkPB24v4YCJ9
sPmx4SZF8E7AFwkB3L30MqvN5/dyBOI31vsvDceL6Qr9b8DIZMqwfJ+d14Fa6TPTkD4/fBMgo8c4
r8Bq8Na9ZTbdL9xd9/tt7TUPygEKSdvYUFjDSzCsbFBWfafQokjZG/eOTq2dbCHigUf5qga8/Feh
BMo748P2Th9e8L9iVuCiMQpKF6T9XhxaqRXGDaihJkn6pF/iEZ0qxdvbObv/qdJjoLCOW11Rz8c0
z07hQMLQIAI6P8JL9UY2jqf439JHHNGONiUKEpWJtGfNnfv39pP7m+eoQ5c0N6h6YpoGzLPrg9pQ
8MZUmU8nYByAsndsaOaz/SIzbl6bogQiXqNU8R8CSDKaeO7BsFfkpTyoAmNyXlLou9HsmlrPPPZZ
ysFdfxBehC8MOo7rvTjlaU8K4IrWw2TU//DEc3W49wVTCTPWhqtM5hXAaZojUtqrU9oI+w/oH1HR
6OflMWcjyYbCNZkwHon0EeXSQLnOcaHx9SZ0czx5VLtv7O+B2AZ3pZ6ix46ooGZTHYJ7afuKcMEo
B63Asz8A32sYw49aQ+ISTJ+dZ0W0dEs0Pl/Es0tB+Q88HjGt+t/J2/pC9zPvWsdca4Q+hiupRpOt
fFr3Pvq4yWE+emuTR1+lTkeBZWi2OGQ4KsMQhwrH2mx9QTRwrfoMFUidBUQb8sx6vNW11SeWT50Y
h/v82/p/OPsPWNXVHxBsUR+FlogjZnO6hVjLnfpfpzZLrx+9ziwpbWd90Cejxx/lPJdBfeUdVSem
Ls9cVVUlbILX8MVWmiHxUV1jX33tyHGluTdgAz+O3BtrTdS9kw1aOOJGw8JsmiZVj7cBxWBsOqdJ
KV3o8iAnYalEa5LGVVVpRDJ6heoLewwEZHDCf5JFJKpwx4V5jG1SKhGLzOceIPrOpQylG5W6bppG
a7aEPE8V/IWvvo/w0b++D8LBcrNwQB3/U37Ar39ymAPXbs+E4PT+hU0ctktparhKoKkmJhKHB1EQ
0tUyNyGuy2VlHNqGKPn/9B7lq3jlu+x9i1j6KBvpi06Ovg8EQ0cUy5mhcKMWSg9Wv+bkTQ37hwoc
1j4S5Hla1VP/a51k/a7BQTzlBFQ8wqmyydkDuXLXkb6fIrU1MsvRVvlZgvWfPVqcGaN7GHgzzlGU
EBuRzDbq36qBePmpMjbT+BXuZlobshVLxGy6IfZSCwelHGPjntwdmDP4Ma90TZYqLTdjDsu7Q52v
W6fJXQ3DWTfc5+WAldSo6CXmQ04SAZuZKkW9QrpyYLLeH8JwMmwBRLgxWqbKyzp/WQMtLQD2vZbI
HJnO140KbKIjXopVnEf18JAqbnwMd2IEIIlaD+GvE7eF6U2GHYqGEj5ZUz6gS1cIni1rz1cHPUhx
nywFJkS6OCz6YIGwtImVH/R/EPKy56/vogopht3nQ44I5GouMLUW3gJsLvBIHdEM3Fi3pNrhsV1g
RBGfzaRtyG+nSADq0zvXH1+WQNOd2l8KyCEeoqTaKnWcue3Sb5NbVtldT2QAa2JakTTXVqi/1Ycl
032SVyhu55wDO06+5fcPIBnOd5MNBM7cWJ3Tni9YO6T6jKeWoeMyvmLSdR9HePhL5VpSmljIHGzW
IbDHlCFSQWJPd8tcva8oB5vRXEkuDqHdb2SCaGIsYXpO1TzfWRS3JBbgwFdA1qh5wq6kHSLjcOuz
QwRfLjSpTwIF/U4bbuqsedkjWwiQtkj67zI4T2zWNnLQua/YSw7Pmo2HSTcs8DA71H5jxGAmhnA9
2H1qeQ24RRVOvmNIRTGRadt+qB2tlpS33DQ3Rob7S72XrSbGtwq0NJ+qiHq3ou3f2xX98c3q1rP3
4guaM1gzIqeEIDiw5Plo6U0cs5lvdw5Z974cd5ykRzZMwcruXCGO/6VVQQNDMYFkYu3Ilrmy9IMm
3JG2Ptyr5nSON9sTFWIXWHqhfufhhv/V2J2a1yN8bLW3+O5XjvwrJOdHkF/HqAsDe+a/NlukkbQ8
66Q6iB/pDHvfQg0aRLdNTM667x+Fx1hufAsqRL3KDmUd7ROAmZwLF7uNRq8SIypCy/+5HQPJwsCI
xJfnAsrhd9xfJWCnb2/eOhhLC5CrL9KV9v50QKzY9NaT40nt5YtBbAaVN3sQPC5CD52rFH1aBcad
b2evOPXNZSjugxb/HQhWmvsZYyORoqmbZQE2WiMTo2sh0o1mKdq0ZhokjDVuxkD565oi0BGdpcUc
AlTiFYAGLbV7K+xb6xyEHoLPqclctDRfxli3V/oQfg/F6jUoh4g1u/8PpN/bmBXmoTYqWtsX8bex
yZQGqkXMW+nm0CwfrDJ9j8m23YyZnnRRrci7wJ1Kv8JnOjaFixFvSDSBerAQ0rfANzTKTc6d49yc
f/10Yioal+4jOJbDHGeHz9tk4tPiuaRU/0v4VVseRamL1av6FcZNCxmPAYQyTMwHy0t/oemrECQ9
7ytgsBWVeeI7bAoyjgUFlTTMgmvrOYXaltpCelpaZj29aK22zRWiqQF+umw/mEM55gdFx8P89q3q
JzkOVgKQ+OBaj2RjJm7SjPgl2O1MSF/kwg4VdDPqRm829vQQ3ShcxMeyKJUmKa/YBH0tGVx2STLP
4LPG3r1SyygtmHD3DSsKXKofDB263sOoJjR/Klxjz+6+Vj1EXM8AAklFnTrcZADmk2bhAjezR1rL
uc/QqoUX0H6YzwaGgj2RppFEnbgM0mkLCyhdvbVpvAIxZByeBKu5nhSitUO/tc2aHI1+3fVRJIjR
9uKo4y0o8ankyUwke94hZivRu0SVMnDntZt340KXkbJf42AJeIpAZLXyndN/wd2MO/kPUfrKmlC5
dj3tL8ajFJ2Z7EP1axjIOK/3FDOLDqIVIm0be/5VfKz3UKS2qHSMEHw6X441du8I5FP74bwEslGg
IWXoEet73QfNRdwQRd+cQDV3EbNCUCP8oV7lOuYvEXnidkQKQHTeEYgB+bvYZWgpaKCW1Ey7buZk
/D2/PUfExOvZHJRdT3kDgv9dRL1IKpj7e0Q3c9YemrLgJX5fi2lOyd+FbRGXCAHFP7fCONY9iRCq
6KIGu6uY0W8RcJ5i+GtT+Nwobe31hD27BEqJFBmwF9M+4H/ly0l56MDHnkDR4tDiLcdYGNbP+yRn
+qF0S3ax4eVbrC77HxafmSXFyU5DNNqDZu4vvGv5vV+yXTRofQOmnJdFpohEtJoV3joeL2e4WOT+
Urqa+gMgwiNASofvI2EufmcQaThDbfy/Dn13XVGuyuMIIv9e2/XuJshCrfiE+aKETCse9B5Pznwp
E/z3fZ0huByoc2nuhZgy1JpYyGxK9YDLVQNP51SbDDf3wLGJoZeVmHjySLTxqdqmmPiRrBRUlVAL
kwTnZNGSS8gyOtsevNI6FkUv716+jzroyT9PoQmjshIXAU9cyVFtq8/SjD+SjNxyzGRiFlalaAbb
Gll7pyEiibl11hUfahIptzfC6PklXQoPWU1iB4OPiSYU1WCgA9jv34bIJ/355eTAlZuYZ6f+2U+F
JIL1RBKmNM4jIdJKwm0/VVDGi8GwWpBSlgue2M7WPQMBI8YevxhhMddv5OkTpiOZ506xloQZJrrg
rO3PYO1k3RCQ0Sy70qzGK1o3KGGh/+y+Bw+hZiJ32XlR72eygJRppuwGCxO+7HjkNvhd6Nh4lJZI
WrHo1HZGZjSgkvYxIPStiMXAfs8ISlX7kD6Dt8BP2AtD0qBG1GoF4zhdZFuRYpgmnQbYQm9RAsJo
goYfpjUiLniRSbTso0jNulMjdNRCmAKEWOTnG36Yqx33sYRFnZS+ZLpzcyq6gjZWN7gdnMIFX/UP
Z6dvqa3mmgmuNtsepU2lpTZyYYaF+Q/rbogA4kmb09AlyM9Tmi36VA7fwkiQRDnlqPyHb6mjqscD
uAwhd/+6mjpzbvXpRoYjrnOTseMEEqC2G39J/HzrLGVA+he7dg2BgiB5Byq/k/qLqYnCHVnKBNot
LIZt1ucrLUzQG+5yZ2ptOknDLsV9AoQKH+T/fdECA+TnMLQlMLb/7aDvvmHNG+OwOKy9tNY/rl7c
WZzPFqomA2ZTjiu9eLSrZ/LjAsmiB5GlVICgNhUFsA3XgoeZ/5VlUjPoCVHJgXgEbG8NdBHV2WJm
DquaBtjL7LvwSsbclIUILUzJLrrhhb8cxVbn0Xn/T4R4qrEeUBg/01JvrDmypjVDWfdbErd4FztM
ZotB/+N9SoSHotVrvyKGGUnMYI4g9hq3zRCrwXd9nXmJ+JoAyQjwDzl+RT9N/EQ82VURf7NQ9KLH
fGmSpD+Yh6NT94vaUb1y09an1EeG9h/i3vRmeQrRLJV+Fq0dN/tPFbio0l0VDPKJSNbSfVn3V/hW
+PIkNQKmFUxmB4PnJ/jaHCiW6s3AE7+6pUYpM5gafT0EcIuauDfyOU5rZDHECM3mbwOalLFTyg0l
ABYi0QQD4IX9wwZfmwlat5fty6iNgu1qbS/8Oftpg2obIJPycgZEcyGHt95cCwXIxR1F0dfCoaUK
OOMrO6m90Rr+O+AK/tOxGJeQDcBACMy+aTwpe3U80XJCI/eQzwzCILepAYg/b8S6U9HSZULJ9Tjd
QmJcAy87msjKF4innozarIEIsX+lQdKI6SoNaYlZbv9K4bjCxH1JVBjITqN7pupdzLUYo0uR1ojT
xd60r9Te8q6DZDw/7F8O49vfF6fAxfccIdWsq4pGreDOB1dehnkM3vaFELIw+afZOIP9iRnmzcTb
VH0NpHevQd7vA7kkukpCg5tN6ZIEDVr1BxGTns/9o3//YoNNGhFMBdhJ4uPMj5U+BIEHQoHvNyDg
V4tKbbfIjvvEBecQ0IPTigoveHqLOfPaad7Iu3UB4OSUD52yQgo0CfzMEkGAAwjCQWQRssOuG22+
e7m2Ks8LramwPdasKH4CI98OMAOI3VzFKtUMjyVJyEv1GoTK/ITi5rzodLtx8YTzcsbjuAI/PlL7
2BBcxGNgz3+OacnALXa8YZ+tTEsyK+NhRNmkp1pNSa3flU6IFNHZ3LSXdewufuW3y9CGNZOREso3
qzamufttI3R+7+tqzYgaCsZJ5WQf+CAEYgG4/5E2yfxRyYhfhPeabiIc/RYol/UNRSFfsmxNbJku
j8F3WbxXUJ7AyRQgmKMtnccb5swdTvwN5DLZPhI1J/vLCZCidDblQjEe6qgnXwf2zEqsHLlLIcua
UQgoPuqw8M0TvtWyGIZ0Ef0WrH7fUwcBgvS7C4yMM3DD28mHjcAdsgZOqAiZAsn1b/BZ2FLVR6ur
oPK3DUOZettuhNU8A6SnjZiFYC66eUZLvqJ4B6l+qCYjjIeIX5pfxpIQDnzSDNUD2zvqHom4x584
R8HtHQgMlOgdDCnUAvZr7V3JKWbDUxt8mhdzan7YTpHptRZ11CbDescPn5rvn5rfHZFG9TSIuTzt
sI18X21z8mzP7tqiMCluxXzs5xmTExCQ7a+ac0NvH9gd/a/qlGrdY5E8KJANzlDacFmGzGkvtYGH
t5EcS4TGuiHoEVGpvafMVGYQd+36xT4QB62N/6c8dvnFcHqZ+TWIxIeMLmRMMav931YAwL8g+j9l
PshQK1YIOGoQCR1nB42EQvN2JfDXA5PxBTYNQx4HYqQU/GjvwjsZGb0FzsTR9XJzTROcOPGjsa9m
v+54xPb5oFTLSZ99QJ+heRC1xq2hrl4BoFCNoNqpV8W7cPY5Ci3WIC3T45DFQ4ytfdXRfjTI9UwZ
bTpUY1ZkEQu8nnTsE8Hv/8eyIxNaflGwsf+sWZJrDp3DHyuXcP7bjvclqaX1kNEVBr6BarEWm9Xw
GABESTEe6Rm9HbnnEo6tmPY/UWVz5m+UBhKiqTJOlcSqjaXGtSOWO9fZACb0R2+jSMUZi9dJKskP
/nj4779IYu8CtE3trIiblJgysnRCTr7PvJcIDCpKR5E0mvDS1SHMbvpOWpekM0VvPt1SGaXEg2MK
CcyA/ycoOQROLTDa7uwGPh3rRzg/hxWpQ1IBVdi0ONBHl6e1l4+jWGPUJqpNpjkhWW/oxAWNQj36
QNVazxs1fEjvcYmux4fc47qWaY6b+tWaQOJ2poxrvJx99QoxvB4WXXYExxn/p/s1cSp7FkffRVzf
8eplKMQ1eQCXSPArhoCWarrp8t2qSFJlBght10gvNUM8qXosazfMB9qosTne1RJEiDuGe2Y4imuY
KdTlvyADe70mWshJfqh55ufqrdmDfBVYYL3WkPpz7+wc44IhW1T+vNHZL+/qPwxjxaMCJ4XGNc+a
xUf4vAZPwPvZVm5tiyEfUs2pIkD0vDZxuWEre2cmOyY5KjsyX5NWZsQZpyrA0MydKbOkTVXR16F7
R+chnizR5z5S5ERVHnF7FVZkTPdwEcKFMnP+LG0RsXmiAFS8Jnpy4tpo2/cOnaiVHJSBausToRky
osxTJhjxA648x+dY2ImaQqKWdyhK1+QhSH2GgBjmKbUdQaWbYEJK8DwqrimzuH9Z6G0IcV+FYzvt
IjYufgRNnpUtUOalQ2tXb3tKVdaYOrprDtq5i5uPm4X0I4T6gtB76kixnsdNbMIjVIvNriQoaX1U
PTNFYI718KEwbEM8XgHZR/sp+U4qW2w+gNMpMywR2xIdFpYKtBpNpKdHEXtyiLbYnJSNXg46mgv4
4QIFBMMVrsI27oF1qXS/kJ0nPD5fqdXm5HaBrCd3FSs5MG5XVz8MH83U/M9tzWke7WN0GS7NhFwR
eQWQr2MUZW/AMyZgSJLZdJ8gfbHy5t+FwTvGhagu27KyUu8+LOtw0u+E4EY/hLeV0eMZeaXABN7m
wmBYYse6QPJiYID+E0/PYo+PVCKRQZJ7yrkaM1KmBq3Fh/BMfZDbMa/v4v0lzUnDZc1AsshQ/+hW
CrDcyZMoQnQxVH+in6KTRZ9dspJk5F4rq2vj1VX5kYXjbZTcJ+q4AV+6HMq9T+B8QFcFZXxsQ3v8
NbAFG3opfyrm8YFQfeEazQZxZg6JLQjpVLqAL72a+dXMbN++WNQimZeuClz+PfFKclqmOD/scwRH
ZFVEbGaRowXBTBxgqlpVy8BUHDzT1+rYr5p9OL7s7fzm2C1Q7VVXb2nDVtFxb2AcmGCgUVx9oASl
QzSf6GSbK2cPeoF2/8F3XELnejvVDWg3xSjME7OVVttBwvA69Zr7FYSWao0jii0MI/18Mes/p6bm
fqZ1DNiJR65P7kI2mlH8ASCl856k7jAxHLK+pqVpicVrJOR/xgL6AyqoY7EW8Mb+Y2I5+73f6EHr
vYQCW4HTBFMZ01HlPiSYcWSb++lp7BtnAkPKahLl0ui+YEEkeZk0TTuTJduIxLxcIEdD0NR/wgDl
JI5MggS06QnW+hkK/JrWCz+o9QKKQXNr1Ly/oN1uc6jQl9YnGqzsf43Ke0re541euv2SSk9gKUo/
Vibp+BQ5/zjqPkECqrtAvyWT1L9YJTcvAHqbjyEjSGFe/R/f21+nJ2BKsPueJfrpK3hbGWwqF2yL
w0ve0bXVePvoybDRT1qPR1JE0VRU1JbDwGNsZyJg+DFqjc2nLfSEt6v+5Ug90nwtQP3iKvRGWeVM
Uq+TjHuMCBbbdSPVNuUKpOqAOkniDP7rQmrOA78zVg+1b/xV+QkBgra2hkwFimws0N3C8Cm4O8Zo
M2xYo/29CYzOIPUcRzXobPqRxV0gMvhf+kGeQi3QH8WlU1dJ1XI0eK8fsNC5gEhzTMkCcKCEqc6P
N6kWZURbhilWQrZTppJO4hSeXVRrMATYLhFBPsFzCz/J0aE/AJaRv77P7t42MLTMg9CO4Z7X3DZQ
1Y5Q6etav0JRpycT2MKpqqjZwwsN0h/IIVRzYrEZgTn5MKGKWDNTHhTRRYl4h4qXhoNJAQhuKL/T
c7k129pmmpCHvp8LwjF1MKj5C2+aV8cbSjmMvKOVIVs1lEg/oBj7DVxmpsaRTWjQAH1/buX6WWeU
OzCOmjPXPwdcdZ30eXvOxuz29G4rbq3+SdXd65u2aWPuDGXiaKhKi7F7uUpMrSXzv2FmtAzupt4z
1Q/TTlKnXy2CUWEXoqDpHdJAfabQbKYMH0cOVkBPVV3j2zSmCh/pfCjZBQYlGBxn7ntbtqBLFRNa
kNKuGqPn8aHUWI5ZGKeulRdthkRS9JyAAfNLp1eqtGeap6HTNYKTXjjrtboRnKA7fg4qz9BxDHAH
gKvou7gxoyMDscu/j7lhtqwqUXZKSH1rbnK9J94DG3hQQbOPnlpDYu8Uxwqra2So+dWQDhfmGPkW
5KwC5kL7bccDIz3mnz0e24LmcnX5Dmfq0Qs8fQaw89pGoLCBzgjwY2Am7Lumx7qPVxz4PzwgIQui
BILlDEzSlG7FgR+biVBfVl3JM96X7JjCsyRNoJY/Usu1LTmb6AKpTYL5OCuxlQhdVOEMl3kUVBXe
3llFFuAoFnRL9tt5L+WeSkNfiy16RP5W2pSiSrDYEkbwBvwyfzl9LzXXMrO6PuGYhlNkdu2dnRS1
fgIHlZ5eK2lvRdhaf0K+oS5lRsxYa1W4o+jBAoSuU75yetzBF/ZXh83GVIzEUg1TPLY9qAyZ8uXe
nrJzu8eBy4g6VUin/yNq29RLzgkxfX2bZehsSoK5vdqkK5NHeTwUzog8xMuJgSXQGGghwWCQGd4d
RWGHFiMmLMEfCr2ro6TUGOmt8ZGg3VkOeDe0Tl+lYkIxA6MgWu7TWYqM8DNkTkXw8x+AIbSq/mR0
lPOXaDnvf+zhD2d4n9CuGuWiGLIYaakfGAfM0k8sRvOJSA75aDnne0E7DSf+05W9ZrY6LurbuTT1
vAVSHNLsZoOT21UwHaVmIMPd+csh1/Gtpatx4mf1c1kaJohnpjVpAmKuBI5yx0JA+c/FkyQGSnOw
s8iFbbs3ehl9+GbppBvOu+Vh0kdV57CbnGJ62yDjQ6oHobZWUjOPJTMds0zBkcmL1Rd/JMqubnJL
A/AyEUXXRCtHqaeZbX9A2ykQgci5qkkJFe14qEWiT/Uj75zrP8zKvP0dR6ijx2buDwCHjLy9uBTI
nYkpokNwWnfJqaVFbniAVoprFJi+UBLxb5nU+5CWk1cVbtU76OJRlqLR8eRJTlbbuIQIgnm9kntH
+Kthh1o5V+w+PQesF3SVNvbGRv/JerZC/Lcclo9G5v1JHa88w7RE8ANc/AFoEk8EvQcwQWJCq0N5
2ppOPL6SLPq/cEQoJ2knvpjVjnlLZ6SIyUTLWA29jQzGerIOCSlkiMT+TFiGJzIyvk9+5XsIF36M
NMxkIOIBe5J/Moc1lDd3ENzg+oui078Yyns42cynsz5PNHhyEZuMAh9yxFOz5XDofUo6NPHM/nZf
1pnZoH9bDxbaUndJgtxGY0DevH4c85v2oEGNl1UAWrl99wWoi1Cef+Rd86eoz1zY/xOqWa44hOb6
BP6EBewon2ZnxqmTYiPj1/bgWCmhfFGejo2PuLed3WLRLNKiauebCf+MHwZziDgNzzOAR4aeLXH6
GWvWE/ZJiUDPPmMZUl/XqXP4nAoTwDDQMwfh4KDSsBGVl7FRXwTz5tMpcjzvm2AKeItfwZusoZkD
Vf4Q28TsJ6SU2/Gf3lU69eXT5Hyf90u2HvExNgHMm8d7SESCu6rSpHfp3NHgp8TlIzCxHGuOrSLf
Nx4G/aA8ujzyBCkd5jBfSmRpCK49UAC/58Aom+lRSBuo8BOMzQE67HUUNjoHiSnVU5y++V8pYUGY
Ao/vFexgzqfolYs5OCR0qI9wkEeddwn4uL7IwQUWBchtKz1TMgcVLzYDW3diK4ob6HDqsIbIc+7m
TdJyIxgt9puQfQtvJgHG/rh55n0UH+8ftTcmqNGdo17KvHHqYlW6TSgtP22rk9A4GtZXQrkcq75x
PKnj8tFukcAQdcuHtlywK2pFgxo9tOYi3HFVffqu/p0zrJW4APJMK1AmB82Wsa8irePnYi2AC6Qx
JZRnxfQZLTVzEFzqIW8mtETyBXyqY83SCcXbnmOnBWFuGq3NQMIh2/sIrm+STQPwo9r4YgPkJuWC
bbnxBYQgWFl4AksfAvw/vZP0MbQx+z91jfg/PGzIwQvmYC3+v3EnvpG8JLviM3HxV3rG5KF41CYg
7QlQnYiROotaZOCfayEXr/loGlFpJFW3aNIm6DZhj37twCYpIZSBg4MT7MY/bngf04wvQvqz4C5b
lTxWqqwmv9HLnpV6Sja2AAmi8IKO1wFFLVa0lv2dcQnA0tvqlFOcK3uhjAoH9LZSMV2u7YYA5F5+
1TgP9ifaKMtruIQuFZ31QcEM388ohWeiMYmTu2Y8aV1hX1CHJIKzPyw1ZyT4M0fyicouT0WJKMD+
CheMa9cisbocg6lKi5b+xJTT8JpECQPEnc1RQLSrALL1z1QW23K6x6oToZPRnCqaZdKkv14ZQGFk
TcKaLxkPnATJuVxYIAkd9pSWBSQjkeMgenz1rC+oRkMtBrkKyUEQUMm9aSEd+oxfRQDZJlQuI2Ou
eftPzDJ71ljndS3NQ9fLvwzu8zxPNpaUjNRBflFp/HBpSImJ13BvHtcpGyXBlyNCkuWap5RnghbF
dH44BxDy6FNr0slmGAUxgjQmXp1W4yEkmuMmFV9kVQ+cVHqUphOO0QDJqG+jQKSON42O5xsHIKHv
fJGYCkhQzIVLL4gK6fNVxvk3YyF4dN6nLpqxnTo+DE5xQN5buo5GeChieOrc+kz8o4Hicka+IOEC
zrP7zdBptaJxGwurMKU0RjCjXT3MSR80fMi/X3X5MpkeetX7oQlr8RvoREHENZwxFXddxBQAsURF
tGhaNxEEPO0WTYYVBxgVtFAJwfrBdxZc/jcpsP7jznjtOCoF1F/41OhwaBNfNqkpv0L70rhHLy/K
C2ZxrJD8ZSJGY1rd88bymUZpiNzxTO2B3re0C2Y6g7u5WzU4i+3QbLCS5mPwwvyc/faUQFF66Oa2
5/3PMWXt9JN8/g0gQx+ihmKq3bhX0amcR+ej1+PFQBM5FwA0BNKVyt7CSRxuKMxgdEZHwlOZbN/I
/4f8ctBeCWYzviDVpXR+behW7XZI7tq94Cial3jHg6R8PI3TrePk1lzX/hByu1rdd+OkMTOYDXw3
RKgWmEcp/FfaWfUqxb8dQs6HTCPfFGuHHG2lEA9R1Ev5pssQq7sUfc0w1V0bk+iaWa6AsyC/hlAD
Kpu/gaRgnTW9e0G2Pd4n4aV1BG8Zzd76704LFF2f7BCJNfgbYGOPMK1+FffDpWovUC8MPENJwCLs
F11rtXb2QaEIwxLxrobepm8XyhhL851wEOrKTExAOI9N6fcXMPoQDX8oBEtg2lXqJvY1DmbkZR9g
YriZPM9cmdZe2JaVdnwJ89j7GL1LIIZfPceYVzvJKyAY+qy6rZAmD2pC+yHUfTk89Iko1rpcUW76
AtPwSUbsqnrLzQhCMh8u08t3gAeCnJSs+ZW3Qr1ehQOTs7LT9U3LWeCI3YPG0kf9ONuUQNFMnuqT
OML8cO/BPyhGWelgLRKwSfZxvxqyZaP9f84W0Qd/4i1Df9qSJP2+jCLn8CUBr9UnP5teE3k0AgVY
tVp9O4bCR6vw4Jh9UlksJZfT0VzDHcf4GeYdWo4sOBG9InChQ6laYVoyUL/wCg62Jxwqy6e3im/g
qztZb1ggpwaxrh70jcsCRtyRcVFZCiYcbarIVrCRF/m09nmqz9vqLcZKLwMpavJ3ep0EV64tJH/C
l+83y5RKKtfCqHDIIfOYvokr+Enfg+V4G9iwIgqFRCrg/+xyq2vq2cdRs1QTgWID1zgvk//K1wCf
9eFQIzvzmSq6Hj81kZ5kJNa9a1HXtw+4HGCcc4Oy+gZGVfbCPHNWYvswNg3+boG78zYDshvAfZJT
m9it/rmTrM7NggYimCbiyHKo7R5wHJLipl39ocNFA0V052VS1xjcgE+lXZX68kjtKeIPqvjWWCgq
wtrHjmH6IyJlJf5+Z2wy9c7Hc7udanFyf9lBhwsWuCD5+aunOUw9I3ZF546uTrk+z5obUISEcJir
/Te4vGNXLtqIvywRUWQux99m72MYJnrCVcmzxxkhCRyup4U+uM1HmCsD9KjCxBVsZok0CPo2AnYh
S4Kc1avy90aHiXLdy8nHj2+gftaMI4210k332SU10oKBnD6wbzUJO8cDQKMseamoEtKeaya+IA6+
qaW9k+PNnbGk16P4GvBBwsfNVb0HJBpZ2zuwwQe+FRcFJPX98aSbZYgoHugkRDW3xawBmJ1nMOLc
rfoXz3ETA3sJY4wDMjmXmcd2Ay5yunRQmBuyiVRhQPy8u9bcNmjLdNtmnZITovM2G3mYM4WIIvdX
+cnbbitqqKfR2o9eLE4mBW64Rml+x2c4ybntmFJ8jqRnd95vwHvi+wmnpZZ2YPeGPVn5mMBL3ZXS
ctGlAGZoaDBVTZn4nGhowrzJ2QPJum/Q8fZW5K7CtA8VV0AyrLNSihvWJ/h4HEtB+aEnekP6fotp
Ti985YXKn+Uf5DsMP1yLnXr993Hf/a5v433er1TsOlNfSu8ru31o/4zQz5vTvXzmAaxqVv+KbNor
Dt/+19g2emWgjmCs3UWK8pXHCRe7imxG1Lia94GplOTsYIaBlyfH+nERcc43UMLB9TKT9Rhlj3nR
S7+PReLd4PvBS7g62YV7WieTK0Ow/PZO3g43HXwnrY6Aq0NQen/1wv1PK5FgrY1Z7zZ+ZC9qnWT1
kh1Mefx+jqZUs1w7vzzmAErMqwsvyr8e3HYbw2uKc4nvourejbfbxUb5LPfWb14EHrcblFv8U58H
fGORjRBGYyv7X3Z0frjllqeWouT3PdZXw2M9kEIkHMsDkZY5AilqZ4Wh2xKD/M/Lwo1RN0K2NfMb
sx5//GMIctBNLLEiIbJhXo3fqHj+dyx4QAvUNmMizTFlq8h+fGF6RQuDfBJnZdObEmDsN6kYLEvL
LBzoY/KGcmcKIkPF9dgposGog7HRGklxuxaWEpmPSCoh9+YV1cSMSgnrM8YfUangADupvaOfg9mV
FMkaW3I+Vx2T+zaGaI39iUd9UJJey5Hxn32wSh7AYpWHrXJNXVI80CkU22ptwf7RO6SPM3+8kmTx
EGorJRLidjCUDsbiSgIECA8Cwiq/wWni1Sp2Nv5E4F4VP8PeaJbrv39qmwS8F7iM3XyM4ay7GWOj
1JL+4WmIVa9b5Ser33pXPlTmzeeWOspavF1qj/K3lRzj3x4c4lwrOxf7FS78mS6Y8rX4FLxusX3d
fOkXhPv1m0bK12OxwyRCFqf9QMzg03lnuDhgueHp9fr6K6fsiKmIKKReImH9dePvx4FZkOPzeYaX
ZaOg29oMxUsnqCrnobrOONqGRLc+uCZhgTw/9tm+vxIxmdD8jfUNxRcqVjmxmMs3m8leRi7/5mkp
rw358C+qZ3Gib7PAzGLa/XxLOIY3l9Q4INzl5qLZbY4PdSCKfjLcGKelD5zhMWjy5ZB+OLtWpE0D
t/EbFwIcFPiESG5lp3qkPXWGzfFy2UvgA5eQBtzpmxsH8NlLv5pHovuJjUwa63R3q1NSdc955P+z
MZB2CqknjYPhboDnLBBZze5MlDbVBuT7g64nFbYbigxB9P4YxOBJWD4sxoEGbSHXhflPSqTmVZ2p
NvMV2KXrOC1feVf7K+BM8BaVnBP7f+LeMTfgkqSLO44vjyraVqoK7LnLT0iga3AbfzxCgh4L5oFr
4NBYnZNeBpofjctbDukwOUQCp8ej2Y8IWOilKfcYfIEhetlTax8C8pjU4mgQb5K2iiUyguHuC61a
xAatiB0yeqlY+kSuqYVUwkFLorKP3wMeUf3qnOOR2G7S8KbqKGrTSJhGKwJ/PPm9OFBJOEHIdyqH
D9IFcB6eJs9wNFCp8m+ZSOeXJAR2z1qadZgBWNv0DwqOLdeuGj11JGFik+ccjnfsIklFt2+1D++H
dQxmMJYO2GkoQBy/lcEaAVBfSuqhLW9ItdlhoAiFwiP3kHFkNblYhh/yqdu0M/MXEypXkLnlJyH1
L9vst5CM2xPBpOnYmJuytV0VT2a1IB+lHRQ4kb4EJl2TuH4jlxlgtNAm9mKCZB+qpZyUwwKJeN3Y
tLlEDxyQS5Cg1iI9vXUpOVC5LTeXJtEMgIHwu2NRBd4ir9m1KFbNqzi1OuK4MRlaY7huBnjIyR7I
0/HF7Y8J0yt6Lavm63kwCRRwENGItcwssOK+BwyumXppthanNPzVL/BIRShyP2SbnjSndRZwjDx/
FofY74rT38T/BSEaaumwgJo3BkKN9WiztAyJ0TwtzLzEIlb83GxOybJepWNe93sfsIR33i2YUJFL
IDiUdz6kiNEtXP/YNJmC0dIAKKYPhzzOhKNpZK4t0hc8sdQspujV2OAtMSTW7kkd34KYpm9/7Fx3
VCbog0kz6XLNopjFRRZkNEf0nyww21aZrCDXJDgYR84Ejfv94eRku1AmQP3w2Sssr1vkpUvVcjy/
m8cX7GPd6KkyGbTfnxkjs80O0sJ4E6dSa8umaVjY0mhtYcMM+/MzKIaiZ8koVVIFv5larpDwe1On
sbrgiNnRbfdc2C9nuQIcikfwpveu6U20NRG5RsyHKxJ0JUOPQwQjovtuTnRr+Irsf3iN7Dykb4ey
J+63sK2EzTS0irPTz2TnNEEDe9g+ybSIF4WwyjLTMTLZCWx+D7B0p+mr282iiemel+xsk0k15LWE
Xsz96bLAXUIKP49TDSzttJ9jCmV3Z/hd6xKMfsr1xR7pd28lWX2plxVUowIw4Zyw8PakKDlCLgsA
VwHMN5C/BoofyU9UpMvvD8Q9jLcK3EPm0NFvFzKRhVGO9GxLWTgksxQ/UVVyJpaMRT8s8PCpC2M3
edGnSBzdPIFl9PrNfQaDcz3MilE6mWL5v/gY5OPXAmgxt0PPZEbCbcvTzo9ildDrIJQ9lU3+tcE9
/Bbf/12A86WVPixl1aNC4+09x9jJR3x2oJl5pKnMphPUyfhDksZkWk6x1t7RUUeBarquuzi+sbUr
+PEAek3XvZArBxfJLNViACMBq8h7vuyI+v9qJYuhLcr19xAlv1HZUGU40knNEyAzHihcqCnhxOrF
PI5aM/QgG+DPV3hedPhQtGFSR4uvBCCUPzTHeQtUb6d/k9Gnk08rKeqYHyI9Y4UYLHh4c/oUuptH
x+tqWGrQR8A7iVwV9OHDy0oPNijG2E4DkK2dVqkgQnqvfiI5JL6RUJFBWdDMh/dCuFW6Iy56XwAj
OcE8bO3pgVZWfM2JTqZcQiA0GrMGZNi3M4LqjpoSm5pDN0UKI5kjnEhdd4zlxK6TIDyenp0GHa3P
pjKqemJjSrHvBMZDx9CzLLS38bW5eytb5aEchQWjHdTK7rF5P1lgZTAJRRpEBw1irkrnBOW+scEg
eaAWfYS6FyKBjyuA3x2bULbG2lMsOHVhz82qbL8DhE43uGIfnaSAF2w4aCrlvqogDzsnKeJyYZol
1+ge/g9UPpcv6ZxVxqx2UV6DKW5vEhWAhT3UUKztcOHqU6ATQZQjstjxktsaBKNFdi1HXjuZSK7u
rKmQnayDmBJFWjXZqBPm43m0ltSalde2wihJwvxqJPoTgqnc5jeQUtSYU3jqt+hJMd/9U9P6HR2p
RyukegQHG4+OXaXSdL7EP+GNfu+5ZYctNEe5RsvE/wsmTnPOuQ1jhzbW0XuwkxZIC1PWGOcsr1kM
K2icLTJVMjLIEwQ7w1YoqwnSrIRy8x54MI03tcw5MCsAxikzto1QhuFCi9T3va54U0+BXUhdJE39
6lRI0lraIqk0D6L2yhYduELYwLysa+qqXMSU9TJZ6hSaYaBTgI/zSKm3Y0eEG4Wwpqwjk6FELPAg
nQMMDwmApdDglUEAGQbPGu3CkXqcSUJNGeqqoJDMFcG1SfzO7z61Ff9rPl4RTln8+11R2lepEjF2
IKwcHNwK2RfGmuagS7pq/VGmvaW/wx/jpJzq7V9db1YGfCHI4Gpby1TkOwmUYzyR/nkfrUN1BYbO
ncJ130ub0DvKpOt061DZDzaNqQBORhMeC7AJlvxYQancxklwotJ9UCA3oCVT6hkqEFKpCqAurpA9
MCgVjzjSQbmo0tUTxnZkq///DQGke7CBf2qxFTgZ5Jp0/F1r6Riuc1Wk7bF/Wgg04TKevYWkgzOC
I2ByEQyRwwcObaR0DOTuNN3P2e1Xu+dMrKMm6myfGjgWqMo2aKqHqYGBr4lmT2dZ0SLYpZ+Yhqe/
Zg6Lz04/wCdiuIC2p9mVoU5zp8CTT7hogQ/lp6klJNV2UwBVQ3rz6xwHjlaXZ7t8828e8+xOlbzA
Hr0C2St3vuTb9aWlyu4bgFS/Pu0w46bpibxQeV/TDjxjAOXRqh4xMqe4T79FKo/Kyw0INeA9V8D3
IIHVHZd15m5MyllSvIMBm+jVxtVCFPjS7GD12YGSit8WYzW92PqZumJod+lpdJZvq5BIcvjG/uPw
n8suWbid7K2Yw9/uhx1OuIg5o00CKS5JjMgJt4zoSmqQzIjpEbFin8Gy/pAwZRIK99BT3a/VZ+2J
udmZs/JrsnwQMzlp9vj75TBbpQ6o5v5wIcQai1EzqKCTCFW9ATgBP7u+b+qx9dn2QP782zDuzedW
d22Z1UG8UeD4n2HBKH0HJ76BKRRFRet9JEKbjZZRGL+5BZSRRUgKCm0vfuV+Vp+64mXRaK1REEve
2PSJT5cHjc05LTbKqFkK4g9lc+2x5JVLM8QFLswQDA01g9auw81LLGcXDnWQ3b3CdgMdHd02ddwn
fIH5LkXVur9E0A5mcDg6htGEyl3K0bIS6iVd7nst92StQkBPojGaUqKPibHQk13kQwCdq0u+bZk6
pwQMKl3RGKquAeqs9C3hfGj4CwoSsi8Pz017BJYDd+fSLSh6xV0DWpA886+NepRsy1B94KTxukFh
FIVrF4IkcnCjZacRh+3SzRVBgJFHq5h/gVXOUBby+UmnMxXserOxRoLNdRQduSaWKTpNyu/8wgyq
eIg4CVzLDUDJLbbfleTK3UKSARX8w3qqAApBuDRcQj9oZ9SJj6igS1I5etqd49UDuAKJ9OsOa+Z4
0Vxc/PW+XEyvdlpcKE/be7ihXE8VLdAr28YJm6unRtChikuR/RrF92mFoNBqnii7CM5cH+lBCYdN
7z1sHkp4xQEF7fAwnw3Eh+2wW5LtYffTLjo9SaCRxQgt7SzNYIHK362ICbB7EW5wh8VRQfj2Jwlh
s73iQiCxaVfAMkwo9UQHAy9BusYABkCC38+qwyS8QjuTNacOtLhzc/GPpFq3DDtow6hxVIhLrOsP
42oJB0H9mMPzq/ZMW1gQ2KfTZkUwECaBXYUMyN7aJdyxtoGXMCUmRhcDnKMo1DyO7BRgoTcKtTo5
sYeQacq8Lm+gMLTbxG0hkp7CbSql/ucNhKHEnHUoymJN3Jhz0pUtGk2QMnaxoxiB+YEDQaKq9itt
Hv8tj8t/Iy1o1S7aVFxzq8zUTr8SqOQQ+4oSrLRFUtyNTCB9bxAjACE+vvNd1tPtK8xqe8PXq9dw
3I/4mngxBiQ30KmqdHJle1hZXY/OYojjBlAdQh6uhSYi5TSSutAdifSpdpnaBBRc3wp6gByzD6Dn
9bMUu7eN9aiIgwhEm73RwpGF4XmXj4QkUKvD5v1b7Ru44hBBS2PmPSbTXytgVgxaJEFkFnN3jSvC
0K9qDR48Qw4YZYMv8lrKued90yBuRh3egmdM0+Rvo56I2Sh53bRsdjjTPideoh1gJVmn2i01/FRA
+YydzLy/snbNiEgMI4d15UYGRNrntaQyS6INnq75by3mezRZOJkEBpykMLTTmZVo0CiV+k1stK/b
UF0Q14ZctQtYJhwpOrdjl9j5ln5RC1RTT8RA6vO2SEWHm7gJeHHyBvvoZDgh4Jr3x7dyi5urgLaO
ZwTxCxLfKYsKjQHnWQUasHu55MjDpfmCnxHStNVHBOmEA2Xl4075iZEXUANI+dYZWJNV6DUAW4Fy
rYBltyQWO1+Br45qAA/+AhOpEDqt/vnoUnewZmdy93jnM3CWSkRI6EfZ2+3JbuQn0e5hqFSwrszv
26MLkjfq/TNOMWXvz71ppG6Rqi99dyPRvflK6JERJDCaW8ZjViwUACQFwmRR/va/chWoTamXqKRc
iIrRvO+7WPuYe/VEyZBOk8ePEpNz1srZrPP4ZLfvv2Ly4Ti5aLRNR4A5HxiP+1Et1hHyqffCaqad
lrR7jtI8MYRicud3VxIetNva3yKQ1dRxuYDWNqvgo7oLdOro4/dThiOMg+c8xrcOk4awCsKJwtET
LoE5Y7SjWTUWmScIIbIY/MA+k7uhIJeLoW8L22MNTTd8fCWlkDNb3ktpbZGzKgMGOiu1BXM2p0jz
r6lShK/ttAFuFpic4B7txSU7Ht4rAaPaiD/BafDCc4DvjPFgbcEs/+BkA+zl56TXRFQuYpWvJuue
Qt+SPGLYPi4RWq+xg4swbOn+2lesdSG0e6kX7fqzVNa3eLOr9Bw9QRO6zGAMYth8hHMohhx8VbsO
zLmyl58GP45QaglRTe9RZ7HLNRYWy8gzWd4ByDxPmyP6WypxWgPce/fvjAArLZZ/EqG7LGKv/Bht
wZEZsUW7kvLXO6ytYkExSco/BOqaD0adOVXGqdOFYH7g3aceS63wbKhPAH4De+9t1bXXSHzOACwu
FSVTcTzfFX8NwkZMuqrqDh2P7NKqaUK7rzoda0P2X1vf0n6TYtB3D1bSL9kTlnWkhGn1LuuC9A3V
1iHSVbEh7HlS3LRKQ9eyOnuH/kJxyVvFzIGEmB1TMVgsetA9t1tBUNjtzz9aX4JeYpzouhdzRw5D
WmqW07UDL2NhjzRj1OK8UXlE4HxY10cqczxg1dVGrEVk6QlX0cQbt+cmVpiwDQ4DugmLSeDKCp/X
9KRCEC/jd69yqcT/MEwPD3PW+FvFVXg0hpZDRIhokMGZ55CMnezyLPY/p1yphVnCYbK9oQgACSXw
oOR+vN8bFHa9OQr/WbaJndlVM5yZjfnjKSdyPpu/z/9t8DExZHpTg0zOx/pBrav1kHtUcGJYvPaT
jHaKvynJ0B7cGuoudp0h/VGw/Y0zK+UszmLbygsBaSWhZR3AYTJ9ape+pkKgZXmDvcN79tHaU4kG
I9BCXu2M/VIuCYjKRWBCLUQAyFuHRw8dpps/jtdosIr4CBuoOdxTujOGlD+D3DpS2D1HwUbl0eZx
FUEdo8B3FubEnMPdlau/nhJPqGLbs4r+/plp4PWQ+bh22pr0GSeO8L9J6Db3EwHOO5YaOzm9gEMq
49TXP6BmHemXIp5byTY9ktKZjF6pOsDZ3IRhrWfAQMJ67R/8Rbndx8ZaaRpgJTC2RiqMjYqyC3EQ
WYNHLF5MvOoGpeJ8JekQU+JzdTXz9U6YhVUDyCeiU5AQT2BrCiqay0xrbt/2lvt13BnvAQ8xtZhQ
fyrMEY0Q9c+jc4ytLTFnRaM5AG/p+jxArxbCs+uf3Z3183tlyFuNvyBnN/gMHRkk2BGF+XAa1PPX
3icv9X2FG7AVTnNIYG5+JtrZdPsBt/IkuBmEuFPy4tV93kiO42LzsgigAw9IaOiBHXFoUwBo/Dmc
9MP14TMhMy2z6hIEgA05oWb+0brmGJhufyrcnL/06TUFXehd+bbzi06IVSdHiXy26fczLSZz/pIb
TD9NqJYi2McGFIW69ApfDcCaySLGf4PxXxQDlUwIy104Gnh6bn0Po9uMBNJhKSmhPFIR2Vk/drb5
Oyudpeh6C4jxUfS30eqyiiqRdZ0Kzu4hZjp5UBfjHda8dPIIO2ccgls3ZbYMlr54syzDJuWQp7kd
dAQQSfglzU0NFSVn/SaNIYXbvmPPeJYZ+gZASgSfuF1vM4Yos4kVP+NmHgaz3CbtPtd47XEu/6jT
kaWPUA/oR8nSq9z4e6AcrVytKMQ6UeBSKE4pWAN/06/SfoDxS6lkUZcXeygU4qloBPx7wBF5LxVU
gkgfLHxvgkWHVLacVjeQVb1Nz/1gqggsKDRhgVafL40ZBsytwlzMiIYwGU67hrRrXucXbnx+lMVs
4eEaI4xk2rrlugzwCJP3XbBvvyNgrdKqFjo0W849Ri5U4qGib8mjllqBtYHSimtQcoZLqQWpFQpi
lxUvH0jtO9X83a7iLs79VQnkGmTRnfOjF7Vktg5wd/KDRuUHV0Qi+V4TgQb28tq2hRS6omVx46Dj
U96iNztsWNoazEM0AhjzA5T4zhdiQ2SyWPoepGHS088w8A+JOgYYkPJKa2l+ResvwAVN5XddPvyb
kR+879W94xcRR0d2frzUPOdx700XM/U8XvTwybrInzujIs8MjkgjWx/kw7LgZXrH2Zcl3tmNBQ4Z
imdrQ8uxCuRJ/7gb9e8H6vHypGbNF/QSmx4M3DI5HhRDXILClFYGbwW1oq9u7PE81gusW2tdWVb3
ISwWRyRh1D70csducY24+0dbhjxRh8KV+xd9OQTiwpyNBIjZVK/FZZOJuzjHlSGmlfu5poogEjNV
sG/7liJm8qivz9ZXkI4J/kN9+EBRjSbfMaFffBHjK5uvu4ukzBjKB1Nf0nm+8qnnZ/JFic0r8Tk6
nUHH1Q7FfRMBlfs3SZ+sKqWOtSrxJVTD9U8SLMYahiN8AepFaiprCN+Lq1pk1r6vgA36PtirHDyt
hu/DcV1Kc0aGAMoVh56Se9QYIA7TIg5dRXBHnjJB2XhmsDak+uP5JivXZB2y0qz+SUMmAJkn46Zh
4TK06z7KjKaeKb6I2105VXjOFZqDPUdB1sc/RrCQsx0rT3lrQJObEv+bdpsSJ4myo1uORy/Fc5Kv
JC+UkgEzY9qJYKsP6MwCsRgzsj+GlMPybCF9w2h9nKBsZeK2fXFH9UNPpsQSn08HwTqz71/NAg8A
PxIhvy2AZeeQJFWQCbEfcl5KMVrtecGCdZt7nVqBPw/Vc4JFjQEk1hwasT+bikqepAP6v+fGRmkF
NSkNJtrCl9vAgA9P9PZ8gGktQB5QHIIoVWooEc7SGcjhFhWEqHSj8rPmvRGkGQ8he3eyll2IAWxZ
hFrcupdS1ioP85VoLbKmDXSbXp09ZKhhH308k5Kjpt7VgQ9WcrUpmCUQcJntzoUJR9OGGaXfHPgV
7r4H2LI21HflDLKQjo21utuOoDoa/DFGUi7sWMJa347tUsrVj8FLjKKaWGsmHJbBnDnjMcKLL6RJ
ZFCQhwIEAHR1IL1EIHxfZdBXZTVYXXESo65BfdXtgypXg+AhbhyjFf1ZiaSmJSgbFcOKdPglRWgH
iUhHbYmjWKPD5OkicXZ9zmDJlfPtnn2l2Sqmhk3gGK6McI0dC6RJHhz5BB/j56daTe4JEoLq8u+x
8SW98lZBlGHIU3Bax5JaYZklyStV8ulQYEfFYHxl3SDRZWgi4K5/L9R51+GRj1g5Xt8cZP3Yf54B
VpBGvmwvAlM61JQ1KuiZo2CznXVCF0LEHS3D+8ICOfITiHAYtuz6KOrL8+LeMHlrMbBW5r6ARcCA
HUpk1lYYkWrpqHqswnn4OR4YdCObr0Btyy0XLJERLR9qlrJTzIzWQP6E+5g1clcuyqyVlkAw7nV+
71Q+p22DVfuX/hRRIQ0RHgnxiIseP5RGIR0Ec2U+vXwz1VQ+DrA+r+1diKvxpMeEqkqxMG7Y7ShB
/8iNYzT5EcV4Cp6luy6DBKY/4J4lNBh6SwGEoJBO2JwclfCoOxDlb25ZeMm1luQzbDwnfvL3WW1M
7zzNkAmZDtdTZz+YBh3HXRsyRTJ05OeELEnfhrtWBDO3NQoIagFXetLD16ovp5HHLg31lZmUS/Zy
nqm10yNvmZzBQDXqmGtH1sEU6GHNyLKqrIPBaae9ztkHVIZbDAkbYM0SlLl7rjcXKuKteDjqiTVx
dA5X8lMeTHiA7UHpO2E0EnaZbhH3OznIvon19OIUc722R7O+74bAJkP0Y3CbvIPJyPyUfGbSPHTM
/WDv4GV1bZgkH/cEqAcdzpqe6IKFIitdg7zeTmLGaw5x0GPfl4pflJ1a4k421uTHKigQOKs9jo43
CLhbH+SBrVvnyLX40Ea32+OB9UOeVIwfIyv6NMWPd62LtLCiGjSQu6Fo3k5ZgAqeqJ8fzJicHMfq
8IxW9ILg5hWvUec7qjeAw9duAUNWbDcdkU8Rfg5eZ1+hRcJ0ioc5zWhwhy5jKQqjP9y9kH+mDi7w
tfzSx0lI+hRfr3EM63tDYCLH8X2wJT4o/+myheMvoQ6Td32D9KDvfaTCqxdChMw01vXJ1JE8kB05
cVz06UiARYMvPhlaBJlyOG0ApTu8oF9QcOstR4B3z1AT2EwDG9BU2+SaA9PfCSPtoh5CNdJypWuW
FlKVSBleg9Z9YlmG84UU4cj2m7WFdnD78VdEr1YKaMokcnjvVT47qXJs9N21RK38HqPGsbSuDoaD
rGDNdk0fGyk38svOQTFnjixQx8LIUZUkDk9bmz/1ergYzD/wSbqO44hzUnQCB3iL3vEWHG3FKDVB
DrMtajOspp+dVbPb1ghq7y6cLh7D1hAM0yX06fnFZiaPpexNHVjdi4n3X4QapN1zmNdvNnoOMHXM
A+S8lRRcpwJyCnTYE30oJsGh2yaIoMXJK3Gl8fnUaD30kQtqGRxbC9sKYn6SUS5+e1rCTFfQF1U5
FDeQ3oVdDIllnv5mQEw0zqYXccKZUbMUJ65ebmQjXVRlVL8nbYv/ApDthaR2C628VlqsQAv7rnQc
w34FTwPpopOpeQYjV0qMQ3rOwrsAFioa44kMIIOWs1I5zJOS+UAMRKzhOeBELZfGfZle/Fd6h07b
9lerxsi5oo89n7dsfZTaUJdlVfQLAy624FZfvCWgjLQGfqBEOiEpRjZ3aS2BgI1ska03l2IjNEFR
Thx6OXrq6vnZdznsvdg3bgthz0ufLa/7akeJiN9XmJCdeHeyh2aR5kN9U6wfEMOwAH1/DqGYcQ0z
su/KyzHqNIx/FMChMs+TcRzaAoY3/kv1zz16JqJ6LlfZKjKzrCAJa8xiatzxEsGH48Q5bls2A8SB
NiDi8ToCwjOBTZ976ymdNSIYLTbDMzDK+AFM3Xz2I/hjOT2u0EIpsioL8gDrCGz8Us+TysPyAkd7
fjH0pFUou7Riwp61xXGlxk9nzO3B0BhDdJzmlgxrBmJxeC+zR+aRBO5fq6/JGdOuN444bW5BS4mq
+jCScRBX1gU/6hZu52HdXjoyW/hsMINtEnWQZWAGVRZj59CXZngF1YP3pPXAB1lI1F3PdiVKrnF1
Kf+vISs6oFQuFa/HBT5vTTxJZkLe2jkaPlXWtLMMbH5SmyhJwHsI/XSa9eAu73iJVdMo2er0Pg6r
aVZmb/BwbciAv5bpDXm4kbSFlMWqp3vfpgnSQ85J2UMChhBQLXPhLud1AW21kiV4+cE9tSdrB9z8
6J1NP/CF/0SCQD1xX0FJUYINs8LPDhOPamRR2jmteU7xGcULxiwzsBWIg2ujxG6SAJNUoP/TraKT
Yzm1/on0gfV+rSANJvN6AU8X6NdIOoLiTlKIYkFBHYqWHDqQy+rA2IfjmZJuQoA+9CsLkEoi9VXa
ernS4XU4k9tQswtoGJ6LiHKiQifjOM6dMRCPD17IUplFC2FM12IiZU9a4uXyPF5Moi3f/Xr0X/LT
4qlikWCD9ktVmNilcRT+IYBNVRW0gTPchkRoF78RifDWaa52oj7TDZ8nB5kPlSCaOw8plOBeFNGb
W2mc90Py+CaZDetZ6yxpdADToOZEPX/ES7UmJ51SRK7UZvgUVuHEzXFN7uLoEbJbtGsr4eOvMapt
9Eg1WuEb/MZ/VWRvfFx+x2BpV4TAiMsimZlvAImzHQSgQ/j7yGRqWC6/cJnsWUCeeJJ/lQqqaeL1
33vS7LduMUhBFJ5oNkSdbsTPDjrCCXo6mXoX8g1QGRXJQCfNvS/8B+btoCg7vrAMJKe8ASOsEkxs
wrHBFMqyYmCYUbIeNkaWLbD46c46n63/PS7T75TDuBwf8Q5Btb8n54uQbtc2y3A0WUjKDAoaOja0
+B6/4S7vFx5T4jpm8yh6hJHaYW1/aXOr4PdKUlPtTeOKPvXVprwPrGcuLapTXq/SPq45lqxvsEKM
7v6pc6WeMXZ3GnotvqMr+WnN4t453Lr16ewvk3vbdsy2agqc/paaNVVZIhsUwkAZZTmd2VQyKpDQ
PwvfcgQr72qPE4ORuve2YheZcJJj7fboVnAlQOABSDU8u8w5esdUk8ikz6Z1707vF52okoScaXUM
CsHv3+ev58zGVR9ue4eMigDovAAeV7JWypcj54TUjPF4t9NynP2YH3Ll8kd9mjGfLDE2cchPdRiV
e2lz+7etkGcC8tAeX4kO2lc11dP5pgHiS99WFkmKG4BsQyEXvvUo0Zg/msSemyGO+LN4Hy1qxx3O
R+Czt22eFfAn/44t1eora8UChKbcOkqrPrpQKA308/CWTwxp0ssFFrLvfnCxOPo2I/b8FE6XZRDL
ND41giVy/43WElItPUv1hJM1Rj/xQrElXFWyIn+OaNAZMmhnc1LHkNTXZkAE4oWxsTzNS8FZvP8v
gkpWRZQXmFG7P9UCYt2QAaD932t/TGVnJIg4ScYBT3QFjvYIH02nbwIhs4YrdvSSU435G6jtOZfq
rwBOijdCt5IiqH/EiBW/ZayEzWGPujmPKlDr5BSkzMXuGxC0I/RkyRSlco3v+6Vu9nLkLxqheXrZ
xSYxnsOp4seReDxKkINwvBsOE2snKOSrs+yya3ZCACktbbwzUYPNG+kbaXLAhvE3xHW0yyrzWoZY
MQkUWdiBzIIGHC8uorwKr2RXisasDyRnIrBe80bwR4jog1VVnEKdX9UW8JC805K8w5TBMeGsGJiK
D6djhRn5Xp5NF+BYxP/rqeJmwCkQk0DonjBuPisszjTBN6JuD2fNkC8cxLOsOUScMKjXIY/dcWPX
r9zS9KvT2vtqdzyCagg6+FXK7nmd7A3eqUO9vaJcXBdl0Ee3hjQMPnIYanWs+fJUpjTX0nGYQ5sv
Ez43fLO+NS97lQVyimGlBsNs3VHzvwitpKc2T/FRgBuXxIFNr9lEdtVXm/7QGPlA0UeMaKKp2FSV
Wmpi4IsfgMC7Vm2HkWasV/djGPiL7cDAOCpXyXBzJbw7lpm1SuWXmePS+Q/WsErUJgrxwEt0c8E2
JfEh+8yig5QITyEnHswcMYzN7dld8OJlu4tN7RL2JxDKsqzzayjdhDxtpKsRXl8iUxqn4aJ28BXb
byJRF8KwYIkbBQmRgRvrt+5Y704X3bCWGc3O2pGGoGQBEUnh91HMSUPKotkSZFxKNNMxXpyjW6Cn
hR6XUGzFYzRh+y7BQu6cDtOuuut1YaH45I5sdHduYComUhGw2JJGZHQryj2JHHZSPKcd9iKFJkfG
c2+x6b4VFVpPKwJyiRwU7NgPd4thp3Yw5dEspiHpYM7P4FmPh+qbjCtv+EH2Eo17MOLwadvU874h
vQYP1+7YyEclwpQsP+hR04GPVv6O9YiXd1R/tI7ujfCNuXQhl7Uaf1xH8rEW14lAMpuhZftEKRPB
b/MEHshbjZQA0mRw+W/n2SXsXxDoBT13BEju/QZlNE6SCXpT5KZUr+KzHRIMTtKD3pEmPbipal7w
al6aZoi8zdc8fahvcbUkQUxOrOoo8y8/0L/mdVczRW724/1Pkj6fRHWoLfhA6TSRuJ1jCK+QAfKK
R9SWUrrKNRIsrSDK0Umu1Jij24iGTuTS3sSdr+njmiVkLqtfOudkG7QACpvpV/0tTd8J3Wt4e2W5
I2+aASljhfofc4UZ/OGbbaNZYZuyQ+mHy6xYzLNeDqsaTR3thZiqWwoyA7Zjr7CSMCGMrKKwNYB9
z2aNTBYDaUEa9TnnktK5uAgvTQEoUJuraLq/lTzNlAL5K4kSpR4bm3LE0m4TyXTU41M1D20CwyNN
8mdLum+1Lzj9NZ7/DdCJjT0NcK0HpofxcD5EewKndeFbN6fAcp2Jwz3Z8iMRF3abXIaUHXPM687S
XxpfxvPwLCBHafJXSx1Ck3t5joZ9pQXhDREISqpgryI3XXnsQlXZsQH0YXN7/dvb5Tkeb7xww0lZ
FxqWCSB/NT5HPHXPRXdY8hyDMpl/IEzCYb0IARVcK6LKij7llm8dI6qIDxjxIGn8gHd0DpEInw/g
HYOJTE7nOwubd5OGMWCFMmm1uy+lTcIqSfXbjn8HduLwAQDAHL2iLjFlTAkYdJ7v2PGh19YtNAfu
Wq7QWgY7xBNqCvKFzF2C3QRByOO8v91pOoozA8NS5+8LKAusiPop5cbVJeQp5b9JP3Ai5rK1aHl/
E1NPKBaLeFpqWobNsZYMfGA4vczxT0q+ttulJbz0LYQdGTaj6nDya41QLR9ujVgylBay91tuZNFa
MRctWJ4ydLmlV0nzNgXDqc7VB4EOKzWAb5qvfTqRU5GZPBfRLB/WCbd6N/mJtYUIOLlD9cqotLQb
sWX/2ygPgkNXxdEA7yYkTuEPwvS5Le878Vdb3lpQpvOujx5r4eB7i0tEXXimUhUr08SxeJNZxNTm
P57EiDZHurfhOeeqlA7PFdxdwP4FKC5f/FTTuvKj6+np5M14Wnb+nbeEa/VmUDUmoCX2DtJzWrE8
adTPukD4bs+5vBwGZVMOXJeqQ6G01AxmMHVWzq6r6CSuH9bpz1+wYvbbS7oHuV1Ev9WBJcKI6n+E
Ewz1umkn6VPdaHMRvl5xLFmfOVibIcmAkXYqF0UW89aZX9gjE/FwXVgYMw+ysLd11hZDpKw2/6NS
YR5hdOFmg3SfoGF/oF8eUGLuu0EORzc3QEJNs/1yIeh6XEmR3F5hlF63oHEVHui2FRL0yZs+UJ69
ouFmK53KuPtx1XeatOp7wMbOPDiAoxNoo79rUPlHCjrLxshrKY0HwnYv1buhEkq6o55vGeRCX5zV
GNgVmeV//HZv/RbEyg+N5XyXtExz0zWm/7Un2BNhVc4vmSsvJQSongmBA5Uq/NZsGnFchkQxxR+0
3XCu3kSEwjLDc/c9bxEAGdFCGL2A98xSXPcoH1NYSMD6Ebo8iSuyTfP1buDI4a1asGadJPTk4tHf
10w1Gg1B9NKqBl+ubwGdEeyvupu0UXLZxM09IYhXcGDym2vXrTgOeGg9hmZvjGygclUuPrDsLrZO
thb+AsL8cL54p61AbjWENbDJzKGq98Macehu2OxPbTW532QDDyC4uKAoCZaAnj76RkaLuEBmDuYa
0eccpfFcJJMYPNDZNwyddIqVSh549DoA+RkSNEblBpktQ1Jf5wYPRIIaaGR37u1EccionNXGilU7
wXtO8FyKKkPzq21WAJ463DQnj1G6fvVO6B6CvYF2JtzjmqsdAX0WWU8gEULybhGh9y64fIkRNexx
eOS1O5yf4CW5QhFMyIEYOlg9Dkgn+154RFq9xbEwfdLKtVvdVQc+ZV7zzOD1WGzCNwQEbq/NCIzp
bJNS9BVO+PtjaA0ZY0Dz6tUxuOAuLDQXhPunTUlkOb1eSRXncRPrqYa/IjtCEyIYOITuld9h5G83
0ZB0geDUY8J0K6R+7M+8T7uhrcYst3q/Y2jwOq6/okpRf84rFgzCWOu5FH5BVF42kIIpebU7bFAO
haqtwW4hL5KG0RXeHWaESfS+5tbr8Eihj6X2kzzucfPPMPCnjngjqLdOfwWd1oUBDxu9qe4/t5A+
S/CdhXqhnzTz3gi0DolzRvWAHntW2lbS/o1MjzS8FLk6EdJdc3hXeHDkYVYVG5l/vl2U0twfDLKw
o1MF24BWUtC0F40jdN+N7iDSwIp/c7CkSpgCHrtac4UVfVcr7UuuhQVs/quGxyPP5odVZTEkgB4n
LUYPQxOYfP2SVo9V54BHJo+H2bzGBsLu+TSTxGxpQL62E7ODUiCT4UmXaUrU8Tm+m8KYDvWRL3lv
TlIQAzYUZAOZE8aGVOU27fG4d+d/QIelBOSEa+ivWySKGhlLK5zlU5ZBYlOIwgZJFjT329paMyYL
x1e8+FsXX56jM5RdsEnP8lQp1lY49HHI+Gku2qbPUR3Wkn1AarpzWK3aA1lq6shjzrDvkijM/lbs
bhAiMo1/9bOtgWraU49splpYDXGfpUMxjWKcVBQzARfbMQ8K+aI9CVdtWtk9tiMgDsdlZMpvkciu
4PD0KZMdX7lq3l8b0aNaM5lbKtrFbx1mi/G0Ntc61aIiQcodVhb3010jFEAgf6idNMGRlp/iJdzI
ya/CV/2Abkyd4IZWDZfeg5qRnCFnU8afUAsmD2bG1feyrU4EPrVUAQSSTH0FSCcSXyhbFDVBZcc/
YnoLdsz1JHnOjedYg/mETBvVn+zbZ0jACQ9xAmJjQ2MVuhkLhCE1M+odW0GySh1dlZscaZdPZhU8
Kd1fvnDGQRNmFwLlYkrYn/WXak/ndVaX5ZWzaJp9/jd0EyEwD1mwsWZxBc3HwBTjdBhUfPopbjfs
mXcIlxvyZg7dsUNr2FMX0z3wjXAEEt76RBUJ/fTM/agxHVZf9nZvRgqDmk46ahOxleSzGx5EGZIN
i2iaIrGpQJtfp2LUj3vfxEtMg9s/m5Mdz+snPDYjGUbKTw1UdtvC3wLRKgyXdISVpzwk76w6nzci
VfHcFI5qInAa+gHKFqzJnmGzkUcNhnXLNS0O0tk2HN0YoR1exEiTpl7eJviGSVcEEv95Tb7hMBQI
jBwEa1Uxt4zKAwbpfoaym5AFT0bEc6/Y45/3WRIPK9RW8Jj3cFTt0rhXfyIItVwDZt1lg+SYO2OD
wv8qKuaFjqY4iM3WYejgJaFbVy1vYWS1KY0Di7Pb2jKvOpeI5tXdV9C9x3BfmIe8mzQvlhWxZfHH
Afb5YosmhbWGTGW6Vw7/RY9BEWDlIB1Z1tBOexLvUmO1LEVuX5/O8wFgFWWgqa9e0ObgPoZ6n5/o
HRQgGIEAcWETQLCAgdItbenBtwRsGcSNXNYJg8aDxinQWvbp79SwzVQwFkTiuNvejhtCRkZ29yYU
YKc+eNx8Rl7Njg+YVNtJ3ZsDYscw4OYQrz/8QArFzx4Eifj4gDJ+0z9swWxdOoZiZc4sYBfPj7wa
TP53pqmfjDQjQCdxQwHHk6S+Pl3IGi6JURyVRZ7Yef2lrapkKUyTOp0IogETlmmuWVpD9guIMWsM
KsLNCyUHQ7BzMB+m/MVSPJSTXNbJpdefCXhEOyrxA7sCIERHVlKG3ySRGWd6bD7tQRnAcmombrcf
fMWVS7kuAoHP2g6OLOGYXygAV6gjU0Iz/V+jl+kK8W8F0eUy7ZZXugLWYRt34ToY4DAUUuGr4HRE
215BU/0EnNV32qpFuwTR76tXFZ7WsfVeoxhEq8Wab5GGNIDhixo5JeUTlcpfunVDk6Yw2MsnzV7C
RTwDeKVfzdEBbMkeKVVZKaQgDYROFuqydQKSIj0XlODgPy4qKTihYyNt13tP0iZiW//ElaLAdQ6P
SS2aETI3i8JTKyg7sJJyUJ6S0JPK0SAXf4DHXN2DV2Ouf8sBJD6Yem0lmr06Z3YJ7dSxDGSsH02r
+/lqivbLXeH4l6BYFPGR60izw9TopQyNtYaCEvjAuypQk8zTVeBV9Da7quZH/KdggARUqWVaFgnR
WrW5/lpgxP9P6rgZAkWQ42omQDg6/J8v2D7MbEEJnNVNDCPCyi99N3vhOOUvkW4h3iENQULYjXD7
VVMDyuIjqzZLXhuiktcjVnJalaFAP1AeiccrNEw2ndNUmnHB2TODA1D1UulSC3b0+2KTYGafIiM1
OL7BslMmTAvKWQkjhbZdNYjlY24yNi3NckijJEXrMu+Hek+VgSQcWq8X9xBCqMyg/U82w5bT82e8
ftue416Oood+Af6Egc0Pk2HInosBFx9St9dJhjJ0oTNwC+1bnTrz568dBiyOr0Tu0EYBl7YSBZ5J
2rOd7vjURz0fn1WYRhUVuMdydaCzcwQgXpuK+nHoJI/TG0QqBNSPZ3t2gfLMfRmn9358llI09l96
HdBIgbtPfd6VE8H6z2bvCwRxiBnUUdg08tDFKSR+vZtAsNzAERQdUH+8fh6PL9SfyObza/8pbMjK
WGFGW0ZBUE0oEh+x5YXC+i3Fpnt+SGnSXZbm0+hjDb/+W2HVLjH91pQZf5+wwnTk3p9PeKtDmnFI
HVKbJ3EkA4LtORsZLZ8OMy824eIrYsHDbi5aHUYFWz8+t9l55R/zkf1BMX7Ye/LKgQRBNRte1q2+
XMy6YZDoO4vU0fLIIvkyabg7iV/Ahar0ymGx80vRk5/DZou8NQs7bWEBMi4QVvs0GXb7g2S0C0Vr
ToNBd7+fSUBeN3asafPlodI9MSy7y4sRyhqwt+9gxkLnpvRJxVYZtQ1Dcr0OVtKtvcC19hEMWIn4
nF/sq7LOq22FSe/O5sBTEoO/36fjXC1aqVQ3rWxswJCCr+j7TK9bfUjqw4QElMe3JcaTtrIgfDnb
3zEyV8z1oN0c5D6nD/Fl8f/f7pRbhlJ/K2+YZNgd7ATz04tXIA4dnfGnAkwvvM9abLmp21teDVsL
ErIwiqNyXkviZ4F0sKm6w/W4fds81R7BT9DXs0Xbbi5LkUwu9r7HTTmJTcV0jRdFpDdskr/tG6KR
JkC5r57jgIK9/tr+c9xZpuV6GCIMCcAlEBza9TEyOUNQv06fkek+EikNBFdjoUCQpITdqw6S12HF
Rs1QOcEy4Eux/+DRAXg/APXrF+mbZy+foWo18G9VyALALfFPqf0ei+NipT4rmWJz3wvF2x6JnpHp
WcIolrnQRPnC3Dr1WF3oseT6XPU74fuNuy6Kif8kHPya0QRE5BZhuFnmKmImAIeGLsLcgOXM9OSc
7Dmw8EFv7B/J6bhhWBydM4Ra/W70KNhLDyKDgV43QZX2QYDnCQJ7IzgHP/rJDnKbeRE7WyX3oAY0
+UckKStxIxWG2zr58oI0cdf+bnOG/HVq9MFIKstk9lMAJS1tPrzvZfi6crc5fddKh+cGbisgIm0o
foBHot4jQq1lmAEyeuLqoEOk+j0O/XoEz3V/5oJ/FlnKYtmvezDT/gKpD0Y94JQhK3kclhhZLvdF
XGW9CdHsMypZtV9KUuu/Rk0k7kgxMlCnjvfINZzn2QivtgKwaUZLe0206fEVT5piBeRTmLwn+ZEa
eXu/milaZk4ZH214QkNuGr+Mlpx1QzBhZbzvvCVK9RrZ773ea5cjXbz0Li5syhEXB1ObXh6FHCUe
cyXzxKHGdTDP+8lzpRVgI/YMVT0kT0iram61WJQggpDuBkC2aK5isy0yJlyCoig/53q2+SzPe45J
D/CJExKYLgKAt234Gw61k3svOqqLcGfJ2AZGoJevak4N4zePCviXBEcYhoGBTgVIan5UeWzSmfBq
rSnAfSLyaCy1nZ/5JAaLdwaGXVbslVVe/EAcYegT6biBYJZJjXOaCVfWFEtSoCpYFRf6reC71dKJ
o8c/+YS/p3AAMGfaCHLFr8AlcVcfAed31w3mGdHF9t4F6bLxt4vqZIX800Fl+BTbduQZIcPv3fm2
gF6FYinHtjiWdaqZmVNPXo9cUij/XLl7v5Hu7JGMlPReXXs1sjGWuLtTVM8sPiYHlazfV7w2M6SE
/a1BmiKSXc0JG1ak3eJr/wuTyguzmOHIlN5egx9VFbRbBwapfnre+mCHujm4xb6kxDZb1iIgvGR4
FEr7FglwGpH+fEsxNcTC5hOsj55wVEzm43nfw0eZfQr0QGSO3PlGANEWiwGok0ZKEUTKCf7HNYmd
0iQG6BQLVCEfU4ct+TkNcNsp+YdZaVVpnPfxWFOPaD1ccr7nuqwoXgrWGPXTeVQhSdc77IXJ6Vsj
kmmFcLOxP1FmLzyrv+I2JZg3AvYXCteNAGXm1IrCds9Q4TMVz6TwKcTLmeiQeQyaax9Lwb91CmgP
R9bH91M9uLqUXRVPjpRAksOaojz5/srBuYi04/3Dn4PtKz/teYHxYoR0cTNLzaM7PgdgvQ/Tdj0d
aSQnjzfqukNYpi9I4CQHBCEBC6+HCzlWLjQPBs6Ramiyu2N8ZdidX1hRD5/eA/BWJAFsq5+jrtJB
7hL2sNvQKzcVkFU9Kn3O3Qq74Vh4s3iNHu1i+Y11xC6eWJH4VlamlX8e6ZlNh8gEeCKV2XVh5Gm1
B+e7cPdRm3Bb0iDUN04679QKhldIuxB76p0HApRpTkDxfEXyCu5BRL/uDi2M10Y76GHVWGDMG7ls
wGS8qCzir/hEupH+pWs/9Hocm4Gj6xgQyRjaMIMlhzv4jk3FToLkn/obCjH87v2DS8L91l2ac4hC
fZZI6soVQNwwppibTaXvczJ0Vhn/XWNpn292ruiUWXL90SxKvR9LpMWsMBztFocTT350SIQtMEJy
/j0qLKpsGv4BxVQn6Am2CmcgyvkCZY9dNzFWpuVOr6kBlJg9Agqdq51gRHiq28DQH2rTej93z9xE
CS8CCx+SbOgtY7ZUMhfe2PtKLY6sXuAzCHh8nSMf2iQ+ENXCQS+evUkJuZitqUfv25oi+R2lTTWT
5Hnfc8Gavj4a4a2YklLbi4APOSLx9uY/d+2ujpmkuThrfWjkuhUtTIC14qo2hKEgtJc3XhT4QLOa
TTQ91tPd+oGviMVD2/u5VHaTBiDqy8p3dirq+XrdGI1O3hJjOYqL4WcmTR1a0aLXq/S0FBpSMq9/
1awcWzfjs4k3MRjXOYllZaqKvsLmjs+bDFS/pX98OC17oWjdZ6vsp8Z0Sr+4FSCLsO6ojZ1gqoiU
GGh/JuQnCpDP8rwUj5X78thqblfGWy1r/7gYa/SWTCyjVyU86ZEsOHrrnkJo45idazSqvKGIXl1D
dG8sicWY1vrqSot0YqnnQ6sBGShzOWFeLgFvdoKFUbmr1PVVNp+ywwJREfnx7Z9UFNVA3Cu3Wadd
WMZaFFspfVKENM9cFAXgLq5/iEydnS31CHb33I77VULsvFXefnqwaGRsYSNS/9xEdQ0QaYBEaUJD
s/ArKIALdzVgnpbkLwIlS0y+9k+1b+IkXYTr2zu3Nrkrk0Hl/4323keKxo45o0Gultl+oGKpwLNu
k3uLJKZAmPsfK6O+rUXewXke12h8XrJuBnVlrvZlk19YmK0ZCUmDIHsFITV0PzlEuGDDYn8c6205
4eQYV+fe69g7YLmz1MFFhgYkCvIJB/BY3/luK41/oVQtCvGSV6nrzL/KeSXsM0vpHAsOnCy5Izr8
2tMrk4/20kNYwQQm0D2Qkf/nx4neOO7bjKvWE1lAP55O+QZEDEoat7QYjTyGCBd8IvwQ6kRbsILl
RrgopGEQJrvN3QNGCZtsTgAujRY7DVANRGBDJd16GqmV2s5bCoQj+jJCXETZZ7ylz5NO9CvoJI/b
yumQtnsKpZBDNsGYUQ652DTJVemRt87woa8fxnu/M0C3a5ON15l7Wb2JOlcsq9BceUDgbOzxvhuj
PW7IGNRIncepynRU7xRIdUlK7+45Eq4eymNrswO71VOV4lVOkvtHI0OpSM6qX7njq5WF9Wd2CO8/
SP5/xxNDxOzz8UXB94bOxGjTO5Er1YDX+drifh5trHqzBqtXFUHD5eMoY6HegogB34H0+mbmV383
cg+yogX6/rSiaKvmBkr6j/VgQWjX6wgbKFQW/uApGKxsFBrEI8729qykaPQE5HudARgPdRhU7rx0
o6do7OrJML2j/GPJKkEA94rnPIU8/QMKosDr7Bqin6u5vu4vxXD7Qo8851PBdS1aShFSkQXE3oEt
16zFzEtNX5/PiKgysykPvIuvxka2QruzpWWXx7B2gqSc3c/+r7zMdPYXfQc7LH4sPqns/geUI5AO
afoVagfAVRcUO91XeGXs5mTxbegtRegotSET901yi8V0xO8RBMl4z0g+SLa2YvrkeAkCK3kIi6gO
kOib8dkuiszihiZ+pfcZKMiAYG/I64lc8jI+7WPtFs+7wvwNkXdwYmLeV6+iHmtAandSaKonP4Rp
wuUQQmrrTHJeWp2uN9aPsx7MD4/zC4eRH1YV/pdqfQKat4hl2G5JreR2zY9/L/C9JMKGJQmGUN//
VLS+vWkh431k8CoOJQgeZB2Qg8L0aoEZwpYRNZS9DDByR4pqo7t9xJxdXGyEwoRYdBOBbBHY6bd/
M+4r2yJPYT8C3T84aYC/nl6LD9kj0Jk4s6uzCw2T1fvvttZzqT+VgOpa1UoWL6xGyXe0ULd/gJOj
4TRacxGx1Yr14vSJ4KnjB/7HZGpGL4AMxo3XrXXvtipv7bu1qLnB9M1438KyCR+gkga3mx8UK6pi
Y3K4yDxY5vTk89w9StWNq8eYtaw8MhLWpxazmny8OulCTQ5tNYUHevJ1Ur7lgXP7AzHj/dkhz+iz
H/upyP+uzE9vvTjdvGj+dy6r0T3fiVvIHLY4xtqzMPAkPn/nTPql2hT/VG66lgm/e0vgoZFHlQgC
vjH85EoQIEapepZOcYfmKRHza4ChT8whGiqlJQL7T6oWtz3PloHuFuzfyqbet/rr0g3bT+FlDAdB
KxrVdYhrEnsomySDBX+fbGPABr37BhAgYkt7A5WbZ1SxHEs04GkWNNgLtAbyQLC1iEXfoB79tsDi
ZZYN6ttuFOMUW6b0aW4NGrFmFEo7JYR/BuV0TxrA73mMNGjCjlyCwUBwAWl948F5zl0sJoqh3PEv
Keyp0+ut2qXgu/mWXshPh7NrGWIaGPTwENINDwKa5uuJHMURauq2D+RqtQ/HJmSQoJjM/auLR1ir
4X4F7VoqiX5wOrDWwJik7d/JRkw0LXTnEIJJzYa05QTeDlxwc0VEPBvIO010ukr+lbsJgx7PGlkV
5T1gdiogo7Zpo1sYLTikK+5TBWcUk4nwYgztFBXuLQ3JU9rlDF7Jvs/x2zh7VibOPzcl2DCvkJA3
oG+g4xlgnh8DHWC7qqYyXNrGdh1/rVOhFHwUMGqsNiSbhjdPUp6j2fTEyyAUmGV3JNUIiRbhCYXL
mLuuD37u8q8cXaLaYc/KTieooQqWBBJqm0FQfbrVnKuJziywDwM+41cCLfyplo+oWOTkwGJXdpH5
OWgpQDaiKJWYXz/DNh6FubTI/EDbTdyUEZnoVDFhjAAVQGNFA4wFytEmvFdh2NBT54GYjOt0YcxX
MKv+PigB0MWa49JVnbPZ2rsUQats3GoZfk4CnnKqFMCyzXsqIl9kx/qfYs9yYJXjO9ZTuCARxpMy
AJAmvnzLu7gezmUn6Q6y/bDR8Wb/eqmy3ueEWlULARrfzYbfZOeUt2VDZ2Qh9Juy4VIHQBsG2VcM
pqao2FVtVqr683DqGW3DYkwMgCF6ZFTxylmqendP19jhjhbN/5RDRy0RBlSfiYeIVXi+aAGzismI
GPmRBXdCctHPogXUWeA0VO3zglfw1zuAr7y0jESHsb/94z8EESnOYOvs8D+IC7MMVKSvagOXoiNd
dLvavUFbKgYFetdms7JWoLRDIQE8BW+sBs70YYtUhyQKvGvI2h4+50eieW4un2db+IiiCtJs5ecX
WgJjcUANuR1bp4HKp/yyNFica/fPONXET7qNJbx2H26f65Y4LYhGSVy+c7kOtIJInSzw4wCoTolC
Yo+V7EvWsD3gN2h3cS3049OfrQ2kLQOQRN0PAyGWJsiIclPkWZkXybwmh/wV6ZC/grJCaNCrBmyz
N+NrWCTce7147aP8rdYGzrx8g25zLfhv8wcm0truemdTziZGoq2IUQ5s9MbINsaclJmVukPJWlKX
vINdL95EUE+7SrrEvzrhSu4v/UHYfNoB6mswenII+oiYNhK8+gXL62te1WNDdIRnUUpRjH0lAsFQ
ed0HWjKIQ8TX3YWG6t+KHz7zpD/JfjeQnN7cO9C24CcwxjzA7WvTPTJMv1XbnAU3Px3L6YhochLU
x8PRJrNQTzZdBa6gXSso07m532kGXnE5pIry1jOIvUIMxn49yIjOXULZBblog38R3i1BT5P5Az3E
0Hm9azSTCwLw3ZgqUl5QgdKxP3Ofu9S43GzetzJNxrHF3vxwJg05iMqBjh9vShDwA7E12vPG/7E5
uJiY/SkaupFxQH2y0ddF8r97C+rOzcPi2KyEJjkEQD1UtRyS8IjnOqwZzhaNBloNpZv4ALnYt4jV
syb+AP5cjvXgrPK19U7hdu+nsKImg/cOKLWXFgnC5wVpDAjRbamQ4iMxqGkgYiV+kq9enIuqPQeB
fRFv9PAlRgxO90mprkAVj8btTGL0G7gpogjyaxhqtPms2zuM+eDllYFVwW/cGmRVA3Ob/8WkqUdc
WtHaPViG9Yl/wO5AAvAfmbro3ODQUYOv6qZgTs3y9o6KEUYzSjSpbTF/OtRv86w4FNHEeoSNLtd8
6sAEXuz4BnGLOuWfKvbbQbdgPkD0iCWQ1S4rmfMQK9dCoMJm+AXeMjof2RmB3hRK6lt3w82c8NIw
01qEzCHfAPnujy4IdWOtuEiXMWLyUrsVKGYoc6wXzkbyclIVgBHu6mzbzj2UXhZ02vQaL4Rsu1MC
otL7TkELhFPYrnN80gKlIC56IS5TM3IVtPCdYxILM1QV/kq+OhW8F3uCXNn2yoiR9CpaEBnDxu7y
4qha2ZbSNaIJ1ry8ATMuJoXgdjQaYOXTA6oivivR32e3nAQrQV6+3VsrjdoId9X99BOmlT4m8Vob
lytcaB6y/xu7WTeQsbpQfjFwekhswFtL98rG8K75ajQdtZXNt//LsY2PLNU6dFn4wU8SfdczNZFU
JisB3D4tcLvmoZsLbWwr0SrDPUjv3Tiq4HLSjnvolEvByVDVmhE6dT9fqWXemAZ8nEMX1st8lYzz
L7BLKALSfkLe/YL1XcqdN3tXQ3rpolmX3kbuYriX0oH21qbrVsEgabfrKLNBtnpKkRS/gAo4/FJz
jvUTA7xUOQPD2Orw885qJtNrwnv8/6uIfidIGt6nFhIfeZs3hMza06o8Dq8rGFN2u4zjZOVbIGeX
CdeNWIbpoVzZsl5uQpwVS1SvWMtIxvQ6tNnF4T3JuKvmXzRjcaJQlN0/v4w0yCzOIN4SNU3H/viT
cN9WQ4jEo0qP+QiwIfB2sR4ZdxCaoZB3WCdA+RTCeRW5FjhUvdStA57bcQRKa3kqa+1L4PAFXbbo
O4BuM6MTpcwZPfPSV7jAt2ioPQRuSujpO6j+URDHyfahyJSw9WWTqCY9n5ZTA8033nPh4RiBds/I
BxEjsmLU9A6iw1LrkuQut/ofZ5MqQY+tByOB+zfZHOpImt85qFWV0Op3DJZPlz2oyInM7SKTZ4sJ
wwpjlb7MzBBEZN7bEk6TFhbg71/TIvvh9IE2ratzx6dw6xP/rLLD2WaWwyUcECF3EOncpOlAe9bo
y+mBVCblcGq9bcbBPqW08OrH6Rz2gMvstIbe9NmscrZOzRGStM3EpQzVnpaCzCqWCR8Sz+18p1gt
RrdpAcrN2orpgCp9xieukde5kd/YHB5HyFeku1Pfg+YZKhPQGghx81lu1L6SUIQ7s4YxbOt4AiRv
Aq8+E2qsSlvd2d6IBLKKjlFK/tQQvK5rBtITeff9eEADO/nAUCY5XcQnIhAQf+pO20LYfWUL/eCh
a49wrWjzgeOGhXQ/Gt4Amu0X73eCznz1P1FnVjBk+8RpMONq56XE8Eg2PHlJ/WUMWYDVtNUOpg0g
sXsdtjue2AqjOuglBeYH9RaY+KTsTUSlySlXJAgztl/Ezu1Dv62Kuq7d3acDQ45nE9ZBanyVVQKr
9zdaGyyo8G4wL277VMbQcFLMIl07aX3Gsc9Ph+gU/wYaYjW3XE/2E4ylNQvP9EDRob2CtSUYchkg
G21/08LitZ/J5xlcN80xiFt25jJcSoCHH9BVuuBfgiTg0hIcxp7mnV5QFEWKvuO2ADErizTIa1sK
Picwo//cL7tuephVAibuwjVbJUgqGxuGSlX3CkuqIMGDtwPn50yvcnQOYuAzs1IsVcoFZAg1ej9C
mvkaq0djzNpYPi9fA3lhRASxTrecKcn5tmBWad4KdPkLYiq7MHu1uCWbIKZxwPwZbJ3F1hWkwlhU
fxihm/r0VpJ0EVp8h6lE19BVQ47MZ4Cw3XRf01rAWmpki92T68kx7snCtl8EnOx4AN5Ec5w8yEbh
vs7l7eWckr/SZ89/utxjfDC+Jl0yYxbDCfr9JMkmX1XwlckuMyLg1rVdrYi5Ci1rjOPzQOM6xDyh
/qfgT02JhDiBlC6jq19yYfHzCk+vX+/Wqxo5piNVAAR/1NIrq7kytwOwEAZNzV8+ycUc8zmkoBKS
GatmjKG3PjRA15t50Sa4HOF/VIGoDcOLh1745Lz0vVJg9E9hwIZP99M44A5PDirh3Ho6g/FxP/vr
WG9CciG+2WqHwmasQ0GVjU87R+p3Omp6HP/r0Iwz0J54+lkr3VsCXjOdy6/gPfYmsMD/WhtkYkir
bChXoa2wtEMimOH6swY4r6e7HYmQNVe+NIEwxTL8lq7I+RlPtEHcKsQmzpD4AscLE7SpppS2RRUi
mXkflYgTsg3a8LzibZNhyRZNPivrFLfBQZbwXlESf4gdJry8gVTK+/QbOJWvVXjEGi5wg1syJ96v
JUApMQzpLZzO4O1d0wlmKKhAZbNk/+d1sRSLY4N0CWh8GYlgp6k5zzlJMTqc0vYNzfr20TOVISLI
lgkzRAt0w+3UlmOABoWvEfUC8uz0QWoxX+7IGP8vchJr89GB4QgxRYFxmcZ2z8hTzTN8jSGB4YPK
aehCx16EM/Yg9nTDbu1+ciw4jjgVcpV2XE1WxijMcIF0DspW/G0tXmisQswDccyM/v9CJlbL0C4k
HuEUHp7UZDa8UFt4sWwKF6IA7QuGkNe9CmK+YGJvx87WwSyebzYps9LWNz5ifNw6Bx6rtMu1lS5W
jx5I4CQnWhK9MICCv93XRAKsWXO+OUpfJVZsE1ALT6WKN64PC0hOXM3B8Ypp9E8/rxVRh9hSRIr4
co2w83E6SjsF3XnruZg99Q9UkUdbhLjuEkkL3hHTIgF9qIIxtiYqtbSwxaR41RmEl7HNN3cs01aY
BKjcNF16oxqHwG/OV/k5CMzVAwFtLnTkeXmQew/fiEm0nOyR7ztwOlIfyDTr+zP6kUBearKnved+
o2ErlFYpt2/KQ+jjuK0pDFWvlK7KTVEb5aTpItnt8JJp+B4+pSyWNVu+xou4ATnzwIzTsjnLIviu
kwvA3a4enVbK60ftJo0VQ4Xz4AlFtDlPSbdqqCADaXrYcKppI/P4ZS76PVWuuhZ3hUQF6IBt0/Ob
EQ/PV3a8gwPsTGQqMK9YQIeNc2JGfN3/vOuvdz65f1u/NUPQwYTKk4lkl8Q+JY4H0iFoL/q7CEeM
mk1Q10xzAlBSLTY+sy1Nno/OQhSJDwVRbs8TfQY+O86v2LGA3s2Sod18iVKXWSNCUMzQiQomIQHY
5s5jcRl1Zjmz1exIg4qGpASuzf+arcb8Jxy0t/UpcyPxkrx9G/ErIKSFe9wkMZIJKaE/t+PwDRrz
k0LhVEFSiHzh/wpn7HN0cLeJO0XsmTGtCtJEpX2JoV1cX4D5FOyYidx8a2KU0zaMVkYEg146B+s7
i6c7DbmRtSpz/Hnf2VYD3vF3iqnADKz2CtLAsENgLib2sHySZzpDo++k6jco+GVOD9BxTN2USZdd
/bZTegYvYIUHjrLw4rxoB87xOhMzVAN2k4g/ar6yOq2vMZaYzaZ6LireW6XOzwbVVcwQK6OCYTeU
W5d495XMv2av+RUYUB6SFhIhPEQF1yhyM5lCUyqd1hr44icrOqVho2nNKk+Fli5GPqFh1KIPy289
xMV03y2zh7oQx/aQWecVn9tYPWLLS3PnMcCOYUIqa0fnAVNjlXFepziiz0TaUzAjUrqQNb7VtMj+
Z4neYRKq6ae4rGB4LPz+R0i0bfwqZ5CFBscdIXMU0KVaNKJIjnCzl8P/Daa8iuePoRuXg5fi9gYP
EPbvK37uf5k90vTnllszZqV7PGuF/JO0qHnXtB9bJbtRSH8bVWy/nfY4JQt0/1XlT5q8cj1f9URJ
J1ejLMD+KG016VJNPAGMibkXXVi2hs+CnfQIA2eUXcrV1WoOQz5jTclp0xjwMfUYPNAfJ1Co/Xlx
jI9PcZxE/NQQnVfgQAxTILtR1qsQMrWixn374zuC8/KAMDlCK9vvSolp9OOWgk/VuJm7jZp2wM8n
zrjiPG4lUEKzJ5NacjDHVVs/yKOyPYncpbn1J4jEPRzW7LHaWXMFh4KJL3w61T6p/Kj0PD+uqPbY
qt+mpwMM5WXjkb5CjWulbH8k9CYl8O8JXqOxIHAtszRsKrdVFdeX3I0V6VRE8pIjKWCs2tZlgwT4
eHpa+YEC2z3S/5BDptfYqQIzG5wOm80zwXYoiV9bCIZ0LB/RGNVfnXKpMPU+nlWCV0FqcfW0tHuC
2O2D8lPOvTDQr/+HCzQprXuqOTVjSNGvbLI3u5Br2wLhNxNwkNFzYDS6SRUt8s1JWfTcKZoc5sQf
JbpGU4pi6d8tiFnRWjQQWtUjYRF8pn/0sOVYlz413I8Nnr8lnY7bfN509s1hyTyuhgD8lUHVPbga
dC9ZH84doM42DVwzmyJGPrchtz+Gs7DZ1Bso1HLbK/puQrqgjokKDm4JjnefKcWoJ0a0R7GJ6Hcg
QzPOzAUwRer+UZez6Y7pdLRHyuXvnleZ/bEqIeEYJ4iUAWsg28ZSChTEKDi0XYaLU0R7CTelTlD6
q4R69rx/tXfttN6e3Kif5WMqXPy5yX7M+Xn2kUVwXqViNuAP4QRRLwYW14yUFcvmgif9h4rv0TUZ
exLDo34Es0Ge4f2SfH1OoLwknONrmTcjCiteFdk73sxD2QiW2rDY/e1gJ2h8/3I8R7K6d84/5VYD
puCQhzKTQBWNi67KuPl6Xf5yDkPMN43Ny8lBrw//7RpYfhs2hOTQcW0Wnu3gR7zOkyLITdTIgmhM
coEonHVjdJ0rZbMiAnasozX9NeUADUwv3wJkQccJt9jFlsHB+wJcD6Sf4FyTis+hh2UX7WfU5Vat
rzOqe2JLLsRHJUgmOZJ1LftPiVphWnDbvtpqyV91NaHfs9E8Ip+4Oog7opCjtyEdOKhCseCVRAgE
I8/8pqznszK06ICo/jp3mgz2pdpU6+umGLIHAKrLoUDkjYJKEge1U8jjxVc79QkyQQi3BDkDK8jQ
K4YU9mAAeAeHfsewQfAc37KvUGU9GELsTCJy9mrCqjFIxNu023Rk6OVh+XPt+I25J6p/g5CRul6m
9FlkLumhT2hXVkOwj20Fw9HEriYKEPVvtzyRlDzAVLaPX4y/xSkuOJS83Hlz6QKp9Rf+eceIy0gK
zgWHCxl92kbu7ab0Lb4PSihcoQnitNQsJRvXpMLGZ/eiyVJnncvBfUKQouNWlPR9d5AmDbdP1m+k
3IqfrSESzZacNdw1nSMWY9I3AtGLJbm5Z8itbOwjD8ff/0PTUe6Q5YMn46klrrs4JooX+kL7dLqO
oa3zL8hs7UeE/MATf0Ejx4VA6M57PUe4sECs3r8vkT8gfEhgsnBdjQ0/UO8+BhMTh/1M4Vv2Jl/I
Gywm0h8TzdzPBgjRBrpIUNLfrdA1g3QMC09jDQPfpQx/UDb1B4shJS7eIp15kPOIz7dBNS4H/f/g
gpteW8F7aVh+3wfk+EvoQT/Wzv996JWdWdfdCfJOka050gCpgiBG0rbXywKyEyIZEkUnV8jtrvik
C1tIKYTU8sJhVDGeV4SCbpglwSW6ssX55p77x43Ynnab7m2f8WJEhGvD03w6zAD+T9kM6/PNmsBT
H/MdbWWsoAzBOb6Rlm/rhHmsNatplUNusn9PKm2f8cacdOKrYvr4OpETx3SHDlfCdvLSfUOTihSW
+b9NnXe1+ieaSNxdDYn/fzpBE6b3Vuy5fGnFnlklmEds490y8hUFz5NArCSKa3Y8wt9S6cdbAsYd
lTTjh54s2CeeRSAjUAguY1Wk7ZU2o+ryCcN9HrYPL7GC1xibRbiPa5y5JnCnV4YGvBB2fFutBFXr
qTQ6C52dKU2xavDvfAy4+TirkoZW7AcJXfS/dU4Wyx5ZiY6DPdDHAyXJ2yPJp1YHojCGuA/PA/ST
O3bCHmfvdZjv0Jn07A/8U+OpJ7ru/WM58f/MoybBoJbSq9CnU8+ma73/NHRCYnDeAEaNm11lKiXx
aHY6o1/Cz4+rYAaFGAmT3NnW1R58a8xku3Cz6zpoSZPqtutEHY/uu3DxGbbcs+6Zxw3rOauRtVr7
ZRaCMQ5NyQwx8IOwfQFtmbccgjm62aFL1nYWEEZo/lJ8LjDA6JVlg9r0RTnszc2XeGVV9M4Mwquy
ew/7TBBCHSJvD6Ln5LRDyKZ/FWtVYg04eAbfHcqaDFjsYbxxOwHuJK1cho9/eds+dTsiAJ/skiOv
l1luPm/TiooMe+/NaJwPc4reUAKAi1HqjZ946M31iCHRVMgYEDiBTeWkIegSXvUqbkMr9N3SzUcN
pE+efw5SC32ODTnMDb0iI2P3EIXjiKqgpKcm3xWugDIQldNS4Y1DbN6vEZInsTnPazJrQ+Uzj0PG
QdvU6dgd7qQAgQjWV1ug45SI+UvlfWHOpTWL/+ILs2TJM+4ck5kI98M0RhFzjkEcE4bHkGKGV3aq
QtrS9UIl9hsYGp9B2uE06F5CaCDby2FOFHYotih36fKGgVOKM9sHjn6TRKqqo+HC365Bx/2d+69g
bnFOMU7eeIkbbubhMspqT5t1xwCTtRV3UBp6JZDe1ACP/tOuGls3CARa4bNL8Hlw8P5L47BzAXsj
XTArSiEiC+VeXQpiqAObuZjHugaVns7YNxhy2SqXIkIxXBTxK8HvPC/P76ytfVZXyi74C/n28JqT
8oPt/Pk8S9T6NOASPo16tbHltjTxkCaaoM48Ufye8N1ht6tVo1zAwx9LjpY44XgFb0QObHyP9hkr
O0hLPmDkh5FMfaRC/clgCo1C+aReH6WBBTn9rAWmjRzXWNiRKQPqNPsy/TgBvEozjtVwKWZlKpql
rwP4cnNdWJHX1q5QJGgFjpJ845C7VmNTy2eWAYsa7GEjqMRFZFtmLpIVJDOi1QHD2i9iNhPOmylc
lrxOp0AdWQCzKdCEbiFBNQKUBYjTOysCoLKMnFODpa4gDmGtGmgKwOerMPY2BlACdVI5zwONfS9V
PL0cZl+ReMrKcP7WDc+2HrydSOCnGbAVkMobewq4YbxEjCPOhKVrG0JblrxA6NTwpw4jMunN/ne2
t6jgQ8U1F94ONYNXexkeHCzvx563VBmPxdUGJgDLZdTgU9vAQjubKXpQkoR8XS1bE5NEyrWF2C55
78o/uCoMIPr2MY5hh0VaJW+r7oSsp13dEiP7RJhm/V+cCpGpoGT+xIqI5ANsdt/z3967AEEaRd9x
2hmb5cLYZgcd5nEgcKuC7piZ01umWUazvnPsqdr2uNYL3YG+9caZd+F6UMjm+8GkWa0YgzjHnwiq
TusuqmADwlUxNCeqJpMkapcZ9To7hUdwq/vL14LaTdKCccfKe4LjJLjzK2Mj+FjZicndcWTBMQj1
QLTDh/sxs7J2AB/F1OWIRAEEHVFV10i3/17k6I3JatUeK6LcGCcliuD5/WXy8Vg0ZzXpOr8BHXjT
Roy77Zru+TYcq/OWhzJWVkVsmmS5PuE/rcEHr7IRU1/nQZsXvLHNz6mbdwI1FmHEaVpemEhKQrLs
dOUbEhBz9NEkEfE3pPskbAgsvPvhl3cCe/OO7EhBxDGaHDJf/3sKiawQZ670GZSKsDc0FY6ZyBkl
CXyUI04oV7mp4CduxxBB+Eh/t2NtOBUw8NldA7epCjYqBBqlziVi39LEOSvgFtBaNnLbyHvqaNU/
bIYD8TpIS8qk9Ek44DiJJ6OUt/+gnOk+s/1OLs252IbrnFaYZYvpAa1IUqrRDy2Y+Kz9aW0BBd7p
srtokG4xu73yr39YqnpDS0YBJuEdlBv35unlQOMFunz45GNHMIghLtkgNWZeYV9IwaYpBryH3IRx
0Hx51M3UHfoXJ8DpiOne28bvHVb+ui3Uh53dg++5N6KoQto2uEzrTdDibv3E10vFwmG2gdCvBqXs
gBiaUq05s17twPZgJiMm2J4whmancxwYG6rEcf2maipl8/Y8IHomiSZ0Gxugp+e5tteJilsNoLjV
6jTdsvEDrUJqFsvzV0mNilGNibzJuiaksm1ebb2D7Ifdz2s9SRHet1LzST0VHiXwLr0iCgEtvHIo
+me726TVc5+91gtwqXMb8GIa9kimJVx2pD+HBJdLGZZblWtiJpBmxB2HESWWn+e7MxqIBBshNjdk
P2pPqDBGzBW3vLYGk76b5sVOl9yma3FdkY5GQ7G9z6zSJ6Bl1gsqrmxtjECS8cYBTRbQ/v7rv9Nk
IJp/WfBher7QKZI4tyLi03M57UbSar4ntmN448wkPLU3jPHNTRD625zuAYgGWO829ubrRiejLLFL
H2weSEIrM1aA7374MkSAb7jRnHniS3t5TXqktl2gQvtDDpuMevBCoxtWFyK7m0GCfDqxfev5EVXQ
VfZ/dSs0H+f0FH07VbtJ0MzWZtfQtiX90bKjANTXz6n0ZMqeS/W7dguGrfVQ5OSpc5Uv+2AMIJgc
bvUk/13OjHnMtVoyiw9xKpn88m4NiN6/MYHOLgJ+sNni2Lx28UicPA+/puttZZ+hD+Jwoh1DDjDU
W1fWmqX4quJ5lDo6Q4U9fGXNVilJj0lnqyTrYxAXAIrwh1hB1TlR0kaZZyZqGPaACCv4j1NmZDlK
Ue2oO+DKyASMNxArYoQQi8wFlM+eSB7tqhbrRP77tI1GUznmQcK7l1Y1Za4AExkDzFB5MG74WKPG
vDV38K7GgX1zCmd4HELi3kUC8GrvfPpTfz+sNzNpRHrJeFpvPF+XSQJcliD5GbYa7jNM95Cb9udS
8cDojbQd1fSR5MLWR6JRiP1LL0w9EVQ5H3Kq+BhORc2bYs47t1snsctCCiE5Ejw2nTlx/uAKL8pK
Bs0bt5pJjrhfyutnAYcEC0XM/D3B2FcLm1haCnWka4lutRDlfrFXwxWRomQjrqyMKBjFxymzDb5R
AuhFhL9NSOfNKsJfN9143Uy1eQBFWiMo3m0ZQGxOxhRQb1+6hnJ82Uh75jvJp9oHk747YUzMI7eR
u9zCydSIFdszv/4CPVndHXTXLRzRvWHN9GqMEiXl2Oej/6kUt4RWefZhYAq1vIAcm9W1/N+seYxr
ITsEU1o8WpHibi4kzHxSIF4Limo/BDdN3fGOzA46Yv4tw8kPT0US1q661sRTDgY/itSbzBZ1i+Lr
Txb8e9C3eYegknSkSyjzmwlLmVHx/Tdvg7ht4iENVPTdPWexrZ76NDYWdDVJ8JiWvXPk+zq2zuCE
A9q3L04/GJSxLLSzlhuD/+L/JZHQrC0PrhSvGIRsTgEhSo7Zu/7NX3lCWmDPGDXR7FKcG5CYy/kU
aypI70NEKF0zq/sSTFArTJdMtXCBkbUgDVUpmwNs7IrOv2AXAJVmL8qNLw6/Nc5q5fAOCztx7HDQ
xsrrqfUD9VizcBPJv93TZe5ZelURJY9X+DN4ILkvdduswrF3eJ6QSiaeL1KTU4NRYXvCgQ8Etsz1
o8V6JxRIfLbPj0JcvBPFgMwb2qqqZHoJ1OMNZUTluuCuuYR6S8wQ+Cjci3PuAexvd+4H/d32WwmE
sEwqHvxoXkMVtHmjVDw5fDqGIPP3aT9pgvfbxEd+kgWkARSLNrGj7Kr0/0t0hJ2LJXX6BV0LStbE
/xS4/BwaYe9zlob5Mv5pkRfcO6CCwX3KiukcdSEPCJJZ0R0jVyGTwqkvWSRwv2e6WXdB3kSQCZJs
8iPHpX1ywmxRSpuMHbqZm1ZimaQJC2iVyyjfAVbVO3XqMzELsW1thPbBXsb2rH6xXAjxpfzkaN6Y
3TZSCLVhdwRo/xREPkyerONUlRTSbHF38ewwAVH/PgpY4uO+dis+JixvTUOEHewvTpuiXuLlRZhR
7gTqD0Qk0n5LPPahJQ5uexCaQ8d4TZnKiWC17lMVoLr75QAqzHGdD63cEyJB55gkuO4jMBjOTa5g
k2YVmavnyu+5Q3L62I7cfCivCvgMOkwokDUEi1W910HnsbxckjkG9RM3fl3RYaAdzloqbz/dL2+H
JXzsDgEc7hQYnD8PljCpZZCC/FxvXK3f0MpxGODeZZs/LYnOboSU4gUXMaDz3sBOOeEHmu6TQTpr
XoFr0uKtDgZIBCD8Br1vlbs3lsy53h8lGPBaP6jXmUkctYv1c7hdOQBYkknlKdBfsYAJw6UbLeHQ
/JWxvwG9QF3yvjwxG0W4aV/q5rnn3rpHxXNOa/NnJGlDdijZqVunVhkgl0t6hfGqhtjgwASAJpRy
ttBm5E0B/nfpYTPl7HLTn3v3lGbrlEDz00BjuaRQj7HX+iWP8uKuYZHZfkdymf5ijtXpUFzl03wC
u3/MemySym6vkZrHZUorLetuaYeQvP6CU1FFu1eJlKUI8YcG0/O2cKgeYzEr5Edw64xzD7EAMZdu
J9P5tePvJHrxTWCDOxjlqvWFH6DYoHXa2EYjYy7ecqHegyvpLlOa+cw+p5hSnFSq8U5vtGDMlDbB
eKjZHUM9Y3DRfamDYgAe6aj6ocHJBv0vF/AR3GkAMyau3FdYDmvXRTfcxOZDZWzV4lSSMbuOzkSg
xuBNAIkhf30BEt1KaUmo6if68HW02dyNtczfz17vpanmcy/hX8dC4bgESONV7eHtpok4bzPhbJmq
L4TYOlWrQDBYWOFsMdTx0Nh8kmB1MLe2BxBsIRmGIevi/HMzEMDWudb76u5ZqY3pD1iWxFCcJBgu
CPvC6/WwrntbuVKOQ0ChvzYRgqVrM/RaaiummbXqPOAeW6xaNMxWu6e7gjJY2leVaR8X5mC5hx8l
7FhCFIXGoDFr/HqI4lZdFF1A5yFUk4rUoXyfnqcKPlUaU9IKCSNBAp96ZeBsxw3rTDQFOL1JEiP6
N3X2zpTk+aWl57sXeD4qpJ6viZ+9ndKuXSyBX9tAul7cDgQqDhKV0yG+IX5T0V0c+Cm32lj/wQHY
IRdWmZKTB8MSH0eeWEcCsoSl+pZ457K9oAsFLhHUkRkuaXGaohwfpaEK4l1DsTm0RkEG2zlrDS+L
SrYpPQyCAMmdH77YnZDHff6MRS1kb26vK7GOpA/I+ft2ep9OVuolFyf7hmW1Rv3RU7/NKNdOD9pr
FUV/yELMN4Snak6I0rflhpIt7JweS8n3T5/fFZWJWOaAKKD71wTintEKHatnb+SPdUecDXSQOmMX
FfqJ5695HZKJLIDjPeIS1vFiqtkB86YzU+7GtvoUwPe5YcXdBfjxxoOQ0nb73YLxX8S9azxJw7/f
RE8k6eUyMyOedurhPT4gOREM4WLI+/LILiVxMvypJYXHwLVrnT8OCd764uib5beOUsChpKmNGNpV
BXea0zadxLtFhVn2P3DpkGbtBabmCYav+6+2NG5+p5ZE/QvtqOMw9GD5Oreq/vA5YWXKJmylPuNP
qLDY4FTKibHUsYxc9TFUOD+1DnL9VjALSUOY8JlDFvZgkyQ3DT86awl05EVCrV37nW8gynZpsEqg
GgwS0IVo5fExxk5lRO87pIBBMjUfU48HTdcKhB8tEvgPqqIqLcF7WsETr7YvGr8VIoGuvnYMxNAk
zoDtv294SILxccGH8or5RNXhA8u8td+/AlAPRt1MM6B3QN09rt1I1IgkMYO8Afj6dFzEqpPOqaAl
1zvjP6UeS/cDpZo++rNn/0yLAArz0Mp7Za6ZQ4cATU6RDAO0DtHGDyAwei+hG5sq6rLt0zW3gaKN
hdne/1KYS5Eol+8tT7kOWxVrd0mZOlYYqWMnkZ0r4enP2onLWTRHFIcSUltaMe+vPXuBLL5IKe66
rTzP494Zj7NeZcUpvjBYgMOoUkNSups9KQN6r9n6YvfnRMBNITfcQwEaD6kdW4SJPsXVJQINEFQ6
UoIP3+5yMAIlsNRVl0KDPR1w2LnheG+sC1aY/QYDpnGBJZZVE506J07f5RiU8kSboRw4XHfIWGK0
i6UnAmwFg7bllYZZJBVIVUlgCk/wCF2ALdmV0w0/rIjk9Z16SREoW0lmEArkwqFf4EkWJ2KhTrh7
E3cYLRlTQbkelkcPaH4Xj8WBy0XVNIJcytNP0MX9HLYV29FW0I0fz7nNstw7pvw08bpC4zk7xpfZ
POVjwtpLsPXJtfZBMaMqKIk0cmmB67OQfQDHaml+Udll3/4UPESjWbhDrzmoLz13VVE5NNeKirUM
eCsafbgvLQIxs0WNnmrtwM/JdBACr4RWgcCMBcGLbm23MBlwE9vIH9LahV7Rm9/ymlXdkjqEDu2h
tQQ5NxbiJNo2+1+sb+SnubIODEuhCaHf5kV+akbpXN0fSUdOGjTKhaugFTl+QuCueYOoPWA7RGVa
pH075NTKJ32E57oCDm+b0m7k5BFCK2UyBHSKQzxBjtGbvw9luWtjKCq6MuehnbTvZ/eRc53YQ998
9tz1sbEd9XxEOYC8IvgQ+YXBUItxu0vwU3bXyCYsFXa6nUoQfp1JDUZdvo+yP5JKIE8Uv7Atlmzn
6hNmWApwkV+v2xaoh3PDsZRSw0juap33Cfgh6TonpaOeI60Kg1Tm7rn73b/ipoj5JyOMNqiMe4Jp
CmahE/973p577Cf74gw73WVp37c+VL2fbjTN4tujfxMW20MpxUpn1G+Ar+LcpHmQFct1uaozxE8K
hasEZlHhtA3lOR18ftqgbJ7S9vgpPbsOXWIkMvI+XeWDutlpWJ89kkGIQzTV4OkamcXuPfq9MhNL
R8tDXgf8vsyWokq7Ofle7O/VQMsk07cLhU12AK+03J4nSF6gHfVNJTiXnirZYmY5k+p09nGTbdO3
5WJOp0DknGFincSKrcZ4w5e9VAiM383X9CkoyL0m3LAeOih1DeZ8D7iPcfrLJlFk9tllsb/6Hc11
1aiS+VQWeDClBYJf7hkEpq77wq+mcY6pAcEvUH9GZcCg3v0YwpWw6JUYP/eLXgTzIbOvpIm3+I7P
fE5uyofD4BaehWYIso7+ICe0QKH4ZSkcX07tX7k6k/X/nfvWLdS+mQLraXIy/wucMVQWcisrQ3IZ
51bacI9v4o8n10kDDsiBfsYOvcqFiIbAOZRmyiA6QFbWn7bsmvNVOwOGP/0iFkeUMf2IwcJ4q1qa
1W7DGOLux45OtsmnTENhn8owwl4bSSWD9MPuVBhO7cKdcII0/H1GMx/P5xrrlR4eaQ7IFCKCNbXE
X741mkNUcXApoH2bIV8BVO1ECcgvwqxOIvOfYHxSHPrnrE9ynnIFdsXev2de1JBbuK0b2sEtBq4M
4o6oIaXKpNm1Btn0wkwuA6Ya9N4nHWpZv0IyP4hehBB8vLbp3769XGlmG6w8WRoHqvT4GCel4irN
ddd2mE/o/1VbVk3me0V1tuS6XLdjbSlgmXcWHS7wU1xYQoSquvO+BqNzTvogf2+w+A2FVRtc3xO4
8obllaqe+2uCFKUcC7NheqJT75xBAeN5i4Hrqh0PBHyiMUAOEtHn5yIUHNCrfrJ9LPtnteTMLgEQ
pdlGA2x7WXsX6bQHFawN3rZaFuW8Gp1xPI3Gy2H/Ro2FpVudI7sjLCVlO9aH6Gi2fdUE0iVHjrlE
TLpmbHacnAEJeTkfkOg5ETDZm4BaXIYadPOHhurXfGUwwQZGnQb0S5n67zAjISpr/EwiF+P9iqP5
g1H5fHWNpGtItmzCIDpaZvDhhecqF3/lWWWKwrRtTaBr6Na5tCjZf7pHGA4VJ+CoT5U338/SSypj
TAmsHaIAyhiUYXn6sIw7uauw7AmdFZdBYVdBxCHJQ0ATD7IUCh2whw4J05mMcAiJuApqxwN1ZaBd
wDvQ8ZjOllRnZT1k6tGWkK1gdKxDQQUnXuwyvlfuBDHLmaro6Uinee/2r+z6k/3h2wboLgpu+WOw
5ChDkCCh/rQDNExOr7OEj1wCvhnHgtjRtsZfX1AY25TnQtnlocEz1rpcYUyHlsdMx1lzByXqZCRH
CacS5/WQLJ8x7QcF82jvZpluyCEDxXsHpN5eEp3e9WymWF8PHzTNbGwZLW3bE2YD5GA1Yilv3YR3
ALFmfQq090X2LwGP9ZQMA5CzKIq+AITFElDs9O8hN7pOG+jgL/6n7O+sI7T7un/rzpZbnac46tH+
ARiM0pqg45mjEUMhS/RhUgR3EHRDuSEng71JCHfN+lZDBl1Cf9Oa6vZl0IfYXAeQqPniFcP3v6+1
1dCij7FXz3ygNRcJLyyqCbFFp4afV5/YlkyzXp1GYKxmwxox3jq59tppfiZNh58Zh79GP+dEFRo0
iNhOv/ZkodqjsPURnlAjTSQewTOo3A54RWbYLUw7CYFx9m7KCUcDU8QGm0PHlnpmQjp/smp1tmv4
6T2bPgGPqCtcosnLWkhCMKyHtBx4rf0x1DdSCnD15JJ1fDrxyOGD5OgWUsi1nuspNIuK+S4xfdQf
WknWjQ8vwfQZgxIO2jU6pbPq2+xXgmFrLor5KyLbt284KYOAqh4QfZ+L+I+KTvIETWwXM3DHLZpo
mWgPSsLQhqluewyCPwnSRtnghr29AUinXxQiMRev41r6Vd7KREsnVI1IZJqAYXfyxv8RY5NB1vQq
J+OPFAjmPsVyHwmqq43SfsZftSY3dcDhuZZCaoVJmgpE3UQ5dR2CESbSfHHT5m0O2eEca64ZYlX+
kLe/U7HbQbtO8CC0+IMVExK8WbfwFg5tWmgJ1Qr220S2aD4ps0Vw53Sqa8xtlxRreNN0KCF2C9Tq
2+QmAB2FugD2uDiB+Mpr1Hb+Dwll8csHTJeSc15xFJLCPLddtEiScAPJVVqRO013GjKkq0r1y5kQ
1zsilH97m/l5xASKaxXy9G9q4k+A62LQjLec1HkoTPTBTiOmgK50XaKUJjypByWKQVsaOz5xYNod
yV7Y+8+CBYhfrdyS7GO3vZZyK8eO0PDSBAb4ItCbypR+SQ80DutVaOEvVUg6iP/E+9F0TMhi48fs
w/ETBAfzwzZjwL63PXdVIkdAZ8OlwUpEsrtojrtwsVHGS9QNr+aGkwitbAukWAqP28nO8tiVueED
C1ZsQlA0hAxJc29G1/9kTleIwWk0calCvCepwr9WSxu66TtrAL12CpG/OWbpXpTpgn3uOpaW4gy+
1orO3vaRpRAtzw9gv+BfPDvlKMCtVAY8MKOaWiSSnXzdpVHrcJiE43l8fl+7gSsRm1VO4TVgdBuy
quuN4Ao853+Emr/yZd4KNHS1qYBkwxoYzaVewFtHSgTUoTnZB32ANTZW+uxpmioOQUozys7kgAFR
vyKvrGKrOMTwUZfkbzSZLJhLd4IwKee6uGSHxhlip6axvUdhLBAowkDihcQU7zKkTlifIYZhQ+Uf
GJLgf9n37aPu5LAKQ8SQZFa5GL4wiXxxnRu/rxvUjGl1mV52C/GbpgVgJbNglxbNIkxFLHlpA/oj
uHnCIKiQzq/KTim3MJnaTNmW0KkhnHyQEjTmdObaGGA7/P7mahmJoVwZKnrYUxVT/Kun0bFaWfMQ
5Uiakssx7zEJcmuj66p1f9XUTWFzWSmLEkuXoaqJXFKFHLBh9BN6EtOc+4OmkApDOgf1aJ5GAEfg
q8vrtQghYiQMzjfFyIoIkR5QGivJPjX/WKMzejaN5YdG4wOLxpQEzn501sHk+UsBxxAU877gv9pZ
y+e5rx9f2KVkCcV4InlQO5SpRAoDW3+h5KPnjY9wzp3QZplNqS69+eXc7ZOvNzxGNvOBpmSjojwq
7qb0PJxjB/wMG7ORdB/LiNh1ccys680D9qv+d3ZgZe6BprbonhR28fBXhJhMy6qG8el0ES5UuEiy
UxGGzex6tk1ewNLruiA7D9agTgkSdxVuQd8F9pgeOOiepO0VxgUieBNeAZ7ldu7YjoBGpmqxYCNf
rtdCPqCSeNCuTcwbEE48Ak0It+3dPMQDAxfSEPkzA4u5b7+sfrkcgxFrMyA/QgOSjJ622881mr+q
lsXp0O3Is9uP4GD8WJhrYVsb8htBSuz12ClbHRi0LmSka4R486pOjTnExAPtK+UJ3gx2G7Id8gUj
IkljMAlGA5rVdqYSByc6LHVEXwI+c3+sVaIwdmbKqRqlbufQc3SVo6uFa1+tlwWw/zdOnjZbt8Ue
6l3TyxJ6DGxDZGhPGhRqk14QAnDlxa1pSAJqVrHNkYAVa+DCblLQuBqskCV1vrgqEeUbwiAcekyQ
D1hRtt0DJfWsmabTTpBe94ANtS9bIwJf1hIhIUq2dR0qNcbV/qP33MptHx5t5X8waxjHe87kUl8C
DJM79XKt0jEdql1kG371kMYVJq1zpr2Z0UEwK6GZ7k7UdNQ0cp/E2qhwaqn4ZebUO43ibyQ4K1Nv
W0GRqR1fi6NH2xsc7w+mJ1Az7uqsv1OeznmJVIAXIjdKhY8sgnZ5uYfJDFKbjASgok4m5CYDEcdy
d5r/co0j0lVAaTW30WydO0hn4N4pQ0ZdOyqIpaUX+1SdkeMbglWNgfRSijoh6LY6nZ2LLsar0esb
0hEVf9u8iiEv7eGnZuafGOOGZU4IKkEZRezoicZNY+Fw1l9lpVU/mfoIGMRomusTsuGRlf/4DP20
JneuOG+7Vz2tLVRiv5sU/QuMlVor8XHBWS4jpGBqqZKyal3Iebbav/MbWo3AFpIu00QfFEZrnSWz
VjyzGgoO2vX1J88sh8cjGMUoSDR8U2cQKJAXGBjHjCMIXstor2dWq0qRcGIr3uaJV66bUXvgGNuD
IHHqd4hZBmIKT98/nE4KHnWOyIar/JEQIiiIo6EuauTalRxDWKMAWCah692GN2rr8pIfWN3Ml089
pQeKZkgvOJDFJvjz9QMAHbHspOqdgIRCH6B2F/60n1yPZH9/6nIc+4GonZoZ4OtX4zIFUr5ZkBoy
2EJeNNZtaUs1oVFYwRTeQa++UU90PBxuJNWPP7M5Ow6ezPafTYVZ0daSuN2f4zCCh8gdVhMHLD2u
yrK8nw/TwtAGUbU9FdgUzm+Kn22XDsHLLYZTnU/XsdLILEhbnV0xKoNCRcp6joCclpE1KrO1INFV
Mkl7DXwnyNj72tgh20NAZ3D2iaX5Y/EOFnD0XJ6FctnsAfpS/M5Crd8iVJXPBQNuyidaDBcK65k4
e5Z0ZDPyEnxmm4GFauQVq19jV0ryOU/qdw00jyXUilo85ClXE+L6sMPFxHZC3wyXj6OB23bMfA7w
lkQkW8i5XVTRGCdTzXM7R6QucMwMKmS36yzo+Xcsc+PD4oJF1u1ve3zNiAqrFAxSPuQ7GEKV6J+G
XYEsmTLa0Cq8Ag/ae/blaRonvpVDFeEtF34WVfQFQ+Z/Dvey1zrDXkCHiqFzXVcoGLOUfOSmy9IO
TCfDHhf8f544N713oeJojsN77xhyrfRKJML4ymRJTCyhbkarnHXzKWsRGrlc0JdgyScawu6QnCSe
U8Gysv/er6/uTstIj/CSCNzyzyc3rr6YEvZN2rvI0DykCaHdNFbVB6/jhysTXF/hBoxyifD4WmnE
rRGrrgoi8BmQaJMyzms+keN2BxBbZcX5mVXV9G+vJ/4x0vi7Ec82qzv77b97/A2ru9V1Hxlbghub
yN3pIuZGEtpzWmpaJFFnKLCO9JpJoB0Dooajzu1VFOgOLIpvFTyXvm+gsI+MiCm9hhgcXUwJwozl
IDGRtBFWvh+0yQPI2sVA9hWU8yC5HjAf9iEUrF0/nWWYT3yBgVmmeosmaV3gjYngqO24ovT6vVFG
843ce96JlIhD26WRx7j2tq2uWwbomE78lQzPl+9ugEIf02TYS1SM7bKydvAbpjiG8VaDl9lh6N8+
CFiLRVVTS3Ay2+WhlRAEdf7N5IqrWzdgvnv4OqyhIEwIBysLXjHwqUZpOgCZwbdh4pZ/wIwjNHDv
0jwPwVkkiGP9clFoqfL75do6cLArPyTwXXqan/G76PDEWQQTtN22TAfy9fova5hcCNPNKwtZWAhX
Msh4A9aruioROF+EQ5Fqr2SFYE/+tZu0wVrSEM4qYYP52iUeCyjEwacZSuVXIhLCiedn3+3lBuJq
RQiVahnErYd/9aOW+9s6mCirMqJBhjlXmxepGEGAZnuY6gWjYXF9eIaR6WMS9qIeYlkyHXjcWpgm
bMvxjMP8VLVAdeNXzoq1AnpjK+izWjNQvnkDOXflRl1LeBJrnqkqm48gWsKZsiSSeHKnaUIs2aQB
IEjUEDHexamA6XZd3wBLAN/peW9lPsWCM1pqijVroNwVAmtJvde7MUTnCEsAdlS3pFFtZJdyhuBl
HfdXGfQuU4asT0FGFcQxQy2OVUva1UPOt7HdMSt8JaGYiHQDv5Ce52QNuGIoK8jEbI3mXMyAOgKG
t7hDQDynenJR30fvs/sfRx/ZlcrJ1lDLA8Tn7EAizG5+fxV5WteNTo0t87mMzbP4lIcT7YrWh/JJ
3GA597tNl2F4vk/Uc1qTjVk1p2zNhFmv+SZZBm2TdPPdyN/ypXGJUpR1WQs1hgDTL0h5+Bw8CWC3
rKG756hDm3vbxctn/ekQQy0gv7WMcYvHmDvoLmoN0dVbZgrJZu7sJb9/Ps2503HvsVRxeZ5LfBRI
kJzr9GLR1zjAxMykFDABdWbdYx/ZgojAA/8SGh28brs7bY6OjwRdX+n74BZ+tyPf0s5Ks+ERumln
D0KRJhEED0ngMg8VcMfSDqrVRJhIwp5S7Slj0MSeDxYuAzK65zynqwPjMrlpu8JrLxnZb0MBnoZF
81pvjRs+h28bF1DEE2ndfp/z5Lu1hfDIBj2WNYgAUlpboRFVpLS6qvI7IkiVvlnz7HbVWjhlYTrI
NlYItmRhVBJEm7895sFt77AyhSjEJrVqT29TqbCE4+cMWOyuiVtVmIUbSVNlJifHw8eSuiZQGo5A
vDUW9jXvXc8DRcoNGesC+EjI3Qvl/yi7wp4HeN1jy7k8fxd4PG+NiuRbhye6FQE1sCCGR6NQ3WVb
Pjceo2SBmf5imRjvuW3exsjWN2jqCAyW0HOKzFVHWIzzCHRLBk3Wnt8izxDvO2g1PvB06cVVC3B8
IFfsQfBEA36U4ufgV2n0fN2dbyzti6WsFLcmpwanOacFO7VM0Ujah76GGe993MqOlNk+LArJPkB4
eLCQ4IMq5V0cjnK8Nq3z38jfYkRRXeFJFd8F9Qvd7NYK5TVVCnWJ7r94ZaQD/7iyEv1tV8r0pngF
LupJ0IJyPWsSaN8PppISYKtAP3iwmWix1ojB2eVv2UVuRz0f6OKnpZngCEo72dMLB6J88lQ/byLa
tl4kJREXI0ODSCvtA4iMp6Qs+mkaeKQTuM0s270SYsbANK2eiNA+C9lVys7UlC0jScT7Zc3qy4IQ
WL0wmrbAX2H+jtPFPTlQ9dsbURi8hPt3DQOnNXZ3/b6wnfLEXA53bKsrd85kAElEgRBOzOytxSat
oDJVvLni4wff43SsOn2Z1yxhkwt6nK6BH0Of4tdh9h1+kjW06DNwWYHtQNjfz3iSKDao6emMsoDl
VA/Uw50dWqaXNAHMWua/v1v54hJJmImBIgEWZ1LMnrihuOSmgz/t0kytS3zsXfP1RNJOOlfuACG0
Fs09zwRxkt10kCHF/e5SSpmfxQiQWNuynftT5PrGzZDdg4NDzE2ZZjZgHQZ3CzfD4DklnAUXzsCH
pK7YNGlrsU3p/nhfmiaXSgsu1tVXMhIMZZVTRs7lzoZXbtycQYaTEAgIbntz3Sl1AReZEDNl+PHl
sQO6wuy6j+ag4O8XK5uUyYtleDjMHHy53fQQdzr8/u1zNOYZgm1PuCCHdopCGonut+sDBaYUEWch
N2b1wTuVrH0UgSpfqkQ1ICFajlA0Qp/1LxlBV9Jtg8g+bNDb+v6wBRt4gER+wSdhqBIL68CJa1nX
FtwVOdW6c9RO4lvWOB5p8wEai1QHYlf+3bYMpnHtv6SCmHkic7qap1jblgShdS8/nWfXcibH9Dst
2OjQqynpKDtr4TEJedqfzZ/EbR6bCXE0X6ymQ8wFaepvI5Q8tZCnv+L58iaiHmudTKAfejiEJp2f
PZfzM4n8vXd3lRH6ejuY18BIyc8xDkw430vCBTOpdVlkX8hWU4sXIR1vpS82pZ7PIfMSngA+xUTd
tDIO4HbqIA0dYyjeKZPf1vvqVp5CpYbjecUgKmzGAfSzYxNjPGHmsu0Q3jb0+dxlo7QeCa8fD4S9
TRmTR8AKQ1hu5qHFhoZuOPicQP9kYqtqyaUCyvl90uyRBd39iCjldVV4jxiIaqU8vpVEjrTuZl8L
03cbLiYj7IfSCgsr7WH69yY+pC3QiqdZkLf6w9m2PwtloB9YWUMYr9Ruj9WALzZcgg69hmIACipx
LqhKonDnWUFNphOzqd6jNMv908KYZzOJfm458vPl07RNr6+HYrr/J9+C6WWIukfKRWPbIc9JNUvD
QjtOk2ItX86z1qWuAmwIq0H8hFtA0+QIExIAYxHmqu0GBwqFcNacd/jGlCJAjc2fGQD6hw6lNn+C
orHhlzOBmfFF4H5NkDwR163URqa4PAQOnKltzBldtwo0ZZBC2tQj9s66FaJlLy4lfiwr0ADggUTm
S8i/ltYzs9svcfezWYCGfumRi2eGPOQ30wNxN3oBnEGRHFJDB1Z7rYQn1SJBoVVSSdLf98oI+bzd
RJ2H/wkywfaWV/jxrI7S9oVKLqr8MeBSTcg/bHq3g4saVjXUcnS2IOJNFwAe8PcDK7owX/meCkLU
zprdme3D7+tavDW2XgEM8wI2h2DeP6+oRDR4K6nqqP9lceX509FWnp22P3oLoVXi7TZyBhji28mI
ds9DqpWr9C2gl2Kj+0fc1dcYjQcaFDgEbCIJ3Al5cHZs0y0r4uxVRa7ZRJtgEKMe9LKbH/KxR62S
swaV/VYdT4LovAn7u1Ogh+skMIa6qP/y5EPU74Ie3e0PQkUbdfgQOr5Hmrf+62ewbZSFwB1wpzIH
hqxywSQP5lsoQ4GOzanOP3GiVMN8+wG5ZC61IBXhuwJIORhw/IUWFETB2WF4jfeXP8TTgBgGWYzn
IoMoBMJIEz36S4FP1j0XOmYl4SrgOXTTPG96DC5Ix8uAaxVQRzYw61IofG8s8iJbMK9pIqoDZ2zx
eLCleA+5JLPXpgCgP63wEYVVjx2GJGDUPLYWw6lKBf3smwLOPcZMJzfojNtFpWsI4qyyTCALLcYc
3EVB3TvDPYISrSyyI5Wuwn9EnjFYOm4Jbeo6Zorh0SWaYcQ+F+NaKdvhZBS738yxqUUu0c8jBiWf
0ufPQVPYP43Zmr46rJNpdR50NH6RSqorsHpCmLDIGIOT4ii6SwhL8jHEAv1rkst3pVPcEnyL8sn8
x+Gb4LLtKHBh82Zdzq2oaEHRjpNmaivfii4/eXusBEFpSQXwU0/qhn/l7Nn6xPhEKBYytimc5TUg
M3rGta6vP5txCe0StiPkYf+7vZSfstZMYpwqTnS1lNLK8qkTFpkOby9gjU7PeohZwrQgiXK/T9h8
lMJ/4ektUIU5Yr47wEsbVOK0EvKkSy8NyDIA0OabEWlC7rv7Y9stMkAxPdqxHKBKFjKvxWrU7fi7
goptcuwauobtOEdFNgydZYagycgO3CkkeNEZdGNdN1VjrAUUaVK+XBdZgt8D8x2lwjWh2YIUWcG3
9pCF2Aftb/MSxiPUxro0Gg0+4+mWvMLfxtfc2ZG19A3Gpxqq9nRb4O/t0lR2MUxBjcLsdNy262i4
OY2UuyjNnBsF9UwrEGJb6gluWv0fqcAGs5h6T5B9RrwPzlqjhaADFWaM/pmYxRZk4VLaDbIEeKxY
7KpSNEslBjQJ2cEicTdp7MKONPpNdDPJKsUVIidCU9f254mUrTGwy1APNXsBo8YucyS7q6uAlzIN
fHjo2LN7B27o3FcPOkt50SfetXVVAWJo/FRifvUKV9XgQQ6jS7bMERYeLkeH1i9F9JQA6sLU9HFR
mcMARJSbaKGq0IwI3zbsm9WBdWpWOK4TholGML8NV4r1ztFAsUMBa5cUGr4M6BAQanKhwrmqNn2Y
TUK5Unn1FhDagDL5uRdlqoL/xL94sJSXtdL3xF+LeuihY6xjCuvhnR+9PJRUC+Ib8BURAfjuTlUy
+BkEFYaqb2BWYPpC3MleMAieFVgYjo3DKeRzTKqzDl4ZicHyHoHZMx0besBNoXCQLy858WKjyI6u
whNS7CSSlDYrnZAyd76kYwyaHcCf8MrXgL9meSiogD/8TDHjHOZ0eo1Jjj7G6iolgmBBGCkV154r
pjmsHOtA4jDDQC+4o/Y+zHrh7ABlCretgf6rs0wH7BttouKStD+AVI0EGjSdv5lGHtBt1Z3N+8MD
rDvwocDG7MworM0TzWImSYiweRujwSQ5uc2xDj6zS3d6zkOMSNS/PFlV9Cq5iwMkCO9OPSnlOwTz
cdyaq3qlbcRLQaS/8D2XoZjEodu+Z2L2dAf1miqwYi/131JdT1smHIBFJY0wy3LGcWz+7LNg0MCY
XonO5stxzakHpaj2PIj57jHyUklnokw72L5kFJAGDRelMTwI1gZuL0Lu7+Ew8CP3UFpCF1CPb7Sk
W8yYzkvS0GMIRPnB+zkKMatMIpI9qKX2rOrKeVEhU+6Z+l78HTcEFSoEp2qwTehnahTTsYjsN5I6
rLuOcQqIS4mZJ5o0ZrnORKM06K4v25ujPzcALq77UTdVwdqDwL1mdA9R1yZCQPUqrgnvAwfn4miz
M00vLEposWNWSws88HJP61/P/G7dOOG41IEOTBXPdk3t3PA72TEDvichEmVzge7UaWGnRG/ct4NK
7v4e4dg21cXGN92HvfzUG7tzV9OOKIIzfw//68e2euVi2uVwJgm4v6Kwuqe6TYZjdJzH3iQIlqP2
/EcCypnMRPNrwmFJ8QLXHWfoiu4yJ+8GdE7UHRvJkrr3rj/O0p4ZLMAZficXJHrXLT5H+NEZyr8Y
FkqaIjCwA7iQ4dwejbmJR/9aLQEP/tIZYRYaNvLj/jCEqQCxDH85zPkTKFP1oYctxiaULkA9CLLX
lTsknwNHzwhH9NHO/UvH+mCI/ncq6lgSjfQP4d/ge/C+OpuEsioSETm4Hv0FrUAqb4X+5KLgIBr/
oDR2rwqiXi87PmCLhbmBpA83mNSPRz+Q4bRxAwCIqqWORTg9pSyrWc/FIyfeETkKktmroYDqU8c6
f+JaJINxmJ5oYKuusoR8w0ZrXtDp26UYsjk8rjNjqUH2d+Y9PGc8wHXlHvvTLLTCf5g90/ch04Mr
K/6/hX5WRD2KuJaB6EfK/PJzuDn0tRcUEa2PL8MgS/v8GbbV2njQIa0+as0M4raX0GbJGKRoBWLj
MJYQUJHtoFndyyqQ1hjiHHNc6v15Y18ZjKtj6tpNH6i7RKLDBe/jK7D39US/s77ZsMHHfo6Q/x9v
QOeItKET0A1IOoDFswtaWLHSXmOg//5w4rEPUsmgwFfr45hJI20y2q1GdU0XH1Ms0RPaQGp0WAOi
B9c6omXw5An5C2EjcJ+tJCtmkbMxVUnaBzvpVtwRuSO6GzZRyYySrknH5zKBKdmqnIekJDBzG6oi
Z+aofWx5kt40vZ1MrRemQffeI6pRIdKGUiGPG8rI7HgBTPsoYfWzIBkh4xsTUkoyok+8b1U2sJ2e
1nyn3r5SpwGxgJzfL3N7oXZ4x8jXGF6+dZAMriY3oCpUfcDwSrTqfsYzHxFBTsk7BdWfRCvPHcMs
6nbhKLo/0pwKyiX6cp4P3g7TX8nrEGUbc/AWyy9NC30pLidfojsC/96cJFOk6iMzWJYO3Hnzn8t5
lusL7mBSDHz/OOJF0D0DXVxAAUJHtu50Bqfw52RfQTpNuJBDL9TqKDPe0ZTOm8vq+JnrWeU/1/Ir
uYc2gUeJrQeniXpqX2uEsTK4ZN83AwEpOMF3xLZYd3guJ5yzanh8AUJus1zkf+7KJ93pdxYHQpaL
f6mzq7kthaKSLIp2xXxJivoMVL+sacEa5QmfDWPvtrLFDlKmPkcya8jRQj3StBgBVnILlsuZRC76
XUPrmvWpuoJWeQyCQBX8xeKkMrwgV1T7LXKBrMAhHX3N/k6vJJp+bD6Awkj2gsPoVgriv5CD1ybC
w0red+NUbCWS2K3FpfFKIMSqpRto18Blsl/NJwalCOi59mYSH9PJAK/HYEKw/wa8sGWXg5/R/cdM
7yAZiOSMwDShPSp3CPbXq6Bzj9+z2fyQZNVMPWHk5jxjbzEryXRkq6xavqj1z6I9Zsg+ct7jOgAN
PXTf9GNA1IST1xgtsM0W3Z7wZWRMOygfQuKjuoDVN1A5jlZLne6VeQGaS6/fCjEfHNmOQF9dbhMx
SU3X8l/rsisDswxqVCc1h800M0h8D9WmgNvaly7zXzqHANXg0pkWAXQJJDnuRfs10+HLkqJNY00N
EbUU6ZDgPsRYrIbR8InSoajQE2sOZCYt/DWtzKdo/z5H0rPcDXmSX+UJETq7301smpODC18NINPv
L4fEV7FO06By/qveVDoZFwUlczBV7uRSc2b2ccVkHKVQtcdaMf6jmxUjbuN0dJHDBQyO4plOG182
pOl9RyQGa3prHmde8q41aBmQFmhC+CdM258UsGBjuWAQ1vQk9zMBdu9vfbDPdPUCumjfkUtJiG2Q
5odMr8IndXKRRCYp2/dnxEyT1GS2bH0ohe9xOPfdmveWJAB5x2rlpFI18ss9N76xKgtsD1Sf4a0S
0B4xsr+Q8MB28LmugFLzCZTnj31RBqrRC9fCyZBJSEq6vFciqBGzA2X11hjRaUUYvwbPWU7fCyF9
cbqWZ1ojgctylhf6NekVPVuD39LDz/iMe7foWLLlk/djE7QFqHoTTQML8kjPbxDgO3l2zu//sSig
jSqyJYEyfjVglBfWqhKgDzxoMmzjYblGDV+vtmzhZ9kMoW568t2iW1KgmTF4JEB+EjD575Ln0ijn
YAwUQNCC4P81N4no0I4SNLzDRZp6KCb8kMqKHPwB3gZ4JXavcjJnOQcFJDdC1S9HgY39UaEy4DnG
KaS6ZffFz0mjW0sv8TTYqnvLd2ZYG0YnDPlA9LgQyC5nd/Lqu719emX+CR8yU1pUV5rnBoxw7Cr/
03AdPs3uZTu2Tw1V+FZAeaDdb9AKsLeNFHDw1dgeCam78lAkp38NksGmePXELyDmUBJOnh2COp5t
MKQid3U1UbufQSH860bwuA+blOEUahWbsBhcxm53AMH7IzkJFZimrQTvczWqKRR0xQcSnnd/VVpV
nQZY6Us6oEgVMRfuRSeCvWhweVujkvt1X+yMDEm59zzB7Dy9lifwA3F4jDhfK25BRszZ0IK0a1yb
/xQdd2GVOrLWSDhgeD4+BsyuAv7Qpsq5LUfOrdm1N3wMWbIEqkzxuFNs8m3pNRyRGj5AGNpXw2vK
ClFCmlHG1uwNyGm6WNGvi2F3mgTnNtxb06zBTi6jVEpUvWG1L/dggMP+SgO71LHzTKHB7dp3j2z1
JdH1fNDdWefRBHNGAm7Y7S5qJP1mrh1B2ArcNqv9Lyd57VGT/wMqHGm6eMD/IlSkhqjfcmbcSDv6
yRVLPhFsbXE0iCUPjoqrLX00ujt+751P9EkdK7rbAje4hcun0BJYzwORSoExPqYM611va9XmG58N
mQ2Larzc9Bqo7ntHdhe9ValssSGa4eAFz4anTGMYo2h+u/6qoYNPU7QmE+afCAaHBJzqzSTch9fG
NscSBLGUZ6RVHPHtKvvplaCV5ymr1wNGtElrWRBntCTzALDg4sTYNRr8/SUMLFYRRk91aBWKJHGH
NJwCtJIsDR9WrsmT8HvRx700e/jKidvjJ1cjh4iFtLzEfVLESfkYpOuj5V7sKNi8DVIZwA0PsjKi
2EvSRyHPIB1/tK34HA9ep5uDXQHrKNqDtPet6z4D7dBN67waVRQEuSv10c38UOIPlStGDuh8WZkH
cJIXBd+NrIU5k0Ua+sQQEjxLFLxj6PUT1Do7CAOlQO8Fn0ZxutfTok+8BW4Hw4Y+SvfL80eujrmo
EivSzfARBVVzFsijcM5qER6ZbsBcEp8dOLet97OhNcbRHiJDo6cGj/gh93tYzpz1VyqIumEb756c
g+sAXSG845SpOqVDIPrM2RZA1xLSMb10qxMg5JD4s4mqzHs74cpFzk7ilioqpo3Z7cmv0ojcdj6i
5d5Xoc7OuYvD8QsviU+xOX1AH5iAPbZiypne3NbthPSBx2qPPNK11+OegSVsRk0h+XqLE8tkIppP
2wT6aTGVhYSbi1dm7MOF/AJ1dNPSarlhuJEK2Z28sMr9LxAx4P/agKI1ZKfi3CvSHssqUoeUaQbX
kHECIwkXDCJY8rEybl1tJXjPwhys9rHVwSsuuQtawNvY3FOnORM4VZI5L9TH2n6DvUArg8GQRZV7
pVwPaZrd4bp8N55b5sjHT/yUEzF7JkUOnqVNlxEw9wpYEp7IVh9s9khkA9l3P3Tt29YL6oq7WArI
sKjNf8K9Peg6r/sr/h45LZvYtq0gS0Ai4HCwwP3AX7wE2GD+ipg6+AUR+ZtJ8UQ6fyCLxQaOvae3
ZuVid2mf6CEakjqMLEdO8N5/MY9zPyqngwfP7U8L0/3Jp+oWCrRm+UDPcjzFutcw16mxeM0MCPDu
oxesUbonuQSVXoq+YlLLZl2etWUsLHyzcSNQxgy9/NUDhsDIj4v9oqbfPWkzUS2+kOEvi1JMfuJT
6VePWdfYaRGpq9IFQiAuVOnliyynp9mlQAdivpqPFLjIbqLC2z3FmLg/j9aD8cSwank6ijo7q3xE
uo72KYgF/43QJId2Z2uwcP1rU1eIeA2fB9JltFEUsDZgY9bz8aD1y9+IfkD+EECgTKr05erAsnwU
e1/yslMmJkqvF4KyEOoIWyF1kTCSWtz2AgTUwHB+KxoL4800z9albRLYAHURYTU1kwiB/NbAGxlW
/3my2r1Cm5o2Wt3TCgalFooEtpsM73Bff765SMWYrkaU+J5VDV9erdN+r16PS7WefEtnmAUdnYQN
/HpO/B+qwHJb2/q81M2V3NnImcCnZKFLSQgAuAUNbZtxmxbj5jw0x3HSXgG52Svw8QVvJEJ8prsW
uEqophGuhoFDtOaIOR7ECbwkBtvMzvvIcJ3jvufKbmI5oj+szB0ZzZEYzmtu7RUogN8nHJza3HG0
Yn9KhFNljL/PsO3GLfyW3IustexwQSlxH2uFTs4UqU/hsLFwM+IahtttaNb19x1aSHzKZGPJpH7H
YHnVgM8fK7ksK9r4EDhYXQE2y5IiP4AVZvu2mB4eYEKbggnf89xWpuhkMINL1JCOsma2sUj6n6s/
wbw/hkhM/IamVYH/sCeCgkXbrhHDoe+hRID4bAbOvi6q+wy+6LJSmivFnPzSFhhWXkukYWKAkuym
F8gE3bH4TsFVYkJMfJyiIv7FhqSzxZ8m2zRhA26mFECsXAmMe6N/r/GZ12sNRpCeWh4x0gzl82GG
nGBAzQvNstpTwIUT6idPK/42jCDF9JjbOBWFdfE+YYg03yxInaS8oRvQNC53T139KanG9XmOyEY9
Dvjmn2B1cKVLW6NRbHlIMmA8BPPHMZo5KXFNAybgFXLkbFf54iIQSBq/6G3unNx7yDk8xJYuDsQt
Rq47q0SO6ecoWLnNm+qlXSgZLqxDWPna2pqAC8QkSK3+rRoWYwujbjh4ZthWih9Da8SGgwCyRSUT
k3vUtC8ylVDDFtPTwwiT4QRMXKBuYcCg+sd99PSUEKod7g9K8Agh1uMY7xKq3+LNst1fWpw7LQ3S
1FW0PtIHu3Q9NcgauzbWT2ookrMJ4wAcfycELgsOVM7SYKS6K/wpNtXjNUsm7e5GUVl22fWcELIT
GCaaI9Kb8hKEskIRTUGleX6Hm0hVctjN76nmY9smpCQlfuE9gXzfNrrV1dnW4lWAmuayw+nAYM/B
yjqId9ljhso12CPHhsiCWh1/3h5dniPYgNZLQ/Ft9sOR3kBxtjDDlf/db/xlszAtRwXyHUQE6QI9
refbWiA2uerRPcevkAr63ZiRh67my3csC8adCbrHkky7EAJBlKCUN392uT2HIXR9AGz4iyRHUL74
0DEU291CPCh6UWdUKzHN/ak/6uoY9vPzlo2X/XZrVnpkuvl/hcU/16tPn0wUBmjlnpHFYUCeGM5i
w0QrSlrgxuo18CxXNWvXJNv/KsUln3wNlyavzYgJT/zZRznhXF9EX0PqcxubrZEsQY5+Q8wdIAYx
dEH33CuT3qNRZ039PexC+qLFPfzRcz0sg7veNGAdnUQiN5SMc1ihDnfgBnyYVxRWSFyWFVI+tBQI
1ANzEKh/e3WydKb8pNoc7pPhEDWrsbjObSplWAa+F56lQyDi5j9oaoJtirXgZirjXer817uh1/nW
kPywc8XEjpTirfGgxvMikWhBrjukQmRG1k0aeIrtGv/pX2kQv3S7wEhjXFubQ8aGnPXRYxAmnrhr
5fBeFa3J+PjEf24RxPvIUlFHrabxJrqPv3Mz5+BaY9ZpB8KH8JFJqYUUSYAjk+l0RsHrQLi1+3Y6
+a0qgPTRY1g5+MHSrZRULBsuH9T/ePsN3k2N5sX/ulkPe6EY6loo6uayWeXuniG407d0oWLevAoV
NstPAJ/PVNiOrV9TQEm8z/n6qoxRGtiOCpq8WlqB//MqSmnHogFyV6+Va83JAQCL530WzxPkp4//
rd2w2HTFfkSVfbl8j6uo/0v3lTgTXd2udQYp23mjhnuYhcIEhoV3BHqJMO5uEL6EmKerEMW0y4rL
pmYk2+QeeP2fPvBT8VZjTSwjPQJLN1Ue3KA5xXwGwDLC8LnzsNQI0bnd3K4Ea+u0Pk9kFbVE54sj
QQuGiTJlBMlxBF03TzCCqMcz6eXtoh1uS8j4T9BrnyxYZql0Ip8b7K51WvrBjGeihaEAKPUTozV9
+qQHVRisMcyuL8novHOIiWg23bo+6PigFMizXVjvm/17ATndVSUJ3PzljEtoIuWsYTeRzg3XI0S2
99DieUxsTNbEvuwp15HZxVmAnTqBSXdj7cf28J0ALrNaL8DcG2+QozHo60+7pKYlvHRvR5Zi050j
MmKfBmWWrGxWcurg9yslQ2hI2LSDdRf3kL+gQppZmj/N0xP+J53V0jj4fapsaAq08jtZp/wdz4cJ
GwwbuFnGkm+6KQGwShbQK/PGnHnx/f1XegglkAxYpyVEljBiD53hzASCbPQODJXI1fdc/+9hIOJy
ZJ/BWh9azuapPNqJN3hWrBQqzTf8eQJqqsBS20RmA0YZ+nTESEojk25n9St9GK5bLuJZCb12bB/U
peyzz985ZVf7YkDxRz05ukOaH8j7KQwBtZcxyvApyCosphT9kAo/sgBkpJ8pKbKwXtYPMPlWMDTO
C5rRhXcS0IVXMdYSEgLt4C/dtrxoLJwZT0PIky3xgHvfjFdCULiAY7sU8UTGeh7CgcQatMf41ckP
/L2LUin/FRdaD1mx5J01BLWZZH1ejTK0oA6TtVo86tcojpodzIp7Xw9WnhGIEFKutTfPXXOMxZs5
odYBkrmb+m+gc7J4XugODtw4VL1og82lP+OvQQ1IgUJKmMRZsz2Am+Zw8vxIPnmp7GnXbsNcX0Je
cZDg2mQ0xGTMDl8Z5ArKpKuVvxIizQDNTKxvWsFcrmodzDoYKUORYK3rriOc2OCYZFRz6SB75DRa
TkPi/d60Zpn5OHwJxmWoNmYc0GaGvs48y5Cxi4EUP1X90LYsOEz0wtnOBVX4WsFpxKr7HmRoHCOt
Usqr+GIXMzV2iY0GgI3jjhO7ywVcixnvVKfZT6DG+D786YgcNbCJ4AheEL9tBuBv1kagodUe8OsI
sWTZCl/AGM+HuFHBuckspZH7LcQqLlxqnInldW1PKH5T96unzCHjKYXzbZ50/mVGL5GoQj/zzuac
YYwqlJATEjNyrEHai1p3hOdB1bVzj3qVDlGkHagROTUGsyYugp9juI3zXQ7FrltYa8sW0meA/pyt
FGfRlLDMgqHiKyW3m6LawYGjc18gaLCqJtUhpdLUiIBiCNGsmffxH6O8FuQEb4yAnNJMmFqwjMXJ
AxjvsHGe/T3LT0NBPmNZp06vnsR16Kncr5ec3dXEYUyZ+OsexYGcDMzQGtCWq2bVxwS1mFYc7XVF
6FWMzBE+Omqtu0ibj2KsLamJhEmoOlpbLnTKGxQDRsv3EYy1p98VoBQyMST8Xr5tLHXmm/l8d0db
tBxG5W915gMRR9D4vWDt3g9IiQT8MhPDsssTDsdarU6VTNgS2Bx4y7AZSvgK0R95S3W8+1Tzxrxm
bK7JjEyHRS4eCO8ZnfDIArrHDoekPXRMZioNUsz9yvMwWxXsxfMGdsLPE8AxSyqAZOHnBct1Ws01
4dMZkul6WXMUpUfJy+GEyAHkrR8OZgN03xMOFq9kdXUfIxCCkh1bwa7gN0g34ikLkyi5O8x4AI6N
bCl4wFB09HeKwURWkB4yV4Sj1ihk8NnlykFdKkpTXMmLjqqyBlQ2Hv9a80ds8Q2Y7y2kG17HAiK9
s2/GlIBq1UypLTg/t9jtAro+0y4mCRGQCoLXnksun1eDQsV23sXkOiHiNvjxEDSw0VpeWFaiRp0+
hC3y3CennUpC20fidwDCLd159Z0KE96CSw/lcbuyvupY43aTcN8mga6nVGwngzF9VsrPOvLI6M7e
yfz4SBkb/Uw5p+nqEujO5/8zUQo8H8U2nffHX7A9edPV5l32lzy/juXy/vGyVk/t+KTIJ2hUdzWd
KnNbvcruCAy+Is0Vo+avUWc1Bfh0tFbzWJJj6dSPPJunQjQp+TRNm9/Ahf+UOYnVViRtFnYeeA5z
Wx8XXwzOcaYJYbX5kI+7SlWbWg9lzKOJ7M/6zIsugshPUu1FuN9TBAIxt6lre3kbDOhR2R1cy6pn
c4L7cPOAijgwe9AUQjx7dlCba53so/PUv9YogsVOLwCib2Uz68mI8PJuDGD5ExLqlB7ozfaT/+jh
XaBuE+TEhaLWdD13s303L1vIlRriRdqS776fYckTHrwo/bdpA9ixyVBdBRnAf140hxQs0G7Ab0jW
84jqmgkrWRRTFoT71GaO6JURNpAuGpWFmNgl8q9hcYAbF8BU/fLz+iCF0jiZTDrsAt69WiYlNeoL
aZ/fBFElkgqmnksrKuSsRCI4OC93lH2XPW2CXH7SEhtdZlLgtG8eDO8cUUp/61yq6O6gEani00R9
KwcxZ4HiZVFSNFQtreJ3ZvNrhYWAvTdlH78N94P7QygBWuNkQg1N68x5fuYAEm3u4SnapZPtPNRu
84YRDgotcb/YBcyHMjYCAlzQIz+E9eFXG7HbVzF11B+7ggYj+F/K9v1Qr0wdVd0Fj3KyzVZaTWeh
mzj0iQU8rsh6N0mjyCXIhaHhnQ2FHown2KLGyoe4oVWisHmhUmGkyL7K47awuAFOhCrY8gr167vT
Ic/wgBQdgFX5lnSULnRCdEvGaoHscrfy3HqlKS2I4M0srvebry9NHqyLmbVoBI3dchfZBIWt/0nU
rER6paV84xyyL7LO2sQpiqX70mPJkTMGk9Zi58P1jI3n+4r1S+qFnnLSJVjHL1siKbo2k0tFfRFG
0JifYZMgQ39I+AG2nJsa88klxXB2S2Ry1AwN/RQlBlPsDiVVU4T0EhkJfWvxJHANVSZ/Li/K6Iae
LjzKuskLCiye7TzlVERg4huNeKQBCIiRyZBSgSv2fChqWldZcHofMsHJ6wjaCcHhs1RyvIDH1IFB
US3WAo66cQ8JplBnP4CEG4AjnhH65j+dQc0CHqWuldumis+DjXcBwrJoYRJcacxQNXj0NB/dASbN
lPfVW22t2V4kOcnlKNpHlNYPwJ4u+suJMk4g5LrAuBtXvkF30XV3WC++P72+aU3PJ6jkcJ63rRl0
nl4QoMJyXm83QqQYl7pP80iWohtVxmrmzM8CzOaKCrinZEtc4XwuGx7XTdPebcuD7lt4UD9mgVCd
Si6lOfaWWcv10iAWOd2egZe2BkSvv+MecdXenobri8/oWEu/wM4dfT5NzsXSFVr77nzOiSlOi2Pw
dm59DmuQTNfSwzQwsrwANU8f7sTyJ6uSDmMhXxsJfEfVRtgQ/15RjfFFjNdV4KmapGY2YbhltI76
IhGYA0cdlpk4uqqtXRmcHm83/gjYYy7bqFAQGM/hhdxID2xNbLPYNImidIjcknFLynJmdqojU7Xb
oTiwE+ND2ihYtGQQmYa8l8qf6hlA2UEsytVNu4VsHPvNpA+B9J4CAuW9jpCnhKOJScQ+NmfsCu/j
cOQ9RywVGe5TAikb4M/lzTO91GesVI8dfSBTvzrqyfPY0ryqCvV56A3ehozQMWd/Gw41bs1xt9UT
Vg46RxOw7kRCkZUzPeXsTuN7yxa5IcpbwOc838vkBJVmK/aZI7NSYaScLWufK9zDkAW+krzWAll7
nst2Ce6BBRGc0lXzm613NIHRQXwXvFaM/WL522qPx+UE2Y16vfaGCKJg7mmAjfIf0SQWWrtIyNXS
r6wMX4tZNzbIa3Mu6ls78XDv6lZzryBX5ft4aFq8Qgr8ajhGId/DK8C2RcnaZv1N3fcyx43egy2q
utTOE1nS0W4yR7GmSAAfpwF+jhK3nlt60AlB1yOFMFuCKa5JsPnHB+PURjwyJfBwdQxWputqbioS
dUitbO8qbzMr7ONSsf/S79jPH+Af5AqijasBkwQQANLlwClXErAakvg3oiA4KTuHPkY8hYHvhOea
dZDadhjMuuQ0BJiesv+ElpX831FhqcO5yVstCP3Ug5y78e00V93eQ+FNqNrUgp9FgUmK/YbrPvm4
0Pl+jMVcXYhy7PWkhXXtlRCDnBWWn+xl2hNKvDXND36z4fSXLuecNhsIqG9RhaKsYRQ6UnRul4X6
hs43Nnw6UWnGZcKtLqqqi1v+2NkA/ICjwoZ6cwuzu/nC1SYrdc15VV/0mwYuJkJSf1LtsIOv0hIj
6si74VBx/dR9qIHsuAB1yYcjDMdl2mW5kAgaATLcKe8toxw4GWxp7KWGFhoVqD4JC72RAyYk946E
cqGE7l/7QqWL41j0DHVT/kdCekNA4aCqo0mFLjKuVcLiL9gomXmUsoqETm6UCn7HLE27HF0J/dy7
n+xap6FVjli4XYvkBXW13IJicjfqGxS4qFaH7FaUcnCzXSMbXBCPQ3co7wmmgZCRXCYJ3QnB7Gq2
Fl25GT/rhbW0RV1pA8RLZOsAX6Rm0bjtNp7cTIaJgvQyvxUozl9FxkqDyCQ7InERDP2x9lCoKc5w
HcYyPLE+sVlFeMzeg7V8edxuvdUrFV0e/yZIQ7kiOpOZUyRxo6ccbaru1mBlquHVVT23ZLQVesdM
OEDwbKauycMRHdu9QpZXFCgOt/U+zvpMKPSd9nsl9FQwM39HUXiOYOADYfggUeyx/r14huy6rxAV
FXaFEwYYb9O+8RAtFh8YqMcXFAhAUd7kG/Xrg9EayMsjHbfSJ45GIGVyUABWO3BFXerM4PPv+NA6
sui60kHNGE0mXEuFx6Tnmhgy5xAQlp4fdsvbipdBU2JG86gBtR+Ul8bSsFTumUMJpzMFuovt9mGl
vXUTtDD3a+S6+p3+zOMT7lIIHSQ8AKVJswqMpVtyMktuwG3awXYpWC6ZtKgBWmPOEZLaB/guNZc6
pr5NrxuUjiCzW/9UElTY3sINEGE5tZ/Up+Dr4CmXCvvkpSAv0VTcZowngjkNAWCQC4QvmrkVMArN
X3rLyJshy5LCHbxvJntVSRbJNVlmc9+0bTo/aQ+vZWCIJrpDTf6ExAx0kLTXE21Hf5MmJJRYXUMR
8s6flwEkwRePfj6OuBYorJsu44zHNbRT1v8IZHtW0DoWJjPRqN5ObutNogLSM6KJB8ZsWSI0y/N3
mKhXe6THFkEH/4BtrJudA9P4RMAjKWbP32dwc3mNHczA1efc+8RQ/SbSMBIySboONHGM/60fnzDy
6SOiLYHqleOYFyzMOoZRxL0HumaVE4ulsPp+8cjriwXLa67DXTo8Axg79Y9RJT+rkHT8hwS9xVwW
TdJcO+ezXmtrohIzYXBODFE7EKeAjV0U+ymqQ0EzDTb5DADHLHo3MUBkAzSX41vyijtczErbXAzg
KlKTr7HGQqTZ1osco138TnvoGp1Pm5PwzYj5kZppNHmhRpp6FkiyFcHliZBRPKqq9CX4LepjKMhk
dqc/ZBrUAbrHP1wa9gEk98V0zkzVxLwRvoRvSrTw0pVQJc3s7a5R2OVKm25Rk6ybZUP+elDmdDeB
ePjGhz5dTeCZ3uRUfvobA0VgiRhJB2CwooA7xFkjtOlJnkXQ8AhpEpELcUEgzVAc68vPtaeq6wyv
yZS4dMGfjqBc35FlLdgyxUHZ1Ux/ZrEIUFQgNxnQTMF7b5in7qBMR31pv0mlnVuWJIi83Zia9PDW
fkVhZgzyL5BGChymReaxynfOOpeUr/bBhA+Unb+nxXp6esFexdLpYXVWdtsL8HZqbDFQxG4M75Bb
1RXMVfMtLXx0oik6xlvMI9lT19wXByw8qwfGMzVnqQ/EX1xGXyHCU3YqrxJUGK2vw3gCdE+Vc8NC
zSx6esXc2ZGeJpngvB30NstyrqiVHZsO2fMNAXNE+jmWpEIThKdNFPvl91fkYETVHqS0HMu75IuC
xk/1cCrGtUmgPvqOkp5eF9C+vI1rpHTGpCVgKrXRgHHANtG/UasVQ6icUZgoK1pEA+6OH2Vct9yW
pio7Rs4dk6kEetbGDUdNymF+86Op3YCMmhjeX+fIY1Bks6vdYLJz9toMsFUvrDbmAOC9Btv+/IZw
KyCDiTQiRoGkfOXdfIsAJoludDCgpu6dm4Gi2dZ1vJXKf7MCvhbi/5oYoIDnUrIhrH8TkMRCpRhW
p13MFqqWjkfw+n/QRCDtzdZGLi4KkHfCRZwG92Y4on8jmOXMDvyeyJ0sOG7aymEKCv+QhxkWaMo4
8QDBHpGQgb62r+O1IdRUrtpQe/dPLoK1d0vIVRp1x2BnZJX9BRg2uM+SSS5lwwZzTCTaa5OVzcsH
Ynq9ZtdcF9aBgy73cNUgT+r6wXIZHCpt/+qmaz2spEE/jYvdGuSS2JLKSXHjSvc2jpxVs8XnLn2a
DK1WN05nIDrhxO6O3XDifAi/Pf2Ojq8SLDrnA8uE78FilyA1reBE2JEGM9snTlzLvYOeqXJfoMsU
xTZLnbUMeYLUp2e/8SIn44G/+wltQe2yzqQ6hy/alI3tuMCmoMasH79Zf+j4SHJ49m5dM/0+5v8w
8jHJhuR7CmQkg4urnhkYGXpMPRHXkvltLGMCRWMjCK9uQhGhSsPQlOrI/CanAh2tnVHLf+stwJ5A
/0Fi9zDGs8xFM1mV7jhHR/aOWR2aNDGmMcnMXMTZKRmwVPSYG0NAxZyS1NJ3ZqsAA/2itohUPJXE
IaYUapkDk31bkNdvhr7Vhz3WDaOPqita1Kr0rwkxyE+htCHELiMF5GS/MiQ9OADmKe+lr725GWjg
c4qAl9e9zoLF0fP8d7GMhMwWp65MeWFl2BZi2DUs8RgOH9N89GcUm/DswADCz/nnfcu22mGyfQUU
eijMxbKq7k8ofvf58P9rYS4eo6YvjkWVBq8BPvjp2QIluZfi7Crkz/YMj3Ne+ELksThCMaGdMRsM
k5FjM+RoWTYmU7cA7goViEaBRTjBRAU1gS97BJe5ma307k6fnoLZxacGp+UrZvVVXNMjumnZSp4/
ptaqJDcR9taQsI08MwG5bJLd3rkNZVucABKBGcDLKPfGvSUPhq0NXq8tUjVGHZHWqhBRcj4I0m0c
dF/ki5nJfpASh3vUIAIwc6AiIydYSeEgemj+vBAoxU79r3WGuRfKEkXoqs1M7ARopSs2e29+zsGi
IcZW8h0AytZMOZb2aRGEByXhhnYAxJqyxSRq+DCpvrrSwJo8NxMk5SbsNQQnQSixfiBlyMDUfy0X
vIrkwyJ5uGaNz97D6X47YWpUl0J9Q1NNuonEZUr9E/DGx/P2d4EtL/7TxnKpSK4I7Ynrus843RQp
KCvAJ7BUwSYHwwX3sgsJR8pXpcbeb33l1GUf+VlEIJT/DTVOXfVhW8Pru7cgema5mu3d/HblF8TJ
F/LlXBW0QT2rMe3rYiIKbyi+3gUn8HgHUlfVFT53sFMl5UFsuMItNa0lgk/f3k1Ov2vYQGeGEe+6
fvHoeujzpR4eGhr11seoFTnQXoU/HNN0OtFP0iA3cvi1LGtp5gQhP2qRj3HjjiBKAqtPUjQq0LMe
UlvTTsl6sDMaWxtRTv9AG5QtjTKgPbNeouuhfGe7TyWmlu0pVk2O1uOmxFSNmNk/6fqxosgqmszW
EziPFxXmw6vIapGwHAi0TQfu3lkMgKv+ja4oUahRkh2pyHQhmdCG0eDqC7QYu/lrtIUUu/9b/yai
I/8a2AyBYF7ANDJ8OH6SLkl+0ljpJrNVj43g0v+IZ4sx+yG0zJ62fiazUmen3q1HUzLPRfiKnZ7q
C9ID/Y2AgrvTfZM0aolLbmvyKn8ctGjfZ6OnZwYw0G3on9nZzX5A9Np3MjUJNt9Xqt0G68GAod+a
she+717z63gdU/iohAbFN4+wYksGbb51BvTETkMLNEShXHXny6nXc9dzPc9kO1poqNTmlrzAn7Hw
lkRN1iaBvUJzZTOg/vWkLYE74U69i7aJZ898l1wDg8CIBnIV6tDRvCeQJfA1NiYOkFmSYhz+8s0m
R+PZM2kH3nkml5zkxx3r+5m/Czs2EjRDLLF7G2iRKvZpDIzOTH5iGr5EliazXtMoPu3gUSn8xBes
yOrlc1/7tS0a+8FX34+fc+U+nW0vB/cQ5Y/bT+t3+0giImZrjgtHXv3ZjN4F4jZE9D1KX7vJYVU8
apJ+RksSYLaE6UPbNB/KXuiD55B+ItvXoxQ41SUIBmjf10CBh+VbEYfFvj0P3zQkcw/4emt9AbJX
E3yd1Mndd55Nnfh3PkxORs+orGFe47jW7rqHufk/zdNjwyK5j74ToVnJ3mli+ZzgVVAQAwTV7zZH
Ipb8kTSNFjK6UVUJdv2vJiSTPjgL+T960ABi9bfJ2aq7Ub9DLkC2Ck3bvP3uOK7PPeOoz197sSD3
fFrB5FSusf4iMZQAGNH3i2Ol3qhbOtiIBPmSAWfHCgOAUVjXLGDSMCPinsKlq2fgTowio0GdKbTQ
HKck7sQNtnT6Ju3oKYvAE7VH5H9hshv9hSLzl79gT8JO7p5Nd+r5kTQ5XdJU971puYQ0rHbundLx
PIwIhoUQ9mUOREL/b3owGy1/q/s/WedG1AjKXgm1FB0nRMSiAmQaZgghzyTd58rLMl5ntVi+9Fmm
pU2pms8axprQit5vRVEuDHNhI/b5tQ3ou+OqwuXEg+mYbOPWnWSF1Gb8rmb2YfBmy43S2iJMzFSx
obA9+tn+u3zEOXfFGLFtMFzV5IXzHD2CAL32YiNylfzWJNaR/2Vmr7sBKL9bPwUsFBHbNCKYGAtN
CBfUpvnMZn52cH4fxbWBSyyufc5qRi7zBaSvzm3Kucrd3KSoa3oF+yVRhOG6tI3crtsx9DbPnxvy
xxpdsHeVnsgld3mhz+mO8aQL473iv5158b+YBbx3QiT7Yg7MQGFDjIYCqeGVem1N9EaI/Jkp7hjf
6CRxQhIkPzCP/yk7fSk45wp2Oys2K5Km4DsUKzenBySfzMDHTBgF4+4ceR02ueV4s8gZoGO9SNOg
B/CdQlg26EtfHaaFqdIwUhRhkxAdpKnMJIAb6N4hJX2wseoxkgTdUNNyhYzDzGah6opnPfq9S2H7
X4G0z4V/TpFVHTBHUkon2Krt0bLLf00x3WLa/7XLd1WCPYFy3Mxq1iHCsadJY9+Pw32rpw1duZmw
kjI4nqe2QlEKfteKqx3j3RzoFciDPo8lllC05AsgilyIy0Mq+zi6vMA/CzfzruCWO+8cNT+WnO3w
nq9l5202Cp59qCFkVOyu/v45pkNv5rvaQrlgWIP/QU+d2BjdnB+e3bFqk8MGhX/NCR66Uu3bCl6N
BnEs8nmZGA6PiNFEWV+Ve1VWK54fbpvMQbmsLN3LOfHOwkCwd18rab1N0deDGTQGuYxb+QGlB6qk
Y5a6s46dchgCmuogSGfgXMVOz4RmW29UqfuwzQNacPR0ZvpnA0YYdQER2JqttjYEfpVY5ix4ib0v
EdKxXzvAJkcrYJTHp4T6ByHRERE6mZdclXldzx7RToXpKtQRd7fLGuhH0dFc/vnAmZlo1W3v+t6s
1cLVbdoljOuu8PAwOAHe/kSVcaMv3TTMoFybY+Zlp9C9XE4QkVvYsFG7LLBQzGz9Y2HpyPzsjK6N
VvVCAzOYMtGjXYWyjvZXXGvbRzD7vaoABx7Mja9xVrLn/szGx3R9Hn7ArnnEd1u00RvTfOiPkIHv
o0DbBcJrugfm0qjg3rqePeKBXZ0+SLVJoU2eHuXfreIBoQHJ3OkPcdCilIoFyLGfjN0jA2K4XAFY
qSyisNHI43y58OaFd1MLZawtI/1KT2s1UKrmhRuxLn1fZOyIWhojFZTleUO5gFRZa2up2Uh3g13c
sdg6jw19p0C9L8aw9SFsg8K3jPnivursUY0F1DAnI8R2LxCi/q0o+N1Jo2z+c03Ma/tu0s2pSyDu
KWAXrGkMfD69DVdiV7VTvmFBUqYP7oXdyCAEZs1f8LPw0+3aM4r3Z0HiAwMqUNOUd2t91Vy5wmYS
VguAJ2lxqtyD+f/LYZNr+tlMPOYPLLsKXDo47zjVlDFklQUMJrXR1TLHvtU79e8U6+SapmGARauo
20Irddu+3XIRCYrTaUbm+JjwjypuyUY3Dsrwe4TKpux0qLWsgR3WdB7DSIiTrZ2rsNzBmu7bfE5e
pPWgih4f5YPCu/ePkfXD+pUZTz2JiGCyI3U9082ocwvQRRqFbER2bOp7ZkNC2PxuxMMTbnQSJijA
uCj75PkIe/YcaEPa56zV183/kMTcEy9OqWW/DcVXPW2A95FvMM/T3gYZj/jITbNOHoQUz6HSO2s8
AhCxYbzJFfP3UELzdY2YoY7PG9EdF7l3yA7xytpfd48JWi8tl4Erpr6F08A4i9P8I1ux4eCli0xf
K6JFgJUxPZdcstHNFUpyN9Of/oaPDjP+NApoLMRmE8so77OnMYfGxd1bWps53QRJP4euE2DVdjwJ
EV47XwX+KzVxixHc7rq1eAJ23+1NqnS/LOn+45RxJyd+T8yy05YU5suJ7LLnYiHVUiiWGkRtUIy3
hfbK7Adu47OTfqNwr+S6mfWQvOKOottV/tEvhA56irgaJVLct3UI9sq5zX9nr9yiKOeggxADX1X2
saSmmnrYn3gbUEg59kC3B7ETqodaRR+A2SElZx78H4avwMLcu+BSSZwhHUioCQwVBr+Iq2wJ6G+n
TZNxjh/m2y6hs+yLaqZT128IonFirtxCxGR4LBTUzC/qZ2o2L1oBNZO1wWmds1iqp3xuUJ/alDOF
rOLRoB1PL82EH4+IyYVCWS9wH2ttJlb/fGOHE9dd7EALyOmeEI4/f1Ns9MZhnpwL9wuc1NJ1wfZN
SrTjmF/CxGx3PwTPr/2O+RI7m7MqlwdfKJXWBzQbkfQHMBKLhWOI73zUBAXv/6bh9Bdctm2vGnOK
zf1PEC/OHPCSA7eWyXv/Nhh5UP8N8ACN+3VJ+Yn0GceBNuhHEO+AR4NbB71CB9fW5cl5OZzCi57A
BIIgRCbl9e7W+TyBNpGH2TYEPe18qYszgyVEJ4vG0FfRw+ABT3vGTLLbbf8iUDHJJmV2W14peu0n
btWmRshDcLnI0/+VNWFt6f0xVFmLFO+o8UVXsjQqguVExFAXKDDMOKjW+fjTR8TSZDpdArYSo6MN
xL4ZOr0QmfGZG6Ro/jFZIA6pGPZkf39XA30rNO4JUO2n9AL/h44f9YgpxutZ2erglFf6SMeHJLD2
TpzzbtcXqH81fnrVI1vSiyjF5Pqy1e9ZwKPJXcjh9pCvvfIqfFkQrn/LuwwNxbWArX6vFLO4YrLT
O9hkmNWB2NuVDPPOYE+1SJPT0OriC5s+0ePG9pLA9z5snjvyKVOCixgp5krYYyvgbDyDSaNSAcT6
13fJ4lnHxYmhS2yleAEkM8334fimyWTXS2nr10D9llOGmNr0SdB+smMJ7WNUDI3lcH95Ior076Mn
RpuPxT/0G10OtFU8O2JwoZUmLBTEt6mu08S9nKgEnz1gpbGhDbq/HOSHNd9wGEgY9Y/ixrz25Ok+
lMlnyLIK1ju8b+owCPB4GL5c65b79uJbsx8mkaKEc8JYwscK4HrMjlnKhrKu2w/ARFmgYG45LAdb
F2+xIMt5IvKBz2o4u0BckmNR12hNAhJ40l9Q26x7JYpD2R9IHmptOSeuQRIqSCBPlNEk4JZ82gvv
48D6F1JunzaOQkircnHKdMCIeUTZKNPNYU31YDA66Ht9Y5AQ3HVhpyOBCzWZJbnyTlppojpV0yRH
BNeYLrwxcc2M+h8kZo1fIlpMmiCKQjlsFjFpS5vH1qYxmz724RFiNBb0ijoC8UXdy2iPZzFTvipA
EWc6deSHynKOjrAvz7S5Ao7ZBehsgBlHkZoRiHm+a+SC2PmUjMcWQWhdsdYboNybNo3cdGBqiYk2
yfk0HECkiDDWbxGRQ68z3k8/2n6/OohuDrWHAw1pmZM1cEqXgNV7otHLxiuObDHDNxCO0MKBDHBf
+x0aFcFdXoQYD8I6W9snZaVWP4bhuG99FPVcOmOu2b61ZaKKiBqsgtzJH9r+grnl65KlToWt0yi5
Hr/l7PS2cuZbkRQz26m8aVQDUSn0pttEIZsp62gP++cr20RN3T9R4evp9jncc4QpD0X7wpHOWKHd
waY80zrL/ht2K1mw9yKJE6ZNmMsTh9P+KJmF+U6Ol87GrcO5SQnIm6E/cQ8mQBSEuylaZIv+V00Q
j2GaVOpFHXyIE7iEHC1S8zZm6m8v5+e1qH3kROUa3eX0S8BDgtAMYj+2cuUUSxEHaxyaLTEyjABt
zoEPWfPwKE6gRa0yWeqqNan+26qFB3aiFeMQU/eUZnBVVF9JnVXSdY3a2gjz9AF5BPzr7dRKr16N
9iOGwqA78IBg3MmwL+mjE9I/BuVoUGEECT6nFftFPNffKPNFzBzfvL7S+8HIBYfDFFEAmvvzYz4p
e/bva44MSp/c387HYOlG6goTXrGefaoVX12/kmYNO7Pd8yS1FNQznUrryr5wrIr4S1U9c9V16AKO
ECOLtaO80cTbQXoGZuKwu7zMyDZ7c+nqQNHT+x1G7weDU5+LIYI3LNSsP8gayOcM/mPLDsYedv3K
/2cAOuHQD1v3dQzH51Z7IfiAXm1A1DD+MFUZwXIictPLT5kS6gPgMhESr2g7t/oCKY0G5VVNUnVP
9KG7sff9kHtV0DAPVl9fu34S08F9hLJVqajsLAL91AzBjqP3YFoEjHNmXnmaH8cRzZJ1rmgK7I2i
IM3/D+h/fZBLnmjc3C9fmygD2XV4lww6cfiklW1dHQcS9j215wDys6qa1u0jZnmmbuZuxUqe6xT4
Gyx/l5rOWAYQ5WzuKGxMn25Sm4aMrZf2/rmN39zfjILLzcxUrfowYy6lm3IVdLsrxx3ClpTGrlGU
Q/OwKrIedhjbtN6TfiaK1xYzKqEvTdRYXEjeVD98hlWwPIgo9DY+wK8y05xiZA3f4j9KSDW60Urp
JMuy1Ko+avsqiSsZZ37DC2yPqJ0BxJheVHr19B+PZ0q8l+gCB5YP8gdz3bZGsAG+TOOHPn3IaTBn
BBHAwpzXMwT09F4d88DlJWH74O0vIgo2zvzgCqB0/EVvqlsPp8/ZMha4iGwIjXTOsB8K5kSslVWC
Mkvu61XzXrks5qkAsVwcYXBtICATA79qNXQ5eRpJmeQlN0m3YQ2bD8pjYIkCAKHV5vW1eT+trz+g
lEJlbgc2IPYtqYJQ58GLJT/nL0PsWS7+7Ldob5Z//+RbDFKGxMCkROixkdG7/EnqAfXs2fI1J6bL
SNxtuEeOt77gIpyGU4uDxFLleT9TdGj6ae15NcDQ2zrkcsOIlEgXeZKX6Tva2dUxC3KxkFd3eZpl
DGWdHaowfuSebugC6Ise3xKEBj/egRAOjO4moGBxLCm+cUTSTCgFVzdwH14+0nWCpGRaur854Mf2
I/aNUNI9EP7VfVQVpovvIt2V3j8XVqeEKizsFi53aT9YUwA7DKy0yq+EGBoFxYRWHgK+NdyHjVwg
3FDKVRpOEhBjeVXUrwGUAOfbeQw8L70ikzLFJdp13emZY+YPneCfiVovnG0tbTUvslFYCO5gp6CD
fk3NkD+ScFC199fG3jcBVWHGCJRv4uLMLNj+ZnZXVRbvAVMqgD6/UzuSvQZLZt/y/Z2j9KcTuSs/
RZWornV4srkIfLAkHX+kjz8IKe9IuWGfpYGqb2hkSiY2bho64d4SXdtHJtrMFv7Jt/5pKL5SweDM
ZKT5yMz722ntGN/bQ3SW6XQHohRHCX60szZkR1wZFBQgHs5dHcxW/KQa94cQ1vTuakiHxlZu7YKF
5wBmGfecXP3rZlzdOGnYphZenl5IFe9BlnLycNbmPdaL2RUU0oEUKQHv8BjG/5hfFOkKgA7nsyrf
uCnQj9nglDku0YMRxNgWmo4yEbagoNHF3HRi8Bm6pQCwMxmPUcM9uoteNYgRWZMwfRbRXUOYtbJQ
1OTfQkSO99jCUvFEqM24usW+vcZeo56N+DAieCDKKmqKKMrq7ef+1OlyPreqDTXAd0aonOVEYvLn
YCoG2rM8boj4b5hUiOSI9FdWflW+mOIJ0zpWd98YRk8oMzWOyyCE/wsfOB9yNRW2GHdjuVwhh+pv
5tEXD5mGST5de3AWx7aFVXARelXhuiJHwlaGUa/Pguom0ewL+INybTBa0kzOqQ6iY+uJTRydnnHM
vf/jHGyL6rpKKV5+JZesx9rqNIbCjz99wboG8Ck7eztSsbC1Xpg/tQqdSv+u3Tpo0Kvxy0fPCfk1
fRH8Mlix9ZHmAcDpNCGuYcdLRtFI1uMw//pX0Ww01hqPSTsS8yxvcZEcFineDZ5ox8Cr+onk8l23
MLtLsT/NlW1WXuL4g1g4E1IWMzgxB2x9KKvvurky2O9++pGfpjai9r3BXY6v5lC4qq5/uqFaobdd
EU+Udy8x5DfiRAi6A2YJJcFz1SNcwDvh4niOlD+tPmuJzwU48PniZipM+PAhL7+fXTpXJFJjxA5F
VT66nH/hSWVsxvx85+EMyEvZil9F3D2F7CxdevO0RSWUaZxHLIvE1P6rw562GKpIlJ+7n3T6+cmc
mXKmgPWgH2JI3tQivStT9aGZOXzjBIuOqLGFlzChTXtW4cUxAZeTiPhd+THXH8z7wuDsFMzRWDZE
cz7+OmpMgTsIsGTEstTlOVzOsNkkZRbDU3Tz/YCro3KzBTU0gWc6o15Fx3apDAvEbSyFoOig0ooW
RxGtED3UBQd2O2y5C723r16ewABPwjrWQ/YIzg/Ay7U/k2uSoh58+S1oOGv0sM8UeJFJM3TULXHl
beaoUT+1QjQlIKf4sdoVwffHs9VR9c6XoO/XEbptVxzdBrCbk1mjiJJ1XMv2eIdgcxewLxI88Hxu
sOTi0/vIyPw+MHK5ET+Gm2i95IpRZjM3kaovgOC1lcUbqNl8EcafZhQzpLxp7KqJbzq1pceADZy4
3rn8ua35EB2AOFxCPMbAxDNgqj2L4ahdEGIRp4pFNQ1IYDz4LaGHH2HVch9m7DmqBbvU66XEM6Do
Pq93oFtzITd7hvXuzzNbgil5y6/05GsSwwQg0SuypfKeI7LdY/AQmPv0x7FXkhlPg6Z6GAH4MTvl
+eoUriCooymqJZv5GcjSIMLHk4S6xV2i6QyztG8LZoZeSnRMHcV49R7wonH85lVLHYJ9PXSRABzF
M2V0fGbMjzBhOJHsE2glFPHWyrdT5eQA08+6UMP/nK3tPIXSfT1z8U25p7tBhz5riUmc2wnOACl4
lk78+aK86yg++Zw++lNh3TYDyp2gfZVIzFsYqK1QvAtdsuWQCcZJ1FEmjoq1ZD90mmblhOT/CkIp
ycjEgyjh0UWp9Zq9KiCufrryY0mDOjZhOLQKLQh3u6R2lNeGmHwcDqPeTRyChWqUPHLDeXEWAr4t
ke/69yd3JpTWg29DtMLK58A6Ek1ubS+s4BI5FKNCcTQnTLgBuG7eHJPOZHcn14VRL9V8axG39AFY
rwg/WKf1FpA1qZ7Nu/YPm7x2uN/x+i5I0kVkixueCWLbXvoD48jTWkvutqwofZDKhqRdlaD9oJQ/
ChFLhfVOrg57f0pn3dhZ1FsqNXF5mruKMH7KreUZYqOeY+v/sJgAkSNCNyfCM6JTAJCWZFGiScYu
YGjXi62eo6+Hhtvbp51yY5xoJOn1YKMczCbT34BDTmiQp3DqGJWBaxlktp+WwwtCTyMr6Y3AaASw
D3wEXn4QyXj7iXRAHImuMqRTbuBYQikKlRSkVNqZgznno286R/XA2LvcaLMwB/AziO/ikX2vdUCD
Xa+Yz/XPkVgEkvF7NfWb6YE2s0KcAQ6pD99RwuSeadM3LUrZ4048rAx0uOx6J2XvLuQ03HX86Qhr
BfhSDBZ6jYZdVKujSlWjdnGkWq2b/qzDdivOOSM3qaIr8Au2NBiweFV14RzQCG1s5PNm+9h3IOQU
2qVuEilM9G8J92ei8YS/MzFP3reBvKTg21vRnqft9SgcjjTpO1VXaFXFDpc3anz7LdsAuXFjZTOa
lmk3AX67WAskEQpH8JAhy5DAFcko47CHFmXjdiRi+GxDxssNDrT14c1eFlzHz15HnGM0hZEimhaQ
0PbKydVtDT9GfOtNdyNrzgNnTv/IosaaEF7gQGdKiFFvNa9x/Vy1Sfz81sfikuOH7Y4h65nf4Vic
d1TRF1WVW5KMVTtcgUt+Om7Q11Vn++79rErps7QARidSYmwyOPUuIp7T2xuAuED7Jg0eNCkWt1Q/
hdwQGBrmBhuiXG1z9rDGpEQwhZCvj41ZtwzoHzUnP0tWgnduCTBkqnqRVBHMSinDuraA969UIZ40
ghkrNEHFhj5oEAAyt1clsCGm2gp4sPnV+6CjNw9HtqkQehEYBR6lmleqtLMz5RFfDLFqG6Oy6OUn
kRmS7Y8UKdFBn/6YDq1sutB/i0BdnCaZh+F+OvvvPphpbnP2+1lodauduxZZABhY1LKrCGEgVyFC
o9AEM4VAg5mv5MMhi1g/c4pdvrAFkWXn8GmDEFg2PKaUTp82ahyw1Ka4tOfuTZFbp3ZrE8kyN5OC
cxIib8l8XKVGM4h7J/QzF7hwSKlym6Chan9gsIPo8CnRmCvPr5sA6QDJVKsUcx6dy01CJP4L9o15
fPHX0K7mXgdPXhtBhoKyXSXTw31bvlHpcIE1iXoQPr7naOETtr1pGJkd4HOcmpApmaYcmvLMvZ98
tf6/5e1uvrkEjudQAX7PKO6S5JS4aaN9v55iDCDHN4Qhdimc/gBfRvMOKgnj4i4zSe04j5kxLZ7T
et09XKHS1wGO5vCc/n8I0w4lyvnqYvL0DRRjaimGIYPpEO1WoZsv4Jbt4Y7KAqJ2vcdX0m7GBvBQ
OZSgIMrZuYZQft5AIJYCKO05n4hWDqiFMPtF33d3Ce0NsS+CWLVd0X5GWctPT273+GzsWTLm4lUE
tD5xQvzneKLON3BATOkytIQqbAkK855TJv6ZMPl+kWjz+WZUiWkP4zJKwlRZssYRj4eBOb00o7Wl
6q3yaR2FjtN2ItZvPD3Zmcym5j7TLmSmt9iwxUs4LVWcxdyLjiR+GwQGrj8IPR61DPXQFf7h/mMm
+2YfE4Ng69HnfSzBhvM4J70xBgudar0s4t7DXKhFF8BtzoqLpA/FQl97nNc9vBIaiI10K9bpeyP+
wVlegbSGCRfo58tLb0REPL20niU+5fUIeV5AHCGw33YOuy4L1gcoJ8HTNIrb89Cc8uaY9lPb6tmk
8qzdOxUVYZsMGJBujZdpJ1Y/Pn2kGTfmdPZCpM/P2rsnAVDtlxEirEojg6jARKUFiJhXEe5wBzYD
hFetH07tq6JoeWyP3tTFmhSXaFXQBDjsGhwtn3xvPq2Z7sI2p9oqr6QoB/W3tOzhWjbpRdqBnU6Y
zlXd5yI5UIg38UUKjlqVmAYZEW/NLlNlqJ7i7l1fWHeYGPaReRJxaRf9nO1d9V9QDzIpDBCXdRrn
pS2HyLmSfQz/VXaNEk6hBEXCsqliZ1FtZm17H4lfJY2d/SarBchFaEdXfEIgq4RCWpEI4ITTdi+9
HbJYi04iH6aIGyK68rJpxBC/tlCDLY5leFoBdU/prx1hpHC89sS0JpV4moE88MBD/HC/T9ddqyPC
iTOcAAbJcAFOZyH6Ymle5+FNqQhHw1brvVDK6KayhV1sSZE121GupTNZtjkWD8//rMxKac5n4tVv
DGs5ojFqB+DZUe2etIZe6NH/FNzVqkuuqs6oSNlpD2WZVwI66lvYRhpHfFR7t63TldC/0UJkdYCf
cefhFpNRTnfkOuG8PafTrOBQ15fJtcyeAdKQrqYPa5e03+jcZV1SoOM+AGyh55NhqUCDyv9uNswR
BCpKVStK4htex3RtBceJ7dxrf1b9eKFbiyTHZ4OEclCpCVhMQQp1Q8EBZGND/7Sku6frbPOO5Keq
adJFj6ZXP4uL317Ic9f/u0Ivi0dpZBqSVaB8Sm9jK/IHEflYH3NFKnG+WmfVtt2DRHuU8WcEL2OJ
J6VOTDUoEZ6ppIkI6bGLhWw5Q97MHFqnQroXe/dXv7CNPVZeKNOcfp6LuS7h6ogAFFUoaO9yMV4H
ulp56snyTw+AxPF9LwGTuX5IpvlqI+8hewu+l6LQVnV4QwFL9nqUynEEN2UlGZ6VGxGaLHPPFH69
ZhRg4H0zFivre5FzgKXLvZWMsLBn+54u+lsqIW1kKzpqolkYwipH0WuJQWlEjfET/3EORcMcyfsx
e2FA/VzJhyHRc4aDns0HeU6rVWImeo/MXBGvvqcU1JleC9uzFp3y4Ds8Gx58x1E+p7r2E85TtYCX
i0H2XsM8HXW2uWoh/oOiPpBRvZ/wk1I3ZtLX5dpUtoq7hnGBCWrBcYl5wzeSg+tDhBqxoSW5UKEn
A5ksGw+xdo7L2n66vKlfCLBW9djkefJo8qI29SBDJZ2XXrbASqjKi0cu+puGnLyvX2/xQ7zXIVjj
CMCfFK9/dCMDcrpZUTs0kXMQR8EG5ycniAg6fqGDKOkVyFcVZmuR9SU8H1uqpywHy4x6chpF27Lt
TXWfMuYzTYPnQVTnkbqjZdOiKihkZ8z/6RMM36/0gOOpuF5TlQOlxrMTglrXI3AiQtsJbslrVzLG
o+O+bTdRngSOE26DbBqUEEGDgMPFKc6ZihMrOu37GR8NOStmovxd8blBN1xzRXiwX0BXh4KdH3kx
mh38vLyxEp2kqoj2z4v8boShu991f82CJwSvEvKqSj8LtO8zalQWljWhM0cTz5dp+JfjNJf7rG9D
IhNlWRA0628JabWZjHyvsaGCt11+Wzp3jY5a9X+gq1SAQQhDx+oiSwwAo7hLkAAbiIM6SqI1Aa/i
JCe8aIMYJg/e9UenRL49J4EQktKp4/VhwQtgA7uuvlZTNcLOCZghAeHsPekdDzQSFnPEmCUphloW
TdnN0coaaaw6FTsQOb+P69Y0uSv2JvAaIr/bgpz0GIL+JaDEnvxdqdgW5tlMWJE0eCLxPwxJwyyA
cIVvHYUdZk1XLVv7N5vUKiLtILQim9m/ZR7dw7AORPaepaYY1T4zaqhk3O4BpJ0aAXSgpgbADBCL
s3dpmYVfUYb/S2gVeW2WkFII4QaIw60Nmn0vMPa+BGFZyTvgi7QLPk6vN6C8e+FYBRxwQsW+5DKE
3FylLpmCedJ2PHWXaoUI7ivgOzWh6QYBczpEbGKwH99yieFsS7+7Z+QVPupGq0QsMHXd+JaJ0+SH
035ducnD3Ectg0ANflScTOE7eQf3cO5QwaXS3J4lq2pUWBuFG06bzWEWJdSh/PFXFuuqSdP0Dvku
RvPTLsx/ZgJ7d0OFwyvxaL0jplKYdGC4Csd76k7pV172qYu+R75O5y5527wVeU//j4zsv7/Lo9oO
P3hOzXLT27AixudA60yJLuNwETAyPm0s8KY9bU0NY2K8ucvXeGY2umm7ZKF7I+Z3jtK7H7p7maFe
M6eci9bOO2Mev7qmaZRwgOvDFG4Si+FVO2+qQrp1EZd/2gJS+SXrloxJEHGPx1tGvPnFkIsBjsj1
KIWbRJAHAOFkYJZi06PA/KoOoX8lC7COr7ZSfUwYmED7QpsjaYPGITUMzQoPmyG9vQAjXirbYJ7a
dMwY60ZUwCl7Wh+Oo0qLMDspkdXiXOA2KpWtLvgN/FKfY0LgFU94a+PYK8JGENhOretCYqk/6kmY
JgMspAWS1RNl5VgEVPqLo5RPu69HC29b4n/n8HOcUzzJGOqJBoK+/mnDaLq4Ci7abn+hnG2sVYWV
nqZVMa6zl4+4N6gAb6chWAVYsjqPU5vUJBnC0rLiWmlasLh/Tdn9fGUPo7/hMOspev3pKptLa9op
O8p+/qu+vg5CfdLuhP2y2u42qhyzSMp3pfz352rdBiBDQhAas+9GZJ4iS7Bqt2d4mAe0CymwSk+8
bTWigm4DaNx4iydjcSfcRYkQvN4oB55iK29LGtUpZoUPmr0cZDpzlpMUL9SumVTwK4mwkuxZtPbC
eA2fvnFQw0hCAQuaJmG/dRDCeZG/h2IAhE7CK1ouUF2Ng1mg56U5oJL8KzAL8pubLw/oCeNb2Y6U
FkqVdj8yqfYwvOufWqj97Px30coeJ1qN4jSoEoSLNwTVASvVs0ACTrAvBH2DRjluRzAPn5y+v1hD
jLgZzaqEXkYSPHJeizEEbyFSL+Rdcbsg7FzjLQbqDVSfS1OCSkxIjWOpAVAuUIqHdG/KXTP1v0JO
icPQO632O3f3AyVsKczYnBkPwnfQSjm2Obk2siGOiT8XAsHXIAs4cdhKmhMCtUpYgq205ymyc8Ne
5zUOPWmtuz/4MNmlALYG8qglnSCQelTTpmFOBuBzqFGnwN8j9038ESpEmlcBq8CvTQWGBsAwDg8i
lgSFOWnlR1fhYv5uFegFBnlAADcnmTH/LnZopX6g5LTT+JQh2hEpBzGH10iy3xKMBmTrmrsABD+a
+0BAyZTjaRLkydG6VgzCCk1QzoLL2BULWblpRjMNtC1EYnhQkluwQ9MjMR1gD2zfJx1vdvqVPZjr
uz6TVrfLGzNn4/4ZtKnzFJCvZ1XAqjPaVv+xhIKXuvYberuRHRL72KldP2pZ/l+SV18pPb/ELJ11
MJmzPVGQ+jZCXSMsl5ytqMBCbEE5963w48WFi9jdYTFuCmsbgWHmstN7apeEUQEbjka80Z5zKY0J
f8lJ3fk7hIRkJLRdevKL2LaKCOQBHfaRSmP9JC5EcOTo4TPX9fB00QefvZgutYHYeqPzsdXbeNsG
hCdRwsmJioMSfSPaupHXmk1yOyS4uHz9Fsl96FpsRBXFzH5ADzP7cex9pM3JuBuHxYzqF2X8BaJ7
NTqHqKMh7q2EevSh+zlX1FeQ3OGuV7agYhG5z8oaTEIhrNcb0fOP0Zx99t0+RMl19SBPf7Gysr84
itRD1bPT5/5/063KnJUV7JPO7/ADgTOfXZKN1LY14jwTspCjRhyuBtdaqEv+KEEnVywu3zAqXZ4Y
yeY/RXZIrqRkGjOLaN2c+zMJJ1IRvOF38nGQgygxNZHr1CCWiX9aYO6zKwPPwJ2gLIdn5CA3X0gI
IOYoIDjooLDJU1k0QVnUgSOhtsyt+N5H4+GPCAa3tVm+kyWpk6OWwR+Q/rLM4ixMgjuILfB++hqJ
u2fAs1uUd5Aeiz+ECveN/zwhMBosGHOU/3UD5leW3o4DYqlnXlfqQWZcE2yCfAj//rx0H6Tq/zX3
LTuS+xGYRxA5pFL+09Ej26mNS/heXjw5k4TfPOBHvgkwsRSHa01Im4XFQQZ1KY5qN1Svtprwfrrv
t+bwXNuHoMCon89KnSaUbf/dM4F4RekQLoJMdlWxOoJnrfbXcjlCdxqs4jiW8wdaJFju6gYKpYxh
Rho5sJnlH5Lh5Se/Ro8JqM/4vyGanHKK3Fvm1AKcSY7Il2kl5GlynwFGF4VOqQammipUUvFEYOvn
2VHfcm+N4oHKJrfs8l0Mp/BTUHdNqEpeuIAGa0wWWR5biGqshj7DvMgEXkXxc9z4agA/1NuU20yw
/JqMx8PCk+ydCUGqrHRFjlLeOPNKwoUYDTSWP33d7L/Y4Kt54Xja3swlFHJ/7f2p+kx/7AAVBm0F
fiYDkDLgDKl5jB+WxITWF+NdQuxHHAZ3C4i4HbEAvFkdIj58uU7SnZ43W2Buze5hKRMU4wQYFsfU
+WUdwZ4xkAhHQ9fDOMSkMG2uCHIUDdbH2YgAUX7Dnnxi3yWb32JwL62d4DXtj6T1l1MC9OQETrw8
FTvxqSy6bUrEQwEZEAHs2Xg1ZcQSS/619Erg3B22FRJzM2ikj63qS5nkNtaSgg/OwqhdXPzAdekz
zb9tC6yF9QNSfeDAfMbaguafgHymkrOLSGVwDn/mMxsAZUmQGi7w8JYj/9SKYgaYOH5CsqLNmINv
wNk1lUTCFeDp/30XwmIOJjB4dn1pTVqMxv6wTMFQ3g3LU0GKRUKrR0Z9v8hQeTXaz9w4uN454Y9d
NBS84ljCuIohgd+uzTz07Ks63CB6F75KDIJaKKZnNRBYgjI3AEajr4kThZUTqGkgAHSiTs7uFMrQ
c4Qzqp5tuF5RBnDAo4Zi/z+rsKDkf7Umw+6k1AJ/aCGJv/M/ix3hljdn6PrgalBmwXvVB6rsmcZ2
yJr6hkJuM6vle/pzX1s8Ej08BJwjLfjz2Nr9RjNVU0kzERPWsNfbn3qDWUP6NgIQKX3JGo5mQmPV
olwMw7Bz+4Z2BR9f3TEgIHq1sxTsxevo3grhumKC3eJUUxspL3FoRVjDZXlPwXYSrtnzutWKmNL5
CtAe9WJ1AFz+2ofRoXY/Ox52fFhc30iKL1PZbvNsRvj0xWB8WPurBdxp4bp0V8RgJyYvV4cHM/+N
u+JpRsimDCb3WHNyPgEC9yXg94wm6CidIyVpKvzkVGCMPe04Bg3+xUCIZAx5hDc2rA4pxqXh609M
JD2AtrT21akx50AlWSaf0Ia5iHGSibclsY+1YUYjxKFkNHw3mHUIhzmcgqGIXIsJejRwD7Na0bwM
WP461Z+q6VOu+35by805A+RFQ/+FKscTP7IX4awVK7mijAp5TDjplOarSrIQgsyGk2NJdQPiTg+i
AVsWSbbDizuMuGMjz2L2mmVCTtJOntPvHXEKJY/sL+rPEvtbgU0d3YV/O2JNsfq2XR1IjnxO59dx
8EzwEuy7RRIhFelIwhtDHngL4YcukiSBXnjTl54HDH+Qj9nWg3bBmDrmQwRLGeagrvp+oyDCzn8z
VE2dfy8UmaHRFzBVpw2Z0UsK39YrALdRRqrEpSm1WTPWpv9R+oBubB29sV527yr+qM+jKBxEFUX2
8ok+B4kc37V5UiffaS7NGOVxTGWlDSV5kpqNUj5Yc2UmkaVsRZhDIKAJJ/sLD26otrJ3S7g9+98e
HLWFAJsfj6PuaogTqshxynuUV+n+Ueaih8/YKq+aq09fTeqwStxU5JVNzeaZLQlC3El/3ravWbJ/
8GaBStIx2g8g4kfAxFj+FluWFoPtuqLcni7nBeIhviFujXZm5FgVIK3e+35rsD2IhdmUwmTrsTCT
beeAin6HTJ8HzJCiMWocchBPknYVLR6mOLCgZgjLhkJA8zwmswStZPJ1yEAIw8XrOqXkTjLf00tL
g7SQC2u0CSx3GPq6SjtzvkRWXW61tzBgLp+JtaSQPWYuO+dKYQxe9ZdHCKBUE1hdvbEPr3INa1DS
rxgDm6xk+yGCYhBU3rjR1IMoNmXt96/U8Lm453j/u1eKzE3Sf7WzPonxF1AYJO6/kADM+kQfa2dc
lm8ebtM01HfuCI/p4aKMOLojDhud20RZ6g8i+pU71TnIU2P6hBn3XS2ldGpnp4H8kvvGidg5u7hQ
nRrT8PvY3zPATxbZSliW0BkuxDavF8sL7tJlHJVXUW7UlAa50y8zjYBIZhFDk4y1aVZSgjDfcNr5
t5dc4rZAYR48YA1TSVBjorvLc3NLrbFtHE9nGtE6McO3aHma9NCIrPVffctdYPKLQWxZCmsXk3TW
7gusYOY4D5kVkJPFeHG1AMv4igDJyW9xzmxYRxVEbbc/r7IoiL43ktq0fl4bl1V4ILP2yLAjpzrp
DclnLl9+MTRP0fajEZqrvk6hl6rbXeTzfjoUyso1NmQ7/UwlXZY9krgDKUuHgWeRbk0z/YjEzxHb
/y+mRQCYW+MKQbSLbDdEg2PUz2ijDIJroac4gabaRA2T3bC075mI7lAts00+jzn79pj+1yYTYPhT
Q8agjf5MgH2UdXzFnyF4dhbR2mZtQHB+LmpqU1K7ryFmmGKGivpA58OHcUucM0yrK5T9qPCKFmGR
/HT1Z/94fqVB+vCzwxUgBWqD5LNNTo4kmC6VptRYjof85+pgWje8NSFc1j3db1phBjkT2+N98/GH
G5pAEscE02JO8JC2KvYvnsogsQjy+95/TjD0dn2/9KAymlQ5pV52Knb33pGdfNORTdKr+r0NAtjt
GEf9uyorcV8N0zZnkIu3jtu+/aw78Dzmw8ChN1TOEJ1QHK/CVQjGOeBSqroPZztZOywL5kPM0kgq
RcUMwXkluaRz+qEm6y4PAi0ccfu9/i/7m4+c1bIlbTTr+3Nf5lwKYQAfnzo1X76AqyziKNtqEg2H
C6JVvA5k4S+eovz0wmmUqOtgjzshdcSP47RVyD+Gn5O+/BVFaBKcZtxEIQf81NQEfwsLNPJwf27O
9tnqdP08U35/9ct6iM6J82M9ile1kTgE2yDnFK7lye1N409XWGWF4OeXCeswbjqPXDiIkDzvqkpX
N+mApy6/QIkLMatylreD0py+X6/tpws5okFl2sOd4z+A8pVxVbZR+UkiV0G20Rn5A1s9bC+Q6U3V
AoX31Tn5jI8MhvzpZWH+Uh8YjI5mei0CFeSMWEINAehFa8N+A4F/heUXK0ir7ywHQIuEgRGNYOrs
HKBfqtip6NZPoJvNN+vEYB8/d6651jcUmTulieBFSYmK9sSfL7gyqkEBtL9Zv+ZR7IU4sceXfqBE
ucFrmGG4GfUGf3AG1oSQ5ywGY2/6p5X6grHUzG/oi7B6f1iiNQwA2TdoznQmC4TXAsqTitE7zg0O
pRSYZSuXqlgfr88Dnx022zNIljperPg/ZoHfQqsPl+VFy4gNoBBU3sQiDR7x2GHnV2voZvqQimBH
BMgaK9URKo1bncVaTiPKAV5C2UvFGDjkCG83JOKNRoMEekW3bc9S35Sn5FeBcCHNzNyO7fkGurxv
izRYuj0E+T7IMHZL64WYv4YO6aoohkrtlS+BUXL4RmT4n3oiGY2ooEk5BYIKL6N2WmpVXfKYwie7
FqzqBviHwXY07nqYjgUrjNgizQDwpreyy7DnCYVCBlO2CUX3tw0L3hu1XudHMiC1oy/igxxtjpPt
Bsst6B84ilIoGe+bdQrLGoabIOZ9VNwfM+onqC+R3SR9BCYVQAgHDEjg5R7kjRFfIXkNWp4pC2/x
qdlByIo3dgJeL2onZpL6eqKGVjwDwOPzu+2OWn9oIKv9kkxJ+0PE8HSu/XNQmFMQprXewk5hzzHF
cUh1xw+Rzg932meqNaLo1QMiAPHHAWk3r+Kxj5jjnYfzw9Aer+HmjvD6nOG7l/eForZHXGEndLRB
rfMbVxq6FLr+wkwfTrT1WHpHhHSKHpbB2z5OO8Mqrii9hPFZrLLzUYiYH3X+yRuw4rvMZYYr5+NT
UY7KsSN9+ICC6pk3XXmKl4Zq0j0gtzBo18zSZXpxPdsWHz6RhJgYHzmMBsKuIFoetdRADcBy8khH
BMW+Uw8otsr4EHh251gFQ3oSY2Hzzgy91TSBKbWAgxQyexHe3oKAtfo0O0Q62ARJrsm2GQts1/QE
PHvcg0dTAXDL1K6MAgyV2EZJGdFL8EpydXbuqguAOZv6C8G+RWHOcFTiQw/pVu5+s17XZlYOtajb
9V6XQPExLqV6czLDIBpGntsxITY/4+XHYFvsqyXU/klayKQr9R6doTNIcehANLHG/F11TYkRISUa
uFEqropQXidpK8qXfU3DWEkTSeAPfXdZc8zFhKYjVseVe9WO04LkkVcqXGhGjQIxwFxbEKLD6mz4
h0QzMsDOFxkFI13s3IQZhY2j+2tcTP78mP9KaQ3BRXlvSbFs68o5ttWfGNg3cUC+YuZS/bjb7bQK
V+eTR5mPtcfPvIYJlPHqWeqe4/BqzX+pLqjA5PJGcjyKlvnKQcCCD2kbH5oQzZRGkkMGl1NnW1fQ
fbf4EuZx0Pcr1yLtTi54oEZjDQ74tM/hJK1Odc/gxR3k2YmVMGHe8cExwOLluzeDH+nSHTJeB7tY
wX5hMXcli92nIaeAEgZmOSAp4eGWWyZn+A9oBIl2L+n9vi52YLxROLA3dMs/3dr9ZBOj2miuMoUR
ZnSdpiT1DETsZ3VapIfiq3c+2leiLLqMECUiuocE/wPsOX4AIJLrmu8MvnXywsBA+kal65bqLWj/
c02sce9uemDeVp5vAx9qCrKK/CBewOcwGo0Q1OqFvW/DKabSZTOYErzPIOBqVJz6tdsfpcKFfaQ5
keWF+yvYQmvRikvuS4gij/0My8mqCFMR9kR9FpmbbD0gv2v7KO75jKPvwc2VoMWhO1QTlHTWM+FW
3Rs1QpUlvPIIm6i0CRRoOW9QNyMDnC0Xb1BWETJgxqaic1ooceFYKL7xUcf1qddS8AguplY8sPg0
xm/2JFws2P2anaEoAWDYSveWZM7aiYnmUoZlnnmSnll13hBMl/drlMyqyM02ApJQ+WCCS3VJIho4
sH7W14V45Q9ml+yQpQj8Xu4Tl8JFTVmQY6D96J8IxgqqHkTxBLtYTqBE7iTU9/cIqvyUk2HWfgcJ
uAztFM/C3mVIs0EJXesd5DEM917lyrmGxaTAdhD8MQ7mfWEYf6cAYwuvLgPMwcd8Uv+GLob1m+dQ
l235iuQmxzS51JNew8GiReHgA1k+aGVsteluw+b18QT4lFRRNvsSh5HCScscBFMVVnXrw0dw3SUN
1yOmezFw8Q4IjmpviSd/rk2tGexJe3O3keakzRbFwweVFLnaX2AznCjRrDWfjvKftD8pm4OKMW9l
bC59YoV5KLO6bkzX3LQ40e5GBQ71BkscMHReh1vpmIb27hPPslqt/ugTV07/9QKOVZpWBt1cKBzb
z9G4vqUd7uaUoGpNvWCLuvvXU1U/1YedN0NXmNtSJ/jl8faJXp1HwDg2JQz7Hy0POpIOvuzcohDw
/fbgwmd05NpfK3+N+w/unuTaZ62mA90srIJj24vrdrk2oYpHi2lYfjbnRfYKX2unhdz83AArgq8T
ooRrUJtdtDRyWPjUpmNqdtGCIZ8L4pMSaPtxLkz6lgdGVRcd2Gyna4apoLF4VqpfGcHd7jdPHV7D
yLevYvX1EvI2IDVmsa2wlJQx0rW8uY7fSxPhKqgyv+uuTHZGY76kH8gLTEuvgMl0iKB8AQw9LYxx
jfstnzIweYdM72rQp/DuvmpLt2R13AuTJUdTIkxZoFwgIaaZE2tITC9ECjyvltTIXpUwPcJssCV9
P3dZa3gjq3ABvuT+F6c1t1ZWadnvq210i5694iU+MxljW+INEuDmaADlAzZplS+MHeQXZw4kgtLY
m1hwkBgltaLImx8lcrCWRM3RLorG8MvBOqsQe6ujq4RHw5EC06OBdWa/+787QWzQDQBzXa98ex0q
UD1l56vAKyV2xyEx3Pe/+LG02R+PuHqN2t0hEEPbVOBwBTr4zxnwbC9r8ugbA/6AyximCWwoO2Bi
8WMkgxKLj3ce8OmJ/Y18LytuvAK7RZkgMloLrxWTYMcVjCZEwnGQvKZdmh49ttrRG6GwQH/G3rDo
uFbHaO9PVKLB8c0SjJ1Ax7mW/0F/D201AWAlrKedWd02MLwGR2P3jg+vU0uncm0lYlp/PYJ0GeVI
AbBKuy7NIhUh95h+oATShx0Ce3oAHf+eD5iFtTjfVrMqeNd/mwlRZUAyj4YUv4zvuyKdDiFP7Es0
qaNTsxhRhEOSVun8Zg74vRMKgJhXlSlnSf2gQ9MKqd1H1IiK2ckprkvBlLbGtkMt8mEqcn2vu+XV
zIpnFZWvpl1kQBu7knbOYy+Ab/EVvmamDskMn42uPJk4curnjkEwxxv9mwG05Yf0opvEdu4QM2TZ
ichCwPfnS1y/uEIJ10QtUzmcDew8K2qjyl/raZcpzFjltLNJuaJFULQstphadBv4TYxi3vSLcVTY
GzZd68iPbL/smBzfx8ekazk4nMGSE36d5mnmmKhlPwxvSx1ciWpupwiny7ixPIex/3SrpCrGFpMy
QArRMF0kiNeSLeZzNXAs7nV3PlNEcqYkB+pv45GkJqcWB30fQb2gTzouoL7H135JdjgAPpfziwDx
2o57sUcRwuOf4iY8IxX8bGcGetGdhhsd7Lh78u4j8q27WYnZtSgXY/BbXuTBvyTY97YtpSjCSOKG
tXH3n1/aYLWyfFXJov94HPn+tb/pR7TUeEQ+0C/q4IzAy/eXaqZUa4XM78z6r+h0FmcHKQy5fPfb
Sk9J4CRvEguIJf0+YEpUFUqw3zlieHIfShh2frvsOHCNbvcsResjASWl5m27/pX14LTNXgN/RACk
MSwPb/OeXEO33kaIR6zJrDTf3WY3dLn/rjAm2/deM14K8yJJM5nOvFt2u/cZSPu8PIPJJF50orjG
NdyheYRIz2veq+ich4S/MqJye1MQQA8TnCorXo61SBFNaNasJZKSdavG6GkseGndpR4/MmkfLhmL
Rqyd/4x3QksWioH/RSscC4WW9S+dApyZaZhzeAk64vM6qDY23WaEgTumDkUh0JFKTMYW0ZrJZaEh
U57IgPqICS8lIpM7jZD3yry+oVM3V9fP8TeBpzzaFCxtTQpsowPYUQnqLqztRUbzx7hxHEPmi/ho
FAP0DvmwBFuN57sIUeryVP+QR9zRfuZghK0o9voO6TrxCOdxDGka0Dn8QREqWCHZ1uiXJYpSy1sW
K+XYf6iXLKex/oEwZsBXZfUT2ssQtmavv7qcEXTLJdafpguPqpjEQ1YTmA/nRABvYksXiTJjPjqo
gN1g91nsO9rR87LNU6viKeU56bQGFQwEPhDJp4etEcEch19X5Yvx2dVswaK+mxc7N6vo3pXg4Ptx
OVgcreM38w6cs56Vx5QfCvQ3riX28MjfFHo9Y3ZWkf6BbFl/UiRvZH8eavvSAi3EWfFaXeN9lnx1
MCuybmmUHAAVu9OFXPGh3mIyNqg+Q6VXiQPXLElxFH5YTBj6JsPKRi0oefP5xH8YPiWEfLxpm7HN
FwgamD5Ye75VgCwXXtJ0qshrLwcTUMazuBtnO5HLB0/JBKagfXiifT1Wjj+PY8NUnSaHcfHIlavg
lVDjGsixfG8PaED78B66GjFL3JxtephAZtVZk8ZvYvOu1M5zYDzE64Eld5k88bcq+wndL/vJiXmi
LNEdx1bqkl2TUHZ5LV+QaQQdjjxFkOnXEB2e8iZmj9vm8Iib2zmWOXt+5iBD59/52hZmPXisNOru
PoSsg5lZYc7uNYDhEqPYsbCUezHe5KOJzU5q4DEgfSOFVGUXTX6jEeUD1K4AQ3m1TBN5+IJViIWQ
FDOs6DIThVVJCyB2FrjRnvpblkAf+fXsOQOBmmkBZ8IG0a1f9s+wkp4kRg+EK0vK40qureW88roW
INFw0Ou/769GWHIhPTFF8WdtAeTxb9R8P/PU+nymI3yo+rUXI4zSdv6dY2//wmyyUQ2tJ8Tc8Ip+
AjB9tD9wnxQyNTz6H647K3b3ocg5tzkuNSK/+SIyt9RteZMUNkOb1PZNlo+tWy5GYbWVX4NLsEjt
qC6FpldhIBsrvrYrES4C1WZV51Lq6QCeVw4lJpb6JD/yOY4EURDJHFr/WInyIOveYUNHRi6fDNv+
jCZFzLaScpRL4QULprnXWpJb9LY71U8QL2yoSN3p4fbI3NVlGDP/+fpryYCmeJCUFVpcBmw/78ie
/Dp7zhJRKC1RrfBZUuWsmySLbOwT7j36uMZjXLFkKe1HLGzb8/Yeg66isYkHAvauJbMKE8+W0ejF
yCvoK/EqZ5R3or6uI2wGyY8Q5LV22qdBuslKc3YAFJEXJZ0iAA8wNo/z89g8cJivY0CEri3jI0iZ
lS/I2Zth302KOiV8ZnHjoe/Zs7jYHIBA9ss2xRWnACNDTOZf4llBS5L0oGpbKTx9vNds8kRWrBJi
2rjf4zhearegZAt8vZokHENJvVt3D8WkiXvl4DeQM6R5avB3WrXRGYxZwBASAaPABHbadrQTX5/u
eSm88Zfc44EhurrK5fpbLTBVtpY5aj2Do2NmW6k8gGyi6tTU4zqomR5HiaWtZooF1fUEWx7aHhxR
NtWheBPElBRUxAiC/T1aRihmQrbzjG+LMUINTj6m/PN+nXQ0WlUwpyERxywcqABk4ejUKb/3vMdQ
zHs18p63s7WZlAQx/WPJazYnIIcUhhjhmChGpkUq7nuu1GvKf4w/Kuft2b8PE5x4CvnhkXr1V9mH
HHwaDrSpwy+/aafLwRVo3eGc/SwTXsmbzUQ3rtPIk3nazbwrgDBEFGrPYnA58ARz30FpDzkU3P//
Y5A65K8tfmrNHjA9m1uM4pv+PipsUeDJRLQoh5rWBxpdwh8gh43Z1t+nlK6A6kFE8k8bV3ZoEUH9
haRbbRwRRh6j0StNpiJXxVqjO0D7/KzTsnR53oP4Q9pMGg+WCeSgXg1Dzi9uaGhaZq61jzqie+wY
UHFQ5bU/jDL9xbRrEwf19neRWmjUsJotpMfWt4YglPK6ws/wu4E6uw+RLJ1Sa34ajX7G5FYwrTN5
CB1e9YanwvlHBz27f4+RHBtVBLbVZCOTfj2ZzV2mdcPqvM916qXd5aowT1l3x7YvvshnMU26+13J
CGjFS0Oml9f3fu6F+2hqv6H7g7wuifhYmd3t0FKaYJzNkqAwcobluVGYyGkjkN3g6MwuhfZOx+9o
26Zj5TSxzwXHqxoc9yxeVXi+VbdvsKGZz28xCF4AkCfpA73/GnFJq+/vsVpoe7fflGsY5rT9wqdZ
6WiM/YGcvPbliRwUmEWfRhaAGSjK+e7mdFv1bON+HcFILukj+2EErOMX8GL+wanhfeewe8E4U5jy
mDeuog8O2DqnAXN2PMjqSqmWHt/hyAtA4ejZN6ibK2jkzxYXn4t/RejRl4tol9q7NBSntQLOGaTD
ieymZZ64l02fiJqOxj1uQ62vl2RxQpr0hiN2xfhEsKeJFSnCqrSVwvkuQuywbPOqtdj1S6bilrHK
cOV5T1wI/Dq/8XVOfA4sJYI/Pi8ISkWxeS4zMkvmG+JabfypCndIVQ6HYAzcPRfdrQwqSwbN+4yC
bhiAAB1woeEw8wx9UsRtjkDYLLIgSM2rJ1mBB4JeI+hgUKlBCwULKnXDYkPEia6aUuodSEACuHQ5
8xP+cqAcsAWo5xP8Bxrrqvd0FR4dk+6M2SpzJsto//ziAU8VbFWtCtsOuWRLESj+3+HIsB1Jggiu
FVAw93aQ5uP2DaD5i7KsZJnvtom2Zk02133UedkMkgE6yB6t12tFCcMd/6O3mOagC53T+bHChSv3
XjWJKap0MDlta52ZviV3TMar01fbshqvusGEpyPx36Cr05wmacmYwc+8TlonOsxuKn5JpvEgyzl9
6AziQYfMluwNeAFq/9T1Txv3+Xplo/nSnqtIKbN5+0FEqrQKqSMntJ07sR1NhRipti4ZAHZdTmi5
34+Cp8UyI6hiRpyhUEUgPtoZTB95XSYpSQY8q2CuH9acNT82ICBp7qxykQVyHyZR4pM7W/1sf8u+
TbfMIqHr4nQ2yHp/m9oEI0xq7YWHL35vJxEBQpotBm0Dr3yMcCJYRRmcoadlBV5IITohJKGlgX7b
22EhpGNosBPidDizTjSI5yD8VVsU7qNN39n5Yx0Ujez/49f0nT9Y4xVfZ5taohOUDQA+YSur8N4H
L0zwrtSrDWCixnuNLv2RMdu0nY33wCxFs41zYV0jx1ycUs94D/VjWwz4VrBu8umaY377HQ3cROj+
maagM/pYWL38diZdh7PdQ0tTniqbkhjTPJO6vt+Eq0RRr6sR1T0Z84gjiSWUzcQRLcoPhaehN4SH
YQLN1i158w0FesugSy+9zNLkQhoM9PgJJhAGfObAIpmqKuR/K1RuQshO/OVko+L6LAwtk04InxTW
WjNzxyRAMHBxjcbNY11NurZh0y5Yguc1dhynYBKdx7lKX8ZVhpPBJxesEJUodsk0d47kZajfvm1C
1VD+t/nu96GzLvJNzoWlue0A+J+aK+S8EzXsp8KeH5hZvUM9B0gLN32WwItQgzdn8tiV99+Z6HPl
bOCPi1/l4sUdQ0W2+MHgYHoIqHJaLmBmV16fxUzDG6paQqBPaPv8B4YLzzpkXVPlKWm6HkgCi9bi
OnNEdj94oGweTUkr9JLubKusXY+OsvQ5i0gHbjJ1VYNp3c9H4FPp6IVOR64kyIevZR25EOJKU4/O
jeNUtSu+XH8q2UK+k89PsSPhZ8M8dJx2E9cqDAEkJcf8cRsVE+sThJxxZPPT8JG6VlWNPhJ2kc2w
4B2o2sSzqMLLdKzBdWq+trp3IVk9tzj40ZZn8Rl9SQlPL/XcstMnOeOynHboF2vNw4S+wabYSmeL
g2eTHNTco4n8u/TOQBD79KyyxCZNu5nSzQoF8J/wHwyIojYKoUQ/wXwelsaO5RQWKNUqjGgZmbr4
XlLvNYDJO/LsonDFaidtBZOuTjXBqU8EPvPc0S4cM+aCXOPHO7iRsBjjO8wnSbXnvKp3skyAfZab
iYmgchrXk/8Fiey5q0991FFZSFA70JGvf4MYnTmC0bA/LYg9oJmaUtKOSawhB88IFyx9UgGoQrjj
Ryij9FBXw/5baik9mKzDv4oRix7gBQdiKPcMkTRTjoAmO+Lpv9wy91UgHnE8BxGshPBb4bEGLLOo
hZsW+xgyF1m6+6ARdKUbHuIVwxDO64/Mgv9xO9zbB1eS9km4/6gRRoBrjPhPPLwTPtw6642J7sQe
GKwiLI7uQVkpqeYHXHskrsZ5WuwtNqQARuvWvIgF2r+Sw+f0RO6FMmK+TASx2d4qLkWHX/8npV9V
XWQqCZ1ioH/rx/K+eFTNg/9z17SbAouNRrJwAvDXOxWSMLJiAj1mVjCp9cQ++XGpT3bsf51swDa3
IOUB2YwHF8dcdD59e3SwRmM7CRfboq7E2UKy4lEFfVBgoiLx17809qLtnpBbydAQOf6tclVBTM9g
fDepeWLFqLEyqcOcxQwjd/lhTmO/LIQwUsqcV6hRDXCP2gkusoiPuTif4qk6aWzkz+C2Bh3o3xHf
+MPxr+snHMN+UF2xXe2PK1CHHnXAUND7+Y6evIbG5pEoGUp5g3V0lmF73w7/vemcP8zez36rbeMA
voPtwWVq8RSrKV4NmTY/K7MClWHpXjYcX3s2psEEkv6czsrRsuDLk6IgbIFBnxe0h+dH1j7XRAe6
GA6hq8jzxUCdO/qBVbJo23efYmVjGDWjxUpfa/GgT8+AfOlv+j9X+2f8ABfXibOsKiREvZ+b/LJP
tJf+r1PGUanZPo4+2YI0wxWI8o0jdBbXq6vEbRtUB/LHtgeNBrD0ITOcUL3HHLXykH3JvW6lL5NY
sRtf54ky4/Bwk7JhR6Ozl7EsVwGlVxyhUIcLF88uhqPcyLIATGYcP0+t2mBX8DSwhUqlUEjCk2gf
OslhsnOHDW3J6dOHm855IdTBo3r9pve1vfE3LxQZ78X7EkitJ1uurt0fpzt8X0CisHGS0hXbFhw8
Koduw79I9UaOl9JxsU2tz5llMJRXdIOcObgjghvctDh3dabDCjZ7agvom7pPb4At52XFzPEOx2KW
+m3YdAeBT9sp48z66KsD/ZiuCH/ofqkUrwCUDAVkNzWMxgrJueJjk5yyq/D6mY+vgl/JATjMnkxP
3kzSKHz/ePx5ggbKIOxYPFfPnYFVsyyKiyf09b8Bk8CqZT3ZZiooVe2t/tb7fy3Fasg2YrSHD0OD
Yv7O6xZJt1h/B6Ukrg7G6hURAlc3+GkceM7VEdbM1kVK0Pff+zPFa3UFbjd/PJfoi42hXjHbcXwO
0qbOk8uqX92xn3rQFwhdbrGPuKftC3SgGuCMA9yZNuswyFxMmE4NLPgkOGCWYf+COwTJEfkKZ7eD
R0m+x3wpqpCW0yf0RP+Xk9tmQYRmlkLLM6eaZHu78cidHUb20Xv4d5Ew/gQpNjXHnkLHkV1BNFuF
E9oq4dPuCVrYycdv8Z6wndh1Bp8vZxJdgYM/vkPFf+Px9LzambCcXIwSyjm9n/NOBW0+2fgUrito
9GqBTLv3P162oTB2onlwFWMkYu5F5p5KE7FXlwMWIrM7y3yO7CXNwyd1vNZy3AS6JKAXALO7f4dn
LjzvlwmoCIA1iAd6pmH1HOPMu+bc29ZoA7jAk00pBLsJeIYwAyCu3fOV4s1QH/c5OCJ0fcrLS6ch
Sr6ogKYumi6yyiw/qNEKRCnzsIL1payNck4C4oVOTH+eZ0X3iE7Heohu5wzlCbd5Oj6nV1ozQyCk
EwNyzuL12qutjfQRGeXtwKa7clH6gdd82KtGCYGSmpp4aIg9p67ofdqdpSomIAaKbTEZbahHo8HB
kPbzOOHxTLJ1R5B43xoyoDLyHz1qbJhzh2TmbD3uQ58fXlrVfQR6T2eF1fBy+4PhaPsXybgyjAWd
+M8s+V8AFhWps8sebQrIy+Mqtg0TqKmrHH8kfxniBeyhQYABYWB80QIFTjZPIGDFIyYIYaLs+Egy
1dVj8y3PwCFJQXxd3Q3sAQK7d9eDnUTlXfPSuCn/Kn6w3sR4C3wKwxL9+3gXzig2BGz5JqAjwD2m
5C7VRPHmx/InxM4OyjqEpqF/naTDc9R5AjzDsCNDA4hlTpScptxkpW0b3UcXswcptXxiSMxstQy2
F3ZX3kiZFeh4wmjrZFuCVTdQ/VqWjI1vRQRlq43kZIA9l+jNPJ5FBvv9aDhfsyqc7WV0rbXzig9K
DHF91jsqnQ3ZGeC3+KXtBK6gKTfVuXMPHwtN56SKJ4dWKZRAB7wv5BLGWb1L31BuKFCt2hLOz3SJ
/UAHfJNAsicvG6loZ9W9HKP+f0rm8P+Ft6E9BY2DKTkwXMnBoGDLeNQd/0/1j3rgxiI/PkXSZMfs
5cNqrW5Ttrj/SQJSPJdek4CRs+GvcVVOKgp98dM+iAgdJR/vZenPGeOBA+7la2htkaK5QJ9GtcKN
Qb+AiJwrCOeYSweZt2Go/0EKFkdoOEZ/nSK7KIOzGJ6KpLQNlzYhBsPECxDMeQFhCfWEdw1Iu9dJ
kIaLe9myL3RC7ppp14sZoqMTbWPZXb5h6hd3byq+eV8i0UGnwM8pkkd1LUB+TJbagjJ5Jp+ef9JT
uZfyExWmLlFUnxiZ/hu94Ic9oSDdn68HKnuMOeNIlT3Cw7JPoy3+0GJ1s59S2motVDa4xETiPZWT
WHUGARCcl5LZb2WbwSAyq6XoydOd7H5qV7avbxeJZKRBippg92ZPFGnNh4KWP/e0DDoheJOqOP8r
T9cIrwPzrSSX1x1rO6HtrlbsLXxYF95VkM2JFfsP9vyNXcJMKJXBHxEEdF9jyXcMIPQVpLxmP8kp
dMamyL5wWJP3KgPwYzjhSMm72xGJxSMVc8z41lm8vcxX9+QbAUVGQxB84m0YxL6zMuTMkkJdkhdN
dFsvxSNGt5ZIgctRMbBS6uAGi0+KtVs96MyiLMfdSwNbpuVMVRf5UwF6g3kZeZ0vWOC5Jnn9fkFn
k19spnA7gGv/rVG0nzqLGZIZVPhTPl7w1mas64OXhY1ZFoQvsOaV+G/gCFXCeV1gRHy/QRd4aPdU
TG1IqGmxYApC2VCJg5Rz6rIS4TbM6Bzr7Iwkx458UJYG+Wety+sDI6utcNESseNc/mNXsPNaRHid
s+IIEWnuMLS0vx9S7vAxz+PZYuCqm/PsuqXdw17KNfIncxhFC+EogF/oDv44VilmbU/NKSLDLbQl
uStuqwiQSUrpcEdgmewLYUk4kYz6tJ3qWdDub5UY1Eg8tELa8bEXdcCkeaEFGO4NxJ8CYgX+Vnap
UuB0IDfroAViLX21Etov/Ze+mh8Epc52Sq8BId5be7GSUnlDaWcNCVwzBk3zhLaGxCsT+OMb5HQ1
QHbEUXI7zXVF5vB6jdMwPVuepB84dCdraUbXPuF6glwTXG4YvtwHlaz5cYB00W2ihkyEpeN+Fds9
eFIdePdXKZCnePHIWMAIuCL2lBNTTFrtNRVEeEfkCYVYVXValEHnDeXV917Kdgqt9tN+15APUXJ5
59gBZRSQUaq3WQ0cQeJU/NNfgBwn3FEfxR1CL5HlHu+nFQ9BrcIaIVw90FAk4lGtqdKvdh+AR6Fo
On2CiH1wX5ympvYOLAJNdFuRDYMfc1IMQtg9KVinCy1lBcrnI1t+mmzlAxXnpi/fBdN87OTBJNPx
x6F+RJ/mFHVPwceTy70c+FbVR7MoSzeX9Z5vQht1wTmx1uXTh3M6yIxKxkjWe0iwp2l61FmxpdK5
MJoPrfJCtWCRPKH+Hv58jflgpElGYM17SmK81q/wUoLR/aRhiw2ufE8e5TTjeTU4ZbOS6/fJP/Z0
9Mk3G9lPBSJ6xY1di11F16kJsk/Ys2H8ns+oEu8KV2W4PjZWRqN8D7RZCKzNNxLaML/v12jRj/TU
/4QFH2iyTdb0/5YwkUQpXmmlzFy8oghPz4GgJhOPLnST6sL16kLs0nbeq5WPXN7EIvKH63yaD6E3
DZgWYjxhoOlDg0d7hTaOQ5qPAtbj/U37V+vKB2MwCQ6kUReZfQT7EF7jm9QnJ+rqYc0GTp7fWHyJ
j7vK1/s1hLlV2k3builIV/IEUePmkHm0Z+Ho/Nnm8vwu08SwAAs/IDW7Xg+/EyqbQ4fZ2yhLeWis
HRxOm+eIYMxLPKh1lI0QMRmi6Gh84a16sAKcUuIbNUicdy0DZMNhUUkNiPCMXyI2JqC0sCA12UJy
LDzp6DcHS5olpAtDmC1PajvMFmg9T/xpnBHD1Z2N9LKbccMweCbJcywjlgFS1KlLXUub4Uj85E8H
fmUSBJCNllLVweWhnyH6+eWQWZU5UqplpbZD/uJ/zHXV/ejKCuW+ATQn/06IcYC/5m3dD8BPSTsU
Vzckrq9QuHxUKtJ+xbHKHRqtQLCiqKY2F0Gi1u9D2LCzd4rNTLUK38+4wYzJOrt1bYaLJip3a4gS
ogqKsOO4B7/k8nOnv9uLJUQ8NA3dEHWLHlH2ahOXnlmqbiuiimdPwLtKrQvvknvMhzxec/pl/fKC
7Co1FvB+1rSOaCgPTrpRSm8YiFwdWOcqc6wuPUgrAzOeQScttS57gaKgmKK28Ijs1niB9pUrPtB3
kX49BbM7Hcaii5eyUnrz1u8uYRsCT5AS7Iz0/ca/61HyrVS9lHfOdLVuc9Rph5fpaEfK4JAXqBVX
48shsstgLqJFlC0oZEhJ3osxrDK07eBt9z5MfQhWMjUM5P4Yi6332rS0Q+VZdTWUk4/gHFaZdrq9
Ov9s4A0xVY33avMiyqgEMmYgcwsoHI2XD92ACyYpbgQwJqK29Ib610g+xBNB+dliDjv+E/QUVNIe
whKm2Od8iojvRBO9aCGQCXUO5y+/YwM8B6E9A+Te6RRU6gGwGnQESOBtJQjkOp7HjxcTpx1Ar7fy
dLZAjcaRe6sEuTWPxxF/wgbfdChZnpfBE3NWd2SjpMQIrhgELQ8lgR4ZEFvMjix0Jk/4z2iYFJz0
ufQYRHXrGVbSUx5DE7vQacoXtChjK10w86kYzuawlViTGQ1aCQoWe+cbdq3suHqGd4rj6r+UERHL
Th6B58HC2reoTF9p47MBTsaxFWdGzL4hsmN//M+aZNlmYewoFJ4+E1LnO1Yu7AzHMUvSFaMU58fa
yf3zq9fDguDyiyjWe8+HHEDQoDqPNJa+R3L1j1GsJGiVwmO+kWXukz2RMsa2gbp7jXhL6npV9u9L
G4lHIzD3/BdNOA08Sa4ui3vNFO7m7lIFBlrDWJhnnW3UQ1bfiXrACzg8Pjsi9ZiDUwD+qrlAz2j8
Dj54TniyIjFbcMAFMNYyc0sW9eVpmeGrcKRqnsxOo67IL41s7p27us7A0hXbExOeWnyRbk9UxUKI
E+QMpQYDB5ZjFe0a0froM2FEp6dmEHfmKb+D7zyA3wrlGBQT9oPu6jSF0CBt8/nKaCwtqa8zXNX+
A6qtqEiFg9inXLhAfvQcTGM6D/At8hv5AmUjVdSembTcfbJAcxP2zJJJoWuocJx4fzLy17J7XH5c
2Rb1URBWJdy4hIxFdvR10miVptCTx2agOh0qs3/sxOvl6vds4JUwCtJ3soz9CK1eIOBnML53tM+o
GWC2CglNIglmHAJHOZu8LXoo0phgJYcSrPFqVAAhPqQZKPbm/cCNx2YyLB4R2IAHj+m7JXGxyqej
j1lQhxT0H4TyMgjKZ3cfacguH+7/n2uiaxKcVlHtsdnvyKTfb/zdaFCszJ6A4QHR6P5avuDwRT2q
+J5kwhB2SEZnPl4HxU2LgkHxP2bCGCGfog3CcByIG9tMmXVG1Gbbp/JHXPHgkbRfKX/QlveAxhR4
u0uDiWt/mUVdrVnmSoynGyskkR79HXVr3IAYbWNxxj/nmtew1Ref8a341SWIeB3OXWPCNzNvG4uQ
hLZmRKGROdtbhVjm1jeff6a0NQiu3cBWKRBQZuSu7c3kAeA2K4b+1R9vwWGEkD4rX1MHNOx6QT+n
VKq6dta+tMYxlloD1Ck3N2ddSYpyfjrpfxeFFYpstEzDgGxfhSVjzMWUgqF7rkIDpPq/8x3dvcB+
7OWZ4EKiBqQEGsS+2iuKPXMpNCa4qnWULRc76r/XFFh5tcjuRLv19ywKtpVuZACrzO0n4pgkbp+j
9l3hmmtkdpHhE6gl2w6VrPpZXh/AGKEeTdXvcgeceKUqoeHP1ZUhgdLQ02qWQn6Jo9sdXsy2gcFt
lLaXxwt6zAwhE/4L1pK3i/QcpsaL5mNxcQGui4abMT1pc2iWHryr5mZYI+DkN3V6DWTQ2C5xKPUa
0bFrsk+Gfcx2Zz3Q0cDZhmchBaPxJTVupPVyGh9LxFUmOLvoEGpvNbdzK7m5S77aJ3EfGYBZpXd2
q2JUJkwfSsnwbZNtJtm7dG4Ynl9j+Sf7xB4VPER+1bBiJyrF9EZwhyM5QpJU7wa3oYKRsBAu/yM7
+YoYuxbs2FhyV0kPpaXCWVjaBMzq+RyNCJGFXp3ObQ7EoEuK2LR95IezKzQOyvIj9XzdqIR6oMRw
ndkRnVxM0jWmKVm7RzkoBKy3igreUHnO0EKK1rzz0izM24cx8ulDuJQbuocNemcpb4KlfEOK9VX8
wCg11LvWlIiAP0cHDVPcvRMn5x6nuEyWOHZg1jjx8QT5G8TSQ4vttefrVOwqc2T1YyPmXSaPiu+L
Q3yXklHSwQegNdRnB5eaYytkSptRNigowntCF/I0jqGCMDyvPrnAp8eq+hVZbzPiGuYRUJc/K5F1
0mdZMiCEJ8ifWJzGXc++YMIotyc+2A1cLHl9NQylTXyEWqidd/ugEunZ/3Sj9FCS3RNFs8f+q60n
WvvWl0o6cYr581/2MzuqD+hpEoJDRVaotgB1bUW41dXK0+6i/SUVyo51ELhZI/zxed0WXehk8J7G
KCN+FGTSbg2uM2qIUrcmlyPrvj7pO3lM+OqsrIQOgEDUEiRZ4kToqLde6dx0esQeXYsCRFOptZdE
kUP/DkkXX0daQo/5MNsmUXzPcEJ84/I5ZUQZAx7dae6t0+P4VAUAynrhEEVZm/iyN0wx2R6BDrLG
DlPX4ll4JoBPkaRZZbHaHA9NLUx+pbgluUMDrXwefnokCubgGgSK0NHSNtD5JvKBmkhYrxxbcA8U
Zhreiomg5P+20RmrUf7FMG2/7qPgyy5NBm4E+uGVqtWI9lxOtLPB75wLxhlriQGTPurapLq+M+Zj
Z6hWU+wlMrQEwDVaf9hO2m1QCoSuNHHjZ3x5M048Cuw8E7pnFsFQsQ76yhGp2rrK8sRiSbsdR9Te
Ek3A+/kRJ74+yLuKclb2I95QDLNRIXWcHefzqOYrdu/VKPYKbBIEaoX7xYDS/TD9gMTE7a0Ivq85
r2PRrlJBbLgzbhKFFJA/uwXBOQwMcHrlhXF3QsnkfdJuq/oLxttSChSpmFU+BA1P4HXGkj9tFF3O
LnAMucTsQB9Ju4zYWLbni276uJElQNzabZ07vWmGUqtX6VSZrzfROJf+thxQOFCjhQCKPIVbOCeL
/R3dFOgY4/AtpWXsU5YEOKbKLekpBSui6N5hNvH3ezJYYeE5ZHYD5sYmYrxqe0aNGMh3cBPEX3oZ
S1vf5BZLYHY9v6WxDyUNk3OPme6vUoJy/kTo03peghK7xbvFQ4sIFojpUvzQV5khbv8cSFdc3Qjf
ttj2piU9ZsiN7f7hLtEE50bjW62ylodnbJ33a+J3vLTlJ+NvpnXO71Zi8ZHOoAhN8x7eOHdi40rd
iLq8bMc8uS+to/V45KyEKYRH0qmOlo+U012WNxlASNCPLdp5Y4hs1HZib4V/L7jagaHI1NdxTjoN
JVZtznf3ZH9mDvnE0mbDTdBv+VlaCfkpNJE89JStXeYEygyzGzb/ZbmccEi9S3NVGWA0qoH6mF6A
x6ONJozGHOIMLTqwI08RkuGSP2YULA5yq5NsRso90Dq6x2K6DqRxj1OokLvZGJL7dxVGnHZVKSDu
RksFTWZwleMgarT24dDPxs4O48HWVi7grMiAf8kDgbjqcTjIPkgIg5WykCKV27P3qKXm0NmrJTwP
T+Ona0X6ntvSyGnPqg6tatE43WDszBDBNgkJvO1+WvLeXAU8xWfNITiWaTU9M9NmFzmp5vP+NgZg
CCy7PQ/wBoLb0J9o27GXEtNdhqW4IjA0KKhZ9d3GXUqv7wvy5BcJt2MMOgYAariAJy5TqfJwY+La
LCTisv84XT9JgqTfpfxTJVXXlFMAk0O/0y7Q2SJE2yaloO9Zok/TFPLH9AG3kysiNt7ptgFOWNFX
S26leTchCZ6E2+o2c6NXxrDYmY9xfQuOghxlmAxqeKvne1FQYSVhofMEHwfSjoAnJsAFw8WxZzcG
0HuVi07M0EhJaiqc8rgh3AJBvItCIkTwxihNdyiFNj7Vq/NDWrWPG8Nnv5tbGoQDQMYS/OAEWlrm
8XBO5+So2PT3Bz8GnLZU0Zq+k7HLbLBAQskU8gnBPqej89/Z/Ba4Fd45iN/+XJIpj7HsFFdJYDxS
D9yLL+FfPUCurp7FAoHoaYX6YAyf6xJfv9M0KC4VlAgRRXF15iqOkMfVZFhKC7cL5GZt7oULk9VG
tdj5uZaoDu9wV30j0hByOiefAoPHCpfwRI6tWjCm4AW9MIpCMNZiSy5qwjwkqlcX+6D3rt1uZtxO
5MOV4WJqeTpufGt+V+E+gsXNS22bkBuycZlERVKkG8yOaeHErnCkhUfNFhIzCM8K98QcDtd4W6cj
po0wppJC7Ja9B+USwDu30/hk7zZXoYW57AkhJx7ttQR7Vk87lnAh0DIa98Fcj7Bd8+5DYogWvF8M
d1INJA+BrqWuU4urHFoTjZ9D9+DLQEOjSOfJ0TMhJnoUY2FBDuN2bYCghQFdYQ15sXObpisPzSbK
F9Il1FuEVIN26QHZmagwTsYQ24vXr/RA0bKhZDJq3f7rO26P/0xr3lTpapKBNZVluEWSB8I9Izcr
4jrAdjrNY/QpOOWPMWyvZ6BaueF4JRLnj1ZlGueVdgC+dR2bS5KGA2Qo+DfukGDueRVJ1SuycjUK
CUDDK87Q6t+2od5NwQQw1BrcoTHB5kgB+moICqK5T3RrQtzIXvZVsbuoqvtUCjxqlZDeCqBeulbm
nTFZxyHq8DFcbxWzD8vIJ1C/IpVaYi3/I9eXokbnsmAcpIENvfGUxH1F/sAUb5VIHpufjD2rfeX8
3hxXgUp3Fr8qBNGQ93+w/SveyUsqZjWtB+ywbpMMyG6DMGHM9sI6ug6hIM7poGv3Ar/tb+wiDzN3
6tc/aC2OZe+GatbR0SC+vqgh3BamxmYlHy/uv9vsP6JVZNKr2vSFPU4FmNWk8EMeYf++q/r3qsxR
rbf7QmWuJB3muY7JkwdbjAsjhuXVQH5uA1j9LowOx9mvZeNIohUX/bmZ3yIrZ5Td/nHCG5ibITVn
5HPkrhhNT8eFaFN4lGLcv/CSTcrSno3r7Rx5DCmHtIwOX86B3I43KXv9ykZiBxVIxuCRUuI19pul
JqyC80t+1qIb5vRoRK1+3RkBaFHyBucG6kyDAZNJkl872E6exu40YVWquZkbBda4I/0DmWpFGPhF
SNRE06o9QjqfsOE7SQol3/+T6tr4N06DzENIjs04oLTzjlEcDx7KMoGtgnl53PMBsy+pAsYPQxX6
vYxxxYaU8CoZYw9d3LtIx6lNYyWbox1VUCDRIJiHVt2q8P4jzuHD389jsk116x3eNmpCp2KYqAmo
ff2CN5LyMc0zm1kuZZiJL0stvdXfzjVZUZWKSdMjSHfyXMZ5o52Y5/5TCXV0bFL08XT0dDkoahJx
q3IOe+n3ZNcpj1MU8CS/fDXnxTd8KHSmEnOOzQe2YCBtErbL9mPWlwD8FGP9bQWktxaubKG6gbSN
8SnmKbFi4s6osmACUArUNEqEU0+kVs7100Uq+aJxFoXlbqG6RHNHyRQHm+sKsU8gmpEFzCY6jEKe
77YGUxD8mHVigIp/HMw9SfpFxFYYRdWPLNDJAf1bLagHJLI7JRyVg6xcJZtDm0rbJwxCcSvjreiC
J/UCyavAiS2nXooArqd3wrLeaXJwXtuQLVD4g+gQ7dR2XxwOAl7ejDgEWJMZqX1mE7HRMo0qhv5J
Qi5JCvhLg49l7CBJLKOyFfyzq3s7u1SST0vtPEOrufEFeoTUDRXBPpGKFZh3wpRQR3uQ6iIVAfRC
KZvczUxaceFkf8rkGTWcMWD9WjYZuRb5jPb1RZxYixYC3093KH60FUFbeySlA5mSyXzx8cjRF0up
hVeiCMb27kEU0idZyoLYD8e71aNaCfJgMbph1Ax67olOP17phxsOXccHfCp+eRTw+6VXbX+hOaAa
ZXwHe8BLPqf3jh3SAQc7inManBXIDmedUH1AAOAVexQZOpGhaqCb7+eQGT5PJ9Utv+HpdQKDD8J2
nwkfGgzP67oD0FH/Gl0S78B1+Tnyu7BiosuGEfZ7Yx8BukzTVQBJTubDG/hH1+t6aAhHAixdCcnD
xcTRsPiA7btJaHyl5HLEq4bY8KKJIO+hegk8T6TiUyeA00aI76PRwg0oFGyW3vYSDvmISFV9l9p1
51K+bs4QZV4/1ztYViL+CXACnG/ED4oKOeYpBGCV3jujWwsRzU6dsNTUgvXnCTwwSDcCwb7yhQGN
gK9502FQTQ/MBlU6/zRQaAiC7HmYzXgsa1yb5JiFz04AQEzR5Sgm1heVEWufFzQzy8miS9+5P5bn
oaPZKJwflR28tXz+20NZcI1f9XG+awMWoKgq8oL9flm53/YvahG4Yv2RFXgQ6k7g+C+Svo2uMR1R
rxm4xKhSdhZCdXZYxQ15mATJ0npkjMkNwBeLI/NEOXLrzDdM9ARO4nHBTBh6UFIDWkKAzwuGpA86
hughmxw93hI/Nl6weipEV99BhZVcwANTqAzR9r8vDarISXBC57Um8TWu3utuCiVDn19g4P/M+jC7
VrKxrOqZ8qSvppl5rZJ6fXLvutSuIaS21rxVwPJiwKULc1MZnSlqj9zup7DsLSgihfx2qqWD60sY
5vL+ZdEhYpKrGo6De7UqVrGz54xEQhTI/+FAteO2WR5HM6uZXF+A07qsU0+zJHeyDzGQMFAeLhWK
tfS+PmMr6qtQSXJkNsDQFZX/zk448+HlZE3TmNr3+9VV6ibvV5cIOjcGOcvVKgkeesvjsExm9wpq
Ia4yWF2mIKiBgyVW/BdIx9C7NATsXMuL3N/dOMdM3JueimxGdQoT113CGCMdbRYSXg4mTasTf+HK
u+ubxjC+e8xp+H4c4M4iDygcoKB4dRmQdPyttPo5C09UoedcI+g8Wd1ZktaTFt6uMUnaIlFDV3L2
a8+nWPcASbzcinfrb7nZ4L9nL5iJu/F/dbA4FToK5W2b6BHKBfOpGz9x/PCkMy+5NbTs3Dn4TtCF
lZ6ZzxjCIf7Ga+fWTcp9p8D+a/7De9WM71N8dzvpPQBLYG7zuSdrOOZ6XjGtcSGAfNbgUR9wnNus
yfl1PFfs1huW8p/JKdj2fxdgvaJpCKqJHDFByLZL+kYsFugz6JEF8ERMSQ1lQNMlZ2kQyx9B3qT+
a5NIfYUooJwUGnOoORqPcDnh9+ykvA2jaW6i1X9iWPGD/YEMUVZD3kCVL6kK9LnjM8bsDLwsblUL
p55FKZaV6p6uR6qnj1EY5IC21lb3vdvR1g0GMdyi1HooDdOzWS812ad7CFlUQqeTF4FkpgsmI4Ih
Umq0opfX7pKjAfLwtPB5EJKC5niftTJFy4LJB0XzOkzDrlOiNl1SE5Hb/bGcrd/t2im3EPzUiYHB
BeudDKnIR6g88MZQqt9mjykt0fCrd/gCCa2pJGhEjFby8eF1wmGuuGUIgCgtlzNUwTXQFcpFIQTQ
4nTMpQl8eJLn6b5K8jpWdU1Ia44TPt73HXsn5uzCOUHx//2wC8xDOhHQbkomPOG1ZCZ6OkphmhZ4
gFVHPO3WicFEFoAFsx96bo8lCpZLM42kPWWtshG15WhGX+O0OUtsN1qWE7HjGNhrZfd7IXjKKJhY
lV+xDtfn1aUcWZl1hrMxcQS/Pqsm18vpqLl++U585ki96PH20uUhA4/c990LxkbxA23VaQoEFLn5
LkKfJ0FEiJF7nrmps0et5La30CTX/0EtmBdgVtDUXklgEPbT7WqYSIY3q48Rg1kAXZwCLoppic7r
szIOyPjWljfcUfDB1ZqOyr6Qzfcmc/o48X6s2+ru6ovQPO7l+zeCZHdBdnV/vQAobn2ln7YgKyWG
HVt4dh/EIC6lOHlKeF+hlhPRMCou6I4L3lirWeAgE2pGyESvTU0EPetB5MLjdI34CR6IofEH+ax2
nfU6d5g8xEmSzsDeWOJjlOKq2az9pDFhZ8nrBRHl/2bBGFoKyB2PcyihKvP0akZQrLTQsRSM5A3r
8JErV4SwOFhhWhJWQ0glOBA1PneQA0p+FX6yGshKaAIUZqpGxCD7Mt90Mjca/c4weMvXFzrnFSws
lVsYUTr0mFB74H18ntKCK3FyKHZJbRkFaOYXgvw2ycFhWvBRz27a+FQBsWbsAwOpqS4GOX0UZOjh
MDPeu5fo0mUN8KhXjiZ7ImCqyAgjdsP/9BGFpFz4AJRRnjSBOUVG7hcw/WtHFrb19UHuH7Jhl1D2
kNsV497rzIhU+Y2CjC3MHh8i4oM60tVrvJug7apjXUT/6WND+hCYEYlcwdUw01afHum+5t/j2xpl
YO4Y6nm1WnfVAmegFzW87QkUY6Sk2cvoWeT+opo5D6GQURSkGf2GmxbjKnXeX80vIVbj0uRKzYal
aKUxJiJgjnBImo+VIQA+m2+2WcswQC/V8JVXNbseGnEyLcCs7T/5DLH+2ernlf/16ePcxSK2wyiI
cxInqUwoCIV4iYmZv4aZmx3yy9gqiyKWjL2sosKB5hfD63gJrDgXjgF0YGxUKngM3JYaDJ6OGKyS
2+t8fckly3ObXzd3pQeMVrxYGYtZVGpeW5DDFxCNY9EW8YIY9M3kwR8MnBtSAKWAXB72DijX4mcK
CnD9q53hJJsEPxrMjFHVIyQ/DkpWtU8kZe/Bqskibfo/alRa2X4Ot6FN+ue9FHBw0Gv9COceu3Fi
UqAYsOFViLbl5BSrV7ZgT78zcKEfLZM45cpN8Ig7YVcNHJvQ0pQ9oas1+bGdx231LCkGo/YBH1nE
Vc4ZQae4bAlVvY+sXWHibk+pijMw1fQA0zCgX/BeoH/1NjJNmdMZFa37eir71TqBKbdq+kp9YPQn
6TD1J2ZZwC2U5+6ZG2BWHCyle+bhgTpih0LczXaLqyQxyNnGpWhHaR69Qyw7VWHbtiP0GMnpHqlm
HdGRaitaO8FbVoBec7n8GFNlGUIvzjaU0VhliA+AIiro8olunht8Whdb9hVPl6TE+NmCOociiB0w
IKATMxcG/ka1gFdxhwc/uaeXma3xI3WVKe95iH5ZEhIM3BsIaTyuEWZRTuyPUKs3QfeXPgZs1IUC
PgyvKQLb3pqo9MJkapYLDLUQBxAd+ZBvv8bLKgYSlBN384H7a9PrzZ2tSzykmu4CxGNK4rW62EVU
KLaEgR2xRtKuIR69QQXZU0YoxeZi28OfgaGflbnY249tNDaQ5yn9ZprrXhozOXdcPjMKYQFHqoDp
Baj3/SX3BM529JRuj+332xQblFP3E1Pc+gnLDAtYwwNfN6CWitpasUYBgME747DyGRBjl7seXFTz
WSsJKCKAqBMxzC617h/SqbtbeX8JR9AHcieRKVjHMSUraApQFk5YlDoDK1fkX0ZKt8ff460tOpvr
NHjXRkGYLdS0tYWSUA89a5tPGsAq5EO+zB6u3/H/wDxAndHIhfo5VJWWBOYJ/m1DK2OuLncwe3gW
kHanXJi5/QsyQ+6RaV5V0zoe4AYDDVNkLw70pnXWb++KH4InWJ49ECPSqo3k1D49kAeHM+L8meE2
8ozBijNnf98dqeJppb9kUwWZR5rMHRsnvbmmlynEUG3W8/IMB3CTFYgCtdfwiZ5vbM9hR8uICQIe
9L34k6+sHSBq4l6KYEdTOzvkNT36kIyHPb3tq4Bvl45T8X/JXL0dw51Zsv/RwzNvH8bhB8z455GW
mI4Ua3g//ZrmfpIdi8CprI6ctIxh3XwInGw2/w7B3dHifdtNqpCN430Lyk8NO7Ho/Vmk3RXGpvii
/8wCDPbycf9gVUuT0B8W1Ab0Yjqwi+UwdxMtEK7zG6La20IZx4+SqfhvFnyM0ozBBCzujtfPu2N/
0mH5w/F7O7XFyHS2h7e81yy8gpvloYjO3SA1HG2Bvr8XNfU876wpG/oKa+v9Qf6YCYUEAX8aDaaJ
an51C9DykzfA+F+KeenRq9fDcVNZHWwX3FPgymkctJNuAAYjtfFJO+h3Ka7yNE+h5n2Zd5NDtiqb
5VRBwTMDV897p8PtaDZ4l9Eo8r+wlaEypfo8FpM10LiDsq+Z5MaIn/7zTJJ1gLYfoZfdgxVi4SeN
tLuIs7ZKKuhT7BrTabS3aa2p1d0MNeTOIierlJH52gXWlo8cEjxrZMOxRmwn7UrNwhuFqijcW6eb
RMPn88wRiM45nlXiNpdw5v6lt6Txd5o4d606EHAmydMLG5UuyzQtgrqtOf0fm8lxGWQ3PaFwX9k4
RP4jHM65dC7LAXo9kbKxEMuY/W4hQ+PqZx07bpvlDvKj1+PGONhcELfSDIFTHMdiuo4it8dbq7k1
wQTMXawVIx03uZx75+73aTcn5b8q5ZjNqeM9PLGM4SfCZbSIM/D54ejU4I/VTLdupZh9eF+3pKSF
KCtf36nxWLDlni/TR1WIOPl/u6nZbatqrjd6kQUO/Z1u0fg3GtHz1ElIuBGZfTzeGZ82h9zpq1hA
0GMMwWy39/+5/1cOaueLctwM3gtiXcX7vp4eSRJk/x5RtNP5MKabEtMgTjUD6Yv1xNhNKiqHJxMF
t0mSY2LUjZzsuxuGx9EdyEf554nmGez27UYB+d3u5ZkrDGSujg10prhzEdyC+y5pfNiUbMTyP7SP
dIKKrwEOJfdAlLDbJxmAp5GtqOve9SYlk36JQnwCsS3PgXIs8b9igybj4874fPKjDQViZLc4NKcs
qN6v5bdUChz2s8iBTIyHMhKYXxFa59YKIX0gbhPD+R0PNqK9xHbR9xmDEg+j0Fqzt0wSIbCk9FJq
+kosJKp2u/+7X3hS4k6kxuYCHc1Sr0NAyO+cUiVXLGNmSmPaEsKyl+o3x/l5TYQqOxLk/wS+DImh
A45uZ1IOw5kBPlwTG45nM2Sp7RLyWu4PUYqLAfYFcpCEZok8/QUpT/a7Rrt8/rXHFZFEDqPvA9kA
4EuXbJ/H4TTVTRZO2Qwo1fU+Wldme51Y7xfGxAY+u0vZ3fDIE3HUIyD36Ii0nl7DSUOZx3yywFK5
6x0cGpUg8EqyZrchk2cRuWdrHsFBdzVljarEpeRgn/XHDwniGXL42cM9aIVW6d06byxBChi3ko1O
dHVt4HD1YeY1TwG+bx4imKSuFuDwtDywgIQSHytjfgPYhZdGHsJqENtk1lTGveSbC8IGoT3NLdqx
ge87JgkorTvmxjGLHPDJdPJvaw+nwPcYlWyM0xNLmRjPWCXe/XwTpLfwALS0eLj3aJFPtGufl20E
lHLKQM300rsNxrNM/o+AXDVsVcFSmZ09JyWSKBuP1HC5qDuFNSAtl8ajNONFdj9yvDL4HpMufSwf
pJCnYDsd8DarbrO9LOxTi9OSV6pC1nJ3HxyUKeACpYUijIDvH4Kulb6wpV8Y7kom3jKENlN0Jca1
RXpTYk8vHp02bOYGYTD34YM8e0JuogKMnliD1lCL/WONYb3v38H4R6kNkgYnvB8yVvei1dnJda9q
WoTU7IeuDTQyZAHcIx2zIq+hT9yUv3FwpnCiDtO6Cf0Cx56pJCqG1EO5LxBe8lDAlUoP0n94l2Ua
uD8V9YW0drdJOHLI3m4pzYJk6q74hDmM+1/o/eTtDjCLqCq09xexfTdhl/HMcBm4FvVIlIOtAmfZ
ZPWiJO/ODdswd5jypcIbH8N5V2VA8pGXoU3QSguUY3upmPq5warXIDsWWgLMXzN5rYJSFtMJpSN2
kQjQhrrx4RoJtkCVY2cVwkcgtJ0fTfge6VUUz8ty/4S4Ihb54OIztY9juje9qc3TXBsUeFDnazws
fc236CDnYTTqd+WYXIIVzmxNyTZZQCJXtcaxNl4eDIEJf2m831hoIQH8GyCRKVoMUaZg5UPwDXxF
RIz4+1ghkV+ywTbzrCI59Qap6e/4zSDVfQp1N59OOXH7MiotmECdeidMDTDLgrqsp6/jCy4vUHZ2
QKN8X1lSANccE+6wOtiZI1tFnw++ktD3/HV7SnY7qd/P7iAWZFv0BZIopDN4LbAXUULjNY2C6c19
yIA4ZPiuZ5pf/FuCgLrcHPsy2fU1TfBm6rCk0WM/Of+Q+73CbJJnelgj0XwRUj6SLAI/C0MyFAFy
E3OX28B6HLqd0Zt03flW3Hg56ctuC91Zj6k+Q/YWilrHZqeRrCQIANBDrfD0uoJxNtJ2uVDVgIMZ
wJQHhqxdFgsbkOFXpVGkdM+pqzpmzKcLs918O6UecMSVyBPg0L+rRT8OnGV2t2f2ZvXlCFQLRamZ
cHY/a5uGZ/NZJnHr2U7e+zM3Ftrgwz4g0gspMRXDSjB1RiPjEybM5mXMKJ8UPxHoKwrMYCLbCKIW
MziY6r3QPmzVHJwrODu4gQ7wxaSydfdrdHVfQg65lGycqSnv3lvWQnjEr/x+zD3fpMxQs+LV04NM
LCIzqeJBqetY8MVtNftyntyICKDFQcmnmPz6lGnTCvxBnKTHx7jW7ne8/MTbLxULET9Q/VPFf0EE
TPLvKYLWrm4WqiPv1wtSewF365esiTXb70NgqYYx2BAiqkl0x4i/kISoTC/QqIgbj8l+n65/sAhl
VnE/w/Y/2AkC9miHPLHCddJ6FOByNdjrahAaVtA7a7RaPAe2nEgtsJj3xDeaTsCCfMiuRtF3ue+m
jnge0GNPtUOrqdVPiTZ/HhD4mG0CA0n7eLk99uwS8e87RH6cxDuTc0IdDIA9WbEvb4QQ6zDq2lGU
MKChi+JqMzD46zzsy5qKoIIFqWf3jkvUK7w1a2imb3zsotZoihGBzc8IGWYQ64fMSygkN02EZdGH
jGFJEMOGBxaOi7jOlprXxqYtgICNK7zHHQ782Ngw/nFZ5SsMfqkRBU100E3RCTFgLuitdfV6/Xlf
45yVSZuYPXeD4O5xZJDuC41/g9QdiBhNo9ah+2gvM8Vwhgotftjgfnhbeo+bwe0/XLI/8G5i8znI
aHkNJKzTtG4hTmITIAJP/7wIFDMaTm2ui01qfu3L5AxzDRRJTHhEIn9xAsrgb+BbgoOmydrm72vM
4YaaiiOUFrSa4Xy70elMNsKgelvtNAeGk5fZHRc9kgpNuZZWAdjMJvXjzztnNuxfyDQqKFUbGlIy
QQIcCryqoFqQCtDDvLs01kEgH+II6jhbs+WE/19TGgQj6w/lr2tsVgDP9+rx7IavuovN3mCUrUW2
Pd5Sr+LWwRCDn6yJvF/syvyHyOqu546Hdcf5mTfsOSWi9foGIiZ/BScsjTmuvyij55vS7yhf7TSD
xHGPQ3e9MumsyeDj61XBRzjg8B7+tLxc3MG+aF3kNy+Ow9rZFVZ3tduicZeKnwo14OR1u7awhl+h
ZFSr+Ms3zNNxP4O2dSd9v9VGzp9+XaGbUPCr/7wMTUibysj/1Em+0/5unXCjhjRQp5ZEsMVKXK92
XoomVxAEJukd0HBnVYD/CTsngfJt9WoCzRUXPXi1W+quEDS/OV6w2sbEpttGjGcMkrgfvvFo5TlY
nyLRG4pAt6WW6BEyH3j4KSeerMCXozDqzlYOTuoYt4BynHJZHbfELc70WWi86FwfKd32X8jKacdU
k2b8ZsmnpIEmrPZU6qoVQrpkSgIrd4B73KakGleWBNPdNdTFm1Y0mLgnOG2hf2o2SAPUFJSM3XXB
wmeWpTATR8EC5Wr1m5AsdqrqZdKY0lh6sl1CDjOjpuP79R3ZIIwGOtq5xPVkg0H38HJeRTuaYg7W
bAK/IIlJuMu56+31SdAyxzEq84b9PZgauFmRvMwFjcFUj6DnAek2gqLpNhvm1VQg5Aw+5HBWSp8Y
gcu3N2dME8aYOsuy/VDSAoE18LkBbTzNilsymQj5wFo45MRglTic3VGdWh7HVWyTXhFL4WXJb1MR
cQRgy2bNA0Y76rxiSNjmTCBYMIa1vhrKfxCEClUL0yUqUh3DeR7v1lUfDmx2pktSltBz42Pw/C7Y
1cWot5hZsLUq5D2bb9lHzxLAgpnEcfuI/U311HSSKfInWZJ7q/pHPMz+9mop4gjbtVMPUnMApVqb
KzqRY7EE5TAInLq7q1ZaIENOre+y8T0UzfLsYdPrTHxynUvJQv75tSpeY0gyw3Nm4bgtc/Mk3OQq
SOKCmtKm7l1YOMFfccjyVaaEMY+wZBrmR/M6jZunp4f/IxI7JubeZ1qog/2ghV3JWRNSKDMk52uY
bqopxj8a9JhRFW8MbS3Y/P/YqAxq7d9E+n7Et9Phzo5mmHXwIRv/wIIjeawjS3WkH5Fi/jnnzlqp
95+o3RTWnaysPl/sJkoRH3fyyFfDhMCrSRtoOf4omlWi0zvJgGnqW4GEBZqIRxDvk0OoDkSw0GSy
SWmAn5VLRvY8OEPy6L07sYGrIergiRjVojOrdw87F0a+EeNBi66uorC1yVYlYx70wGXFlO4Wi0Kb
vx3Cghblzc37bs1cT2IL/eymjPqxggXNo2QW5UFZqV4dV3q3i/sEttzrLR/8Vb0zSMyjAGiEY5Ku
hU2saCgjaWENRzsmDJSM0E63CeByxwDkq5Puk2RDgc4bQL2fVJK9Dtd622BqXneD1+ASH/GOvll7
lumtpNWrTZ5CpxCGFhCnWBXcTF6ku6YTRBfVcyWH4PboSV9J//in8fQD6II65JazZ0ath+cmEKP/
zhUxOvLSynTAsJHEIQDTzMxcB6LhSQ8lr7Aa4++QzSvd2pPFq5Z+4fcYPo/3O7g3qaUvtW+6aks3
hKNuQHj9xSyXUJkwKsRKK7fbjo5y1AUIfZlezysN4RpqMKr90NkgPcMi+7LcB9940u0f8LLZoE8u
QC3BHqiGvYU7UfW5njwLUTZbO/THlVkW6IjC7bDskdE6ZZW86W4i13E/Q12AHljfN7u9YH/fBIt2
5ZxhoR8a3PAk+YyCEAyAP7baCewo4xICgh7qxI0mZE0/0rEm3+coeYgB/+K5ip614ecTTlZ6tj6b
DDo3u7gh0Lh2qrsHFDh6z+QuLztjXFvFxIliTbufzG3l4/nBLXbttHkQ16RZjHXoVfhabdhVj1PC
tEhfsB4PJzkHX7BJ53ptIZcNR6QYez8qDh/ZpeAAsGrveRKNIQSXiIijl1n3Js6RsMzyA7vvujYO
/pioF0E1l8uI6II54k7W4+oV8mILOWPkr1K8QfpefumuaoSBRIF+66q1IRl2itc6blJDECcnZOnw
TQEyToSEEOG6FLh7JGel58xYAL5+JVNvIpAOW1yOEv+ong8Zo7/nHhS5T8NGNXdlOuRxTbQSQrVm
iTpJR5zkA4AVx16UFoZI4Owbb488PLfthb/ifiY5TPFWIWnUQlIyu+epk6U9QiEVVqOcOHkWQJ2U
l9KYT7gv/B3wkzUmqsMou9fzLmtigf3XdcvcWuvRU2MibnIfpbfsurl33yT6jx6MrXxIeRMCIZyj
kAqbm8wS4b850r8bsVXr+/f+qbavENc7ErBFZDkSI0vTM+EAmpDgTp2vdoGdqmUDx6zjMHP9B14q
5Tw0i+bpgmoHM8EgjcZKWtdnn/sj6UuR2BxvLr/kO6sbbuCw2YIxhsQua1TRBUxaOD7InrsG0FLZ
1L6skWsPb2Dzn5zF8vQ6hDTtLaG+R7N3+R2TUW0a7jfkj04Kbb/ttYlKeQmPY9gfpkBH1p17BJ7c
fMWSmDs7odK5VvASN7rmb+zejh0UCyvreaI9/wkX1xlJ0NqYL8Ihic3Odj5HzFOilmf73zmr8nKH
NpbB2WitDlnbic24bPcuIpTOfpqX9vYej+4bMNFi6cyKkigVW2f7SFBSCFO3i+KA3Mj1tuwJYM2D
pZ47EIvKyy3iMwmvOz23VcbJ5DIorjj4+H46W7GlxVH+JCoZ/hVa307ixLpqwHwMu9tzeo6+KY/Z
mLQlRY5EqVibnS4rbQi1v4ssMTZ2gG4Ce0XNEWkPb4yAXv1/2D6qTZMc373p5G2gdHQaSGW4wKtZ
7JutNjHdmLD/nyNLv64gbh4taxurvI+9EFt+Krod6eY+jEzjbepvct9ekH4gWm5hwdjxNVEo1N+k
KSRYNEZ0kvm/8mr6djdKhQUgKHB3CSc4W9fyV00/8nylBMHMA8wXCH2LGvLuARIpNAbL2/JHozTW
+5adHAQ1ANWIoCscD4SGeiW36IMObgv1wDPz6wBnSr6fR4e9PU9DKJrUqGS5wZA7T9f0CgVmsl5u
brCc0IR1qj0TWJdoo1K1h1+SpYDlf1rNaZyir47yRiZxfJBiOtshpgf0cVRuKWzVkSk3iqopxlrO
GGfDnEhKiQeYgAFJ2EO30RcGCuvfgRv/Q6WkNQXUVcoaEfdEhlqx+MS5uyAic6/jF361LbDitg96
yMlDpDCh7vmSbqxs2T8ip62UR8EYgWBp1nUK+DlVb1DrYaqrn4MxmgLZcYQ5/rmHI4Yh52JroYcr
rjnuDzkSPUFpFoBnoSSUP66JvTDHXE4qCfjK7R61KY69cB2z8jS6LqXMNIZ271fNDy5pqjRGugfS
N7IZxeVzPThekf/s0ruoGTLWrgGVJ6JMpgNrqt4/tORColJzZ8Ovu5jypAGGyJrnWk25wC87NHAZ
cbo7FuyanGtT4iQkS+Bq/dPEocgoLQrPv6F2Ar6R7shZTKRb+BzFPvno643WSvVTE6szY8ygvh5x
BZpZFymLMuzeOT/KBnA7dY7PrDprkEoH8xuYObLs9/0W2TDVNcnyhQnnPIkOz9lVImG12AowR2LO
ttFfSj8m/mci22T3T0s8RdVILhNiwY/uieCHjBoxlirbBn0KPAFZ5aaAzogh/1sLr3Er4xAXlCRd
l48Vn8VMH3tX27H6MoNSDWigaYfAXwXBQOi7JYHPePapMUGt7VG0KVtNNXjmk1nKzf0pCthLzF1e
dP9G+VSR8OgWhrcQzP58R5cxrBCQrsfzSZe8TeW9ZTFG7lnEkMXdky8KqA5xAADrDXPoP3h7Plfy
z6083HK7spT5AtiL1iPvr0UVC95RjcFyOvKCWwq3Xs0JuTo3QbzvgsTmIc31j5YgP2KB7aKmhRi8
ZcAei9XsR06wAsvI7uBca7jzcKQpjEROWrteECuvxy0OCVlyOmtZzehPlA6Y7afpQD1CCH0XKOyr
6mApvYScPenlfxPW4Id8pgOTf0vz12cx/7epkpg19yERUsQFh+rXASgwWKIRctQOCqr0MvPtFTru
tB7vWbZ0+XNOEIt93Yn/Vh+yXjRBP/kNrjdpVk/zNP7REbRUykXFUMVSRWi8nAIQ7l2w9NhfLI1z
GJkdNk3Vfr8P1aZkmGU1oJCSqdMJ9V7Z8f/Pwx0TCGPWZOIBjYvPl+pDYS8Q5apvLx9YWiOEGX8C
+gy+GLpoed8WnOkLHoLdF0BqskB2xeibhS4jipCSjFcVvAuGdA8SbAUv9RB13VgkKDEcOLmUvRJI
Swv979G2GX5M0YpOLJwau8i3UbCiFLJUZw6O/DJ3qJHLqOYgcdnF5erDgV7j8ENksoC1D7duprZV
dLL3N7g+AlN3+zwo9wRuCstHkWmJrXRAdL1R7fN77GQOoTilmV95S/vrthvvdqBW+fJ2peHJHKnQ
5CVVP1o7zfBWpdxwHuO8CyA24cGshddHhaLye9JgJjGUKfFHtVAjvJ9kC2z4F70xlao8JAZ4j6Wx
y+rbgYJGdQUMPAPWiMty1KgISnPfoCJYHnwK3mmlRHWpoXq+hCHH7NK6kt4pfjN9wEmKY/0Jjv3f
lF5S2vTrIqIayNN92U+4uRxILX/CASRrFH3aBLne+rewgydqRLcepJxYyfK/Y4EqO2zOGzYOaqPE
Uz7vW1J4Isa7MRcpjjTIG5BYZtOl0FS3NVYaklt2BMtdiGpM9O48pPyoiV4NvijQjDXRV6iIZjkh
7VyE6XYQZxrS+6Q/btxixKAQfLZ3XKDhloJJakKearU3rdrcz5HhMaKtDf8Xiiwu0MVLhY9QAUQg
Vtuzxt1MDGL4FKsny8JFQ2IicoX/JyQ+EwTDTNuFzKoM1BqoyMoqya/HAq2qt/wdHvdbq9Ofp5wC
smuNHHU06WaSoA+War02bdZdhomjwQiNzcNWcBauZEhFZF284gW0kD9226YtGHegda5Qo9g8dKU8
KaCos9oZPuaLogiXr9Ufu3i+EwuNDwyKoIUvmr2btJnzvfQGVp6SwBfkV1l5uqM2wfeh0Z69suRh
0dEqF7Ti+w3ePik25xUVFaA1gBptGKsHFk+6SakxA8Qoip/ewGnw0vtbeEAEjeYhW/7AjoETay1z
dhhSh/j/QyqHfm18Eas9in4rm4HfTvxhla8Rq93+6Xt3GIsggsnxi/EWSdX3eqkIomt1YjUfOTqm
K/+Vja2+MSYf139HDZUarrCsv4ju7DTTWYHf4O6/JOdHR0IBwvTrs17/n3ffMK0ImBadR0Nx/mxG
Kq9nWZq3j5AzWRWw0Ro/0lZFCa/UCFMS7B6kNAwR9euumZteZQ53vDaq3RAnJmvRDt3ExOA/MSm2
ZDgUFiibAb7TQr1Lva8lfP4ieQXjIhYyx6wBWx6SGT5hUcZWfPE19eLHVRR81GlOfGsf2PhHsjAh
j4qjaEI1iDYbK0cGMJcpRMLu5/f52U0UQnLJAUTAMya3a/82uMI96YX0QmJ5W7UON7lVUte52BPG
k6/MYPuLpr56d9hy8n9kCb7JU0tiOLVSxTwC8MHBOvUEi1kIBTJmp82WEpCQGgDFYqjLGk6p0kWb
VjOOQCQOhsf3keTbsPOz2utefFylPDLBU6AN/IulsYF2CdUZcVneYKlvl2sGYCwYmVRPYE1zEMQH
85EgGbtNRlGfMIWzHTHs9juUQL4YFYLWnbsuT3z4VmGSsq3In3sQFld8eANIh/JJmVOmccc333p5
OJMc3uiEp2Kb8YKN766TqeSdogHX2Ew09G3EyONGFifXh+D1B3RaZcp1/wc8wEKjSa2SpGV03+DX
XhlipE99ZVSP56dD9S7646eJCKwEQsUoZjfRHvgW5RlfwOQtXsnfe/5VaIm1Tuy9I17eCpomi25l
PCR7SzLhJk+F6CDMtbCjZ5Yy3zbjzj89nx4iuJgVx+1dTIHo7WJTallWG/cLVGfmnJwtkjo1imrC
ussAfOPkRkz8xXRbq3XakEYgT5Ho9YvW3740nnyUHdoLtbAFMb0piY1vCzo7zusqKD2ALMwcvM1E
mBHD/XS9m8X/4r3DqnWi6HPY/qVCtl43HZ3YWXx3hx5NK2yCPBB4RL8DIXvGVmrttdoSVnxFiiwc
pMhRBu8jRxhHdwq1wy5WRwZ+JydoI5hx3b6CVxMDMrdSMa9tm1EhZ+8tPnYeYBPswLBrwD1uPl1S
Lm1IgV8e0z4CKRO2Wjl+WMyEUaZGR+YTu+3puvzq0HzbsZEWSU4omD+H+VPEmuA+g1VC49cBrb3I
ZekG3JU+ICnlGNa7htzkVKzIw+ZAKL05iLPWXlAdwuzaRP+KpfukfWRx5vAD5nRueX+R+7AOBBH3
bizNGqrAW2FMH8ET6gn5p3Zs8rFdCXQZYTuis2vLrYlHXusi8V+1LKJH7cnMzQRE6gp7kIcXYTfN
T3BzkubA62ON7Pms1iT+u5f6i9uXsGDapxTvtoYmb0n0LJbGClqs35tudMDZrrmdZxNpGx+xGOmf
X/um9n6+x1xqhbPmQK7p0jys6YjoPq/GIa9Zd5nMGEZfC4DLb91u5Yvgr8U2/dxC+TVHjcpJ6F3o
pXd7A3Ogik1hEZ0Z7RPfF6OAUjV3c9LxRaIqI3LtIbDi8xpcYeSXK+kSigj7DMmetVfhElbSHNvu
PzxPRt+W/fg0IKxWiaObPxaipvW+IjCdIBAjTKqou2kd60oFjKQ0we0wRHnZUHG70kDumkAmv3Y4
4ba3YBhSnpWFfKonXOs/YeC0WrUaB3f0b74q++n73hGwenAvJU28XpM4fMxIPtN24K6hCgAQakIs
NN9Whpl+oSxBu4EqyZfrmPBUlo2tfNEPc4Vh/Q/vtn/4IUystNbs0SNRKvVV3Q5m0N5LBPBo9JqE
jEMpaZOcade3lSSIUxDToj/F3GMd/mxuwNvPUNxZyCu4QipYsdvyYfTXdURSIUg5rIXBEt3B6hLQ
VlUHxg/POXTTVM4RAPnFnluhtrjsuZ0oOj5tbe+GFNtB7fJGNgfgSYPjQ68xhK3F5ywr7LvmCXKU
Ghfuuws8DbCSAcAoaTx0hdhddVM3qG9JSC75YgESY37d3tmoEWiuAHG6u7+VT2oWyMd7tKAfSo2d
KS09RS1qnfB1vgY0ygBxHpkjgqxA98rvomuu8WhPY25uz40PTCB0mANPR03IHPthzhicYRW44PSU
F1SdGF6PpR608+bm6paj5r0GacsH8v6kCfs6+/SmZXpJwiykxkp4Sm/yJZYA4BV5pO5F+pVnsOSh
puGnzYaNtckSOjcJ4LTEr/dF1N2x0ouGwSqLqZxAmDARtIVz33iQO8/LhN/XHfCPWScdGDTECJl+
Yjr5jlVwOxZ+f6Dfge98MDu5ZCJ53u+C/gS9BJQOPiqeYdscpqH3k/oE+dr5ETOrVW8ItWNuFHHI
Ub/RQb2lBgl2Ox6aj5zxAV9r4tTxbc7CnP5MhwRqLHnTPP1KAVLetwQI3JS/aCE09KNv3O7Vu77t
LYg+793mOolnKFU5bX565iKc0g+ukrvFaopcJgv15y5M8kD/4bJ+wGfiG3dG4GbkQ1jkefUSg9bM
/rd1dtGijuVm6EweCwlDlFxOJh54vgzQvCCF0B5xswByTZ2sKrsF0q7Vh3G4wHzU528oORSkz9hS
y/6yab2Es2Zgk7Ei8s4OWVSnWCXi3yhgKObCYK+BN2R5lvHdEE8p6+ipakLALLwg16IJDx7Rxkrj
/A/jtSDLI2CDtVnY94f3fRt59JfDH8BS+Zpzj+4pfSgFlagoYeTMX5WEMT0y60EtSSKAs+fTLfqb
IwHaKzoqwQK1pf8fbiZ1GVLwCGXM7hUXpyemFeAzKZdVOGqGdbdUGkvmPmSBXnnO5450fAAMPvCT
scvopZ+Ze1/TDmF8qv5/jIDF00uboa6SfsUXThGedtPrtIjrzQQh0xKZKt8Jh70/WHfVf3+33ELZ
Ywfdho/k4eR4Sm0BaDudnoyOsKNZtbvzEDzlt3G5AXwESG3e0RWzosP1eAw+Oofh/781xVPcXOfO
A8La06x4FL/hj3p8SBQlkJ12vbUIZykGXgGKHsHK+1IV48ZLBYcuaFRkJfd7wY0c12FIFygOUqbv
IdXLFe7SyABWfrDGyy+Zbt6PM7eZ6h4uyIkCkUGCfGzN2siz4DkKF5sSbdXdfSWJcfq1IS6um3ph
moSFwQvXtIg5Gg/olM7zzGI1pj1Mj94LFguYLOJrXJD2J+RgK2tqj9GSordCbJdoGYvEekQy3CXJ
3/HxH8UngPIRIoZJUBTNZkbnBeHHoYEdFSiwJ6dV1yyQp+H8Mpzbh2wV8d6A9eYjfSTKwo/vfm1l
DwPQg+mmOeKp/P7tjURdGvzvjOwjXsIONBikaQCnP/3n3dRbR4/bL9YfjDEN8xUL7wVOv2DF/drh
QL2ewu/L+Xze8n5GylmFwRhsArU6i8MgZunwtB7B3S9bN6jzQ+eyIasqA8ZAYMUVHWq98PsjyxC0
cKy28/EaqoHsZ+6LRlVdxERynL20fKBVQLOPMg9VqmzLXJfgo/BrRpeymlD79KLQyOEWAkBYSQCJ
Uv05fIRNc8Krk7Z2YoId3fBPtIJJiVetD1G1fLyTILKfeX6FYxUMHR4tO+2UvnsDwRXmlvZ/aY44
VZeUBCCEN5FCEPHRtjVP86sLAkISCWwopt5Og7l2rxYWkmiZjQYBkvynHK/l9KMiy2XZSQvOUPoi
0KguNzOUE9YTgK+QW7G/Mx/AypdHtYM0Id6iVvWMLVgNawDvmVufU6tJwfgsczgrzkfAKQueZW+q
TNgw7CjteIR88mvIuMwBw1uUNMFgUV+tms0ogT5E03/w0fJnpWHYRtvSyaisL1yOug6Wv0jnmLk9
ZiIeR4goGUI8pL6A9ngBx8nsiSaX4PGa3/6JoPZcb2V1+8OZ1hCiNpzE51/2gutoGp9t+scBhPxF
/PfYgLyq85Uc7ym5HA1Z1XkWnJ8Hksx5dbqezXwBOZbL7AHIUg1ZFlk2i3kZ/GOoKeKKIh+6Covi
fHz4kDWFXy5NlIo0OGnmjIy/fPuaTohFRIZ1sVIilnY9LIjofCatIdBO/Jz2Y/HvCUGIwuUjkDXw
9gep68bxJ5p3qs5VjzisMApnEaqoNl6fc3zECBXaPD6Zp7LUeG5YjNjm18QDFSAQ/drILGgK2sAF
bRLJJsDzaxH+t88qcPBZ+P5gJfnRKJg+09OkluoNBZy2yhruUlVua2EBnyB+g0nKaYHehO80YD8Q
Ntgi+Yct67lpYktrc1ZlxMaB4Q8fGY6SZCJbqUglCbaUtThD/AWjNOwOY/VI4PLG4Ii+nJheHrEF
iCUg75kwSvpr/Ay2ZO2kLNCZ7LJdSnih63LDfs775Smu53QIYO5Q39ZK1ga6bvQMaxxqfbJp/U30
QQ6srT/DZwajhZWkE1kiVf6DDfmFmzWfdkzWkcKJY8Vp0V1OSYgmDlEKga+pXNuwNCosNFqwFOqq
dMMZps9dkI5umCKtf8jNXBYNDg4LL1BdjqmQkbizW6C+RnWLmPKPYPD6kT0qqzpPN6jhadbcNaKh
khTQClXNzrJHjs/KG9lRtY1gw5Top88OupJtu5QgXr1jpHaVDZb+WZuLArlyFarz7rz7XxSlqaGr
NKoClcSfRIIsOSd1pHtXMZ+G6OBnUMGOre8noJG1rSqpsvf7tnsL7aSMtg2sTgHFRtHPvmdBOp7i
BuqM4TttoJcZB+sERvvPuOHAebq84cvymCDe6HgzXEBRpoXMorxzL4XYtcUXJ9A9OqU78TUB/glZ
n67DWQnvUdWjQdQhHuenFkrDmi/mA2qZV6NUf9DsnWyZdnMLoq+CCBiSjAVoW/uN6vLJZ9Xg5jLo
UgTA8X2Gyni/TiO4hrTQ/T5ymchoP5O/qF00IL9DXDO4aYTqJQlafrrT+3HXKB1BbtBfH6TS81D8
Qc7afnh3gktFu9a25Gh4TN/FVf7PQ2ZgmRTVx2oEblV7hw7omjvIDSpsOaNBIYxKJoUS9n9bOngl
XgGPWlpZfgnKex+bgkAFymn4wLRo0p+JNTDtY5mUPb/RjNCmBbjyqDE7ngMl5riy6DVJuzOB0J0F
f5lmNbXYDSr6zBPXBi9OqDWFYLeGAWFwl0exISjKTIoDajbW2YadO1zdSnsUuHqnuNjQuI2vT5F3
ESu9c4nBWkr33h6Fsp9huQTeH34lcMKDwUtAcMTp1k2WeAIYZJBl7zo8M2+TyRw7zNPtco3d6BKw
a386AhAK/jJnmB0dRrm5/dptWhvHwHu4ud+XILoVd+pon0Ta6dQTeDDzkWlyz7JtxfRItad7K1u+
z3fuuBVpyKx8EexywNgKtBTX6mjEWSrnbei8PFj0lSrqWTQKlgnYYWvoFjKR/r+IsGUWRt2sRuln
t5aK9fPr3ZfiRa3aMIwvHSsYWgUI9LXSNUiuG+lp7Rq22Xg9e9OPDP0rYwvF8UmbbLNcQj16tjBn
RMMMSWGSuveNKeySy6vx3zdHStjzDQiGr8DI/mQBYs3eTHsryyd2BjPqi3twF54ileSXOH3+6/S0
tvokgOmTv7MtOzfmEb+Ldt5HprRzwcEIXPz0UbtClOcBB5wjwCNmgT/D9rr7ahZRC7l/P0POt5PI
8jW9eWWj6+ca3Fj3vH7nIm+7xotouqzM/jEmdSrTthLsX77TvTE9kqKMlO/eqp1R1KpiHcOKC/B3
p93/99oi/knj2nDLgFVRoExAIQDfy4zVUyaNa941Yepye8mlhleIc3rSSbo+ctvDIgT93D4jPt6f
bDjy8+XZPartbKxeNMDNJlE06oJjygRyVPRdT/DoXzMGGI8lthrbPXoCA/rXuKyYuxXiUb1I65Lc
WGnUHtgRH2Ssg3FZgq0NjPTuOoF/oej28uRZFR29gIQB/3budHcyR5OpIpWXp89MRa5RscFXUG8X
P2G+G1zpS4hZv5Ya0U+ZMmv2j2573XMV+raavtzUBvT9ulL82T6kMIMlKgdRy2CWezDL/3vZbUnF
LgWjIc0bac8wJylMEAePrjeDOkEBsklu3q0tw6KtTTBWcWAWe8cuR9OsfeuWgp4wMZss3AuugfyM
tlPWVhFvuZR031c2J2pdHyBGNi6ns5a7/IpliP/VQXNbne3aKXnRo38qVnXeNce/GifGoqF9Ggkz
A97gV7lypkk5IS4ymmz6AVjQZImuNGJl5CtZt8mhDK6rcD5uiZDUpZvTvq3FIhHRsy7iQP64qspz
lwgSmI95he8CUlkLTGC2jSiWATLkxSU+Ne/3vrHjSM3bNNuQvcralVJzkiH9KzsMVCL8WpFGVdxi
ygDtcQCQpRFrl2LF04EcFfADXdK/w2mribNJfDbe6cNSN+qMAEBIT07grmI0qOUTCXr8nAv1e2Hp
ADZuojujAbQaOv82MXYGF12cWpa8Yg5+9FY2WlQN3T684U2GvjzR7GDUUYN7PAAekJYfDwhTWtea
5Z2iXsgG+yBsWNF0z7jqE3w3jYxg7Monmh9XNkfLJLV8D0lrrvq6He9qDcrA4ls9+qYDMTAtyxla
Ihg4aco/+2XKounSeSgvPxoePrpwcfTT2alktFqA0//htm/W8hnQc9/bAfbeqznIKF6L/0mXRPi5
W/cJLvlxPIyOs1PrN+xEnRwEeo+vX+oqVtsPH33nxN+hqf6xif28ZGAH8o7MehPL5WeMXTD7XgqO
j9EDmX2xj0TUJl7Vv5uhgCGqxzI3RpxBytiW6HxOEQN3OCvXma61cZ2iLlTB3VK5IvWoCzL1IZV6
5X7to7I4sjxDiY1zKlYyUvYj08W/k+5/pEAdBjU0QbzTN/+GjAzNBM8nc59DfGF7G9JKA2dx3fdA
QwKOUEWVj36Kj3phaYLorfPFIHKHHrAtGBeeexU4U0Q7+LOLoNSUfZ8+niCowApTynyTQYs3wpaK
AwlL6QIljXjPLO37HeHs+QLIMEN85IG/jBpfU2g70PVJLB4vsvG/eTJDjkYZJLVZicD6XaJ51S38
JobEz5a4iMAOq242RLM5/OLnGh/Z+CauAOHplyQ/XcjhKLac+CVtY0PqAx7yuSKLfSTRwG5AOKrG
bhSis8diSlYw5BTr0hvJF0lC9Sr3Mv2sYlu7P8NstMpAJHN679NxL5xgDvqerMrbhRAJmZJcm2lm
4wOmDKvInQTBVwi0byfcvfOI13omyYe9dOUkJNui8vAmbiGX67JgpPJLdLGmPZI+HFInf9c/Kcjx
+v18OvrgCjfle50U9APCRbVqdwJ93qJOHk+8SjkEN8J8J4hlNEDQ2MfK4YY4bQn9JxWENvnnt66i
JvPGkthjgyB9Lhf2tML64uqUVAOMBKDoF70Yj0kY66CTgcPNB4aBkZrhUTt5RaNN+0W3YiOBhBAP
R1jtDc2qPl+Pte0Czp1K8p8hclgH5666spzFRJNyPufwv9L7E5DpdtJ0KomLYCzz9AwkoxCyiyvS
cW4HZfZNT0PnPJbxH0D/+eD6gNoAb2KTAtBPKMGnsZt3XDMzCFTTordZiqndZkbeKeNMxlzoyqVy
aP7qdX01Ye5+1RA1ySyK/sBDuW+9w4ye/Hfu62bqdakY/GME/wRBO2qleCa+LGLhc0iyCZxuvCC0
GgGVART3pImVvA3Z229SIqlSNLeNZwzBquKNCA0H9Juztbbc8h7PxlEMRwABuXdiCUr4xmYjchyM
G7bgfut2/aQLRiVmbTa5p28pEYyOiNOboodmuI+f79VafbtPlTg6wmEexGlHTpOej8RbDd2fZQBa
+cJhPeV/nteioopyZggzaIonPKEpQpzYFuhAl2YB4dKoMaZGJ7Mm8f3t9+DrexWZ0t2Rc3zkUmL7
84baIW6xtHipg97ateUoN5oQCCA3T25+2JlzSZiJDPBshTIGbfrKquh0Nd/Q7T30Z7ZtyMyQYqUk
APpCzo9kqwce1IpQW6dtkRnxGqvUhkKGqHYbOMcjwzaajptTJEpjJctKorLNTKGsUYsv3eoyHpjU
na4FRkYyPDQ0z0lOpUrbjVypzCYlXGC8vsatI3zIqBl4Gb5+DbkXIOlNbjqzoIWMu42EVYGWWAKL
F9+tX2T8DFMGqTrD6qP88si4Ap+T8NfPOw4TRDYJuLSEvjvfyzjwddOzgDhuTVuyk+3TZz/kP29m
S6avWKyRP7QfsoN/Q9N9ryqSWJEiOfgCRfZNRTPjeCocr9kbeEvw8X2iMYYN7u6W9joO2Plndm46
ZYX8kl/03mRmmraeMkKCd7FUQne1HQhlC/K3h6qzZy8xA+nlQPXF5uN6i5+CGUGrjJhy+QLJUc6Q
LgSSDJh2jSdvyi/92sP6ZoZRUUzvdYHD0bPrK3LBeE+rywuGCLgakwJTLfNqxlZpIujS7fCiDGsf
X01QASPQb+3A/H3OHPNAqU0pWVQVXGsoENipUEaPPWnhcS5utHLkbMtb3aXTVsyTp0v9n+j2RV+g
XdSTB0m8c3X64k3Bqqtd+GEqp/uTAr7AMlIczW+++ERDP4Ew8eE85cdcoehKgxxCVR50kmMccvTE
TMUEG482aqA/Nc93dczyf7yVr97fsd0PN4xtuSBUGJRyRrsCxKuJH5LnzdSSOU6d7pIiOFR9o6UJ
Pafrx8JfwNXRmqBvhDQ44cfDUepFZY/Qecys4ee3loAFwzueFUFLehMC5tFbknaibGj3jCPNBibX
+2novIjwC+GME0ycN02U5RSJXf9uKOQWrCnAacCVnmjtGSTt1rbfl3T33SiWlnadE8FfHeo2GtNv
KrXqAcq2n6i0PdbDQs5A1XtpmPUHGSTH5ZCRNJpltFSZwSWOEtLHJgeS3J40i9HUWG1Xme+vtscC
kdWeeZbTYWVeXgqn4d9CSydjT9L3Sm79gF4vErIJclT+I71S0TftGak2xNw/GSgIsDOfXEc/KvSr
alVNCnhsXhqehsUmgGfPD8HkwgNi49NX1ckrTGZJyjL/V0Bw3dA3vPs4jPM93oEgCYhQ4dGueQ1+
B3KJHWTm2JvlHHzssxtuWDzfQp9NrhyvNXvmc+Z49BpdAo9fHwFKVQRTp3bdeTwAC2iDi2Sm6GIg
vKlE79fZn2VhbaL93CfbCAgbEdgH7xrQpuQJGqDPOEJIwwwXVjKSjUwNf4cqqnrrKBX0mJyWkuB7
KiyGqkrSVxzmLDPzlgXBr1AfVkXGYeZ5uPDeTJzskbDopQW9dt9nklFgQAxcnepPJjIboZuvaFig
JfvK9wfwsi0WcmBtqKPa+F8BilZ2XkzOl7oCgGlDgEDc2vxlDzmrZlR5LI25nU6kzfS/a8RiHi91
Y58bg3DGMD+zyrFTvMctNJ9jb7eLg9hqyHNb1ZQ4yGrb1llYSJOBK4Fcv13pcPVGFZlq4SDq2GGO
nUk61lAuDFzxKFwTC0RgcNx1Oo4wNSy1+vB+5J2y820NRZRbvVmSytUnvrBcIMvQ1ab5ofUt412U
ch8z9JVvAIA5WUXFWJLT/moUjEMXztn0mqtaQFUHKbXOVejnhEJYxKr0VfuNtgBO7mVCEzWhJ1HO
xFtJ7cdQJ8HW+OvzXlv5sLjC341gqoMlaHQjcEiWRgFvN/qxWytyolgOTEHiV8NDbTt6mNNjliG+
45c99xMbaFfm4HgtTE8A3z+BVY34j8J5ERzzVFvugJVyLTRTuBS4kZb2ItGRIziYUQEQhF2rcy5f
bN0HIGoOZMPxMb6I4vIdascr2PtvbBmdpCzaStY2QI+q9kYHDgo12pBmDght6dS/IDac8AnfjQcF
eXMY4ninqXderH2CSDCCmneTO9rveLm+f5R1a1LZsxgKgID+mXUj+vWflq4Abn0BafV9Cf4mXfJ/
24i2wn5hfIxJst1gyWnyG4bDlUZLQhhyodD/j6tWVfgzGoKUwKhrQWJ4gVp2nrm3WiBJROJSYiig
ASJJPBVRuNUVueFewWKat1aBqO0gOU8C8dW05uVukWkw8H/unWOhP/qV2S6YmBcKSI7iOfNpwLCM
F/YCjrjKHHiFd2tUk+o7bca5A3QpcNFgrXNLbYIXecN4K1h7kYekaSWIzf6OqDJ6m0BRIX4PZWrZ
xYAXBJiP0yIgoPnADIqGntl1kHgbhfFMZ+TJwggVxy4XYcdPnhWMkSb5MPBpCfUxBdxsoBCbPLe1
2CLDb+9TaKbqVo4FOrCXw10Nts+Wfr02zxfG5EIKVpxjbyd5/XVVuzR6p/AK7H0AQ1jMQu4zv5Jh
X1xltz7zearjRxl0g841I42N49oB32QMlIlix9gCsx0hXyxR52gsDD6Yp/pn0TgsMe8L8Re0fXMI
EjgzJUru4lzQe+Ibycduosf+0s4TsuUrkg84Rt/ZzQZKt+Wb/9rPIGGiBFuWDitXPY0tj8gPOAQ9
dTnR6qCgb06xnFaJXjrFNwn1KcS/7RMxHM9R5Q3TWrkPMPXUH5QCtsf2IzJM8U2B+kCDL9j+EDy7
6SIbIi3w1N86fwjjsk8hHHjHEHE/DrxooAUL2iUoP2ROdZYLlVy9oJEuOxrRPlQJ02mUs5Xwjo+y
I8Emo1qkuY4vAJ9xkaH760Ii6KDNGz26wfXqp8GJnMOgeAvcNylprPJKX5JEwFa0Y9llwkI4canm
HXN+1fA2JF0j3mQYY5P+Vz3Vh6QMxc3B9wTTkR5wgXwLdVTf3+67HwTCqN0l0eWpuVGkXFftIz28
6m7ZxqytAy7xZJhEIjG6qi/pY9dkyGBj1bfU3mlUX+sz0+OBQU15NaDs6WAnqenckmnw6WEKU0v5
cbCvbM9nvhXSJShVAfaILgw+p/KpNrBbYeMe/BbMjZPspxmpYCIL0yILUNdnH3mww6b4CzH8gHIq
kyPykJFSt39DhMNOJ31ODtu9nCokl7icoeGJGS/fAW0pJeDcXAsPyFpKWMO7nDHeTPz+7bjEMHNL
cImGftIx75IKp/UmEufi3Vrf6Bb7Q9cdurHsM7UTSdWydDf+KKuFF4Gi7GNLsgb/Rj36zj82TMVw
0js+thYQdGIh2LipzPHP+g435xBumyDBBzOevwvJbZYeO+I4ywTULxXGBo8AoMt2EoaRd2PPaKDB
ysLkMkHN3ww+grfUuoVpfXRdSlZYFgwm6hT2NzEGKBI3nVQYYUQ8OLWo26DOjQTsLmVyR+5JxZQP
DqRO434AXWDpP4/TFWh5frt0vuNdb3vVIS7aaIkpk0XPan2nkF6uuV6MtCppWSxfS0NoIJIPN1+E
+fwDch1RdaqKwzchkQvjBWpsaNGpqO05BMAsJGYST2BOwlS8TfENJNWoHh3/Ar4YIKELRl8DPPTF
P65nmpLlzHM+HULDGwdswGDce/9qh7sTzhUn1bMfdrg5E3gJL53cXZz0LZx2VS8DAyYDFLlgtrKj
n/y0nTPfNw/p8EsEUXCAz5sETM93RwD4W8yHtDoAMdb3HVUfBhroHRxovAAY+7xZQMgtP36K5jbT
ipOQ+NEhxRvM0K/TbogMpv/66MSnyYFBCvnQTTKT2fe0lciZ8IXGHnbAn6KqgUETRRL8o6L9KzPV
6yuDo7LrEaEazSAoqi9BLk5uyv3P0QSjDsNALrnqQ/PI7oo8Q/C/L+iZ7eN6fweXLlB0agbq1lZA
MT58qq5tjA6tJ9VVGx8H/rr7q0f2kGYzzF5FxQUFQAYur5WVtKasfOSbYzCI7UhntlIeOfgYik6H
A3OgmZV/eFB8K4rJUd/TjrLdMkdYh3v0eIzBEGCBXrY9/7X13Cqxm559fhSG7CLrKC9HzhOWtY5K
5FqACE1XPKy3Wl6IOMT+HQg0iZPHv1BYwjyZiROHiG1zffD8bMJiBrOCUW2ySMD2TAmu3+00GbdD
jEdPAkxieOUDEExQEaKr44cKlDZLcRwHCAEuObRq4nDywUVZpcpuAPNDVKtXlKaSn1ZGlPcnFuaU
230TPPHN111pNowyLk1kElOYhKP0u3/fX6tP1tRVpAey2mx9WSYmAjP7k98sytFDTRKVQ/MIR66A
9l3CaJniVjPhbsuU4vJ2R4donK7ww3Oa8G9IRjA6OWB6j4YaG9OmXdf0tgYYav8D3763LjVZo5PN
JL3EljH5QwGehaYPgF+l4W8NRMlVW3Icxq7xCuhcckBJbEwbbXTfhurKxF3DZTEQjXz1it/gRcWF
J58gEdv+g1LnhtPqT6taFUo4M1P/qO+JIlmDyW8uV6iXfu9q+AKY7LQ10ndy8UD68J4Q0+WAficu
P58Xx7B1q72WlA1KgHVTMhUlZfsrW+bup549LRWSAPXE0fVKSUMiO6WWWNZMIVyKtzGJlso+DLqQ
0QSpSaQGDMY3Cm25/XZskyF3bgeSlVbcnDx/oYuHfJJVAPu3ehIZ5iZOYemqyvOP05Bl6hmfew5l
V5RpDsar5i5gLg4qcomHz5PqMhk0DDfXtsGo/jCSsp941s496BiDw077WSPLqjoHFwtp35mosG9L
DB5AoSpIhPPzz297Rurg7X2igx00a1GuNw8P6r6fLVUrZcQK/YGlpReujybHB/TltbxjVGsxC4Lt
DbcGRvVlu/lE5xRmqQsh0MuB4vsXrkc59DlFhDuwdLOETxpQYXyZFwTabTwFV7vTbapfD9j/iUaP
8ApEQcYSTWxMeS9gpKjdmkD0uEHsA30liGvPEia5uji8cG/z2TrJqSKXkbCgtt7wfBFADA+bDE9D
DDuguZ1yN+TlL1Bq6OkLAi2m64X6z1cvbixis7BQMPHk5xO7bgCgsrve1diCC5casDRhg03h0dON
tUq3lDojpSbOLIxee5kS4rB8ZhYNf3EIbgeegRAcsPJ0IQUdIE+mjqsFLHcA76FYTEaQnN05YY/0
BtBsO30Hz4ODa9sQC+YK29Poppr0U5hmuDZyricx8ShaPYFNvMZnoCdEmPVLLqdvcvmKfa7CFGqT
1zO0ThFrdkh447EuxPO1TWNB8wNs60j0PRkxwiFm1ZqOGGK752wvnTPP9FOssaoFWHWjzM6mLtyi
QB4Sq2eQTOQb801n1hgd3LCzrf/HDnDgmXXnZj2wV1LEnUf7pN4iC0XNYSnkjMMaRQCZ9kztrFE5
zAlDF4SvtWFnS5OIPgL7Zgo3PmHZk2PMxdBDEfT/0WkBFgZ7G8GQ75tAdkyX3TiT9jGLtlfvwp7u
DKnTcBDKeu1uQL9bfsyx30vq7nmvIKxiw1jwhboixIX6O7JwugM7jIAd8NuRWsKiSJ6zpOeR7MQf
gpqiQm9I7msszn9a4m+6xF/Dv02T7QzQ6irXz3xzRippFuvFV1ovysLJD6l/Np8bM3Zf32ABIhy/
BPFJ2GUDNx4JFq6wfg3CNh65o8LDSi/gNo36QnIBAjPLkumyWfuYNqIev7lld8pNgzobd+IqZ7+S
pLecz1cBFQluBuLI6NxEFNwcP6ZlFbRsGnz4BvfK+6YcF9IEFKF7F94PgufUn8I9ByrT4xjvNNrF
LzA9bpaaeEMmW2fFcUOLCHeDH3hIB5XaPby+Rv2WB/fZnVrbvNkOaCdMZPU/xng70IoVF1tRQNQD
BzKoNHKl48yzdZ5bmYUvD2tYWCdFAkLmaXxA1Jf2cqcWT+lIKipaq+ZucfsH8YvsaunAKfW6qwlT
7Jn873WsS2LgZTwHVg8mJ/nUCtx+hrlxuTkVSMXsm6/dOiw+VlEkms5jPtuAqUVEF0R8tol8DkkF
UjgIcu+6H1L6+f8J5J3F5YsYHbACdQs9m8pR73cSFmzKG/yzK/7WgoTdRpWmMlc+k/7sEJJheBlu
x4XVvgnIIBmMnuESeECh1cGJ7thnC26slOvv+9Dq+UsilpXXv6duw0deO0NfB/JmGiE+CRodtUwg
6KfhOqGVAQcAA6dyyDtGLn5P49k3aXBx84J+OVXKJbZAEipv/h7ieT/KFloZdy4k3K6lVx6dRJqr
U18EIB9rYEGbq5Tr1Uexwz2KzemaNwc/c6DbTYqFC2iSySTrFHpt0alD7EOZ7JEeC+LI3l2x/UbA
bVwXo7K/vy/ImE4PNlKApuAQ2BmsCLKAHvgOc+8jX0jrlmH9rhYE4jEdx+ZPrIb3zxk+Cyia8D/V
UR+SHAJBPDCF9x5uCCrezaaUveOVS72Otgph72ab95pvtT22yAOVd6FOCtxCtfqZVHWYtNsibj/l
THjXRtVqgWr/tdxrFfW9Pz2ZvhpmoFk8bX9zG5S2uB0uBktq3m238cnxcHuryKy1FLu+B/xis05c
8K3sVbGMWPx7xNjY+xs9qrtdpdU7di3oUtsT53hvvkJ8KKHGdoa+Gpdl2AjGU3mvK3NWE+S0TwXf
WqlHJHV/Vki40L6AGxrwVQY4F3Z8Z2itoOZruW8SsFWppI9mYh/XNZlASIPyl2l7Ltzh9e4Yr/26
JuXDp/jnzTjcDtbl6Msl0FljF3ro4SfjyIGNJZ4VfWY0ZnkAtTu9OeB/PbwoD9PCTbJ+y3L5Y0HI
DTXcodoioxtoJeWkVnCoM0WveExG5yZRtpWQj6OqItmLPjaZVOr/waC/UVWZ33mCBO7Nr9RRvYtY
2Eh31zXLQTRMEtDXh+nUq+sMdWXB0ivMQjIt0Fav5RRK4v3B6HhxY/6DAMbljvmSifWE8Dtg/Kbr
CivRx1npeb08/zC3v1IePrKkFuB0osUrgUlr9ejLhajzpBgO67Wx8OpsjQMDaTD3iNX+jsP1inHI
DIQ4MyXQydSu9fmLWnkr755irhPMHOnP+EEEp/Bja28U2UQF4X0XooawWyJ1qAt+xJiOr9SvdibE
+G5vIEGuzjjcb9UhMT/G+ScgLNA7vMtj//RyJeiGit4XMaArjnMp06AcFA4qTQAwB2BcrNfPxnqU
KMhrg3odIkG5oY1Gooh7mgOgw4ab34ujHVJk583qHr4b1KteSjOA67gV+N3z6uV0znYQZ2TQc5mQ
09lyEvfe/sYHLrx+U5S8gA58+QbEoK5uMLYfNc16GEHwXBfZJnCzS3C0jab8XN2ejCWaDUOPjwP2
Bc12h4oJ7vsmnnXqlrSuaRyjUPllmeWLklJMxpARTQOTxmcXANu988uJql5KAxy3h4Zv141tdI59
2zB4NmrBQey3i663a0K2gAwhha+kymkxWPcDGxkoNg05FxYu9LXeRfZe2uxd3EWKz3DyarAT76iH
vQ+NLDMXhi8WLuR/O+6ZsMn/yMZrkEQ6jGd9tDlaqvUFk2tC4cOyHP3MjmY+VyKSvz7+03Ug1Wrz
bBCwaz1HvCKXrFMOLu4nOqa5hb/JkD5t3pDhdnx7W1CXcTNW5vIWE27hwttweJZkMcIWrdySUIhA
sBF5+NR7RSK05zrzCK/oUqWAdaZhQ1ykLQZ9QDQt+J/rmRLqeqlYctt4h+aE1gEoSTqDAATpWRA/
m0FEE8KRFs7x1mZTjiamgRU0JjYnpgh3LHAAdf7Vl5TfJiJERWwJm+H2GUt+Y6lnVly7mda5W2+9
z5/X3vb10el/d+URIki3THpQ2MhsXpt8IpwG1TgPeE15x9WkaDS5XkIvX3mMjhtQB2DQIShO5rvD
IG6aIYeRm6cY39tH8K5Ah7JyBRbXbUHrRHDeDx1xAkS6RfJBbLuwr773bvFwJC6wxISsALNOMhHP
iOCR78yACF66l20zgLpvkW6Gq62vyZAyyKX2B1iKixi0JgZ0M9bOUjUp4OTKLmW68fyF7klgnJUs
hagDd2vi2TJJ32FybqIuLhpoaErl8GHKbHQO32cw0SVcoTNwVFwIzVaWBnjfdSIMH2VkhUi191dD
tUMZCQzxSsBFoaRXeR+mtCZh3jwPfpBCN6mpEvp8WaY/KjQb40WCcOayuxB2JJQv1sSQMWpf4oot
uifc8WqGeTq4yKf9gVmtxmDQCZzrUhJffaG3Vaeo0FQdiXQiGm9mAZSmS/Vdk6jxHV/xtyMQVHfr
fhbaryGfaFmG2EOCtHfpOJjya1vjJ8r6rxFigs/zRPr/YvMhJWCIEUkDG5FkgJQCIGl9pCFT4mNX
AwnhgqplL/y9ZLBY8vJO9XYpGGXtjaq6hLTpq8TPLQZhxJCZioU+Yk0rNVqzNHA57ModwivR1b01
QMg1z6PcI3zj5AzDRAHC48yXO/jB1JXKJsCHSZS1VNw4B3G6Kks1thzYta9X8g8g52VVi/0Swykm
K+dHT0vERLSNKYjOrd3DzZ6L2NW4/JRMUre2E0yKPk0l7T3dxHBFFe7MEj5HTY4xiZUhozC7Olih
YGiC9nVghqJb3EmBNkgVN5sTwjrAUEY3+CIw066sKsYQ/skMRIQwVc8hqNPGajylHrHI4DL6UkTT
pLEc6zj9z8ztKF3xqW1m2LMnNdpnT3W/b9tNjuczec7t7frgULhWZzcpg0EIvzjqmVOdjhtP7IDk
UoxPCrah68pAsEH/X+ylfVkaWoyY+qFpdY8k+If6aI5G62RUGqt8Kw5sjVsYpk+e2Nz1Y6vgqicd
dmXqb1ZYz1j/mweK6hZZRapAmN/ZsJJGDO/gOlqsRWY/vjKOUukX4cihldQrXbY3nxkMHscp7Cfz
W9gttZOK0f9jZjAt9cNQfKDHqjiAPdV0Y9tLHg1eCXrF2FxgCAVnWRA5Us7Ma7g2pJRgjVaDQGzr
AE2i7/PWnB5q//ADPdCGRc2HSBsci0Ly4Jq9rc0IBedOb78bjhgXsYu4AagvfB+Io6qIja10f1RM
ZrpGCkCsw5zG12NDC8VXFZDXczmlM0G4E+BMxMSYmSmB4/L6WdVLl86HICv/e0r8RQt4csQs0PdR
JuLJ+tUsY0fGbZwZQiBitReVuqRrnp9jKc6CvhzN2+2jSt1Mj/Xsly5FfJKQF5RzuP9fmUNzhK/H
/FZaZ/g27wdvQ/sWQHUcQdFmUpMnc9kreLBJkSeYN2FaE3JYq33HtVFecyMQN9R9d6Q7h7uHMXs/
ZKDMVrlwlb9HRCghJ/UixyZe0mxbGOlpDxt7LkofPC9LRkWZDiMnzQvyCSV/cGOk/rIUP3B6pKuS
RpWYrzzlvcf2Q9qIaEqELT7b7Y7D4EHUXd/R32Cpmn2Kv5XIMsURH+LQJmEkpkQ06hbTOGPzD66c
VUA9CePUC9pqB9f6GJSurC/BJ2/M7Gb6sfWSyvigDVT1MFMKSP2L57wDWSqGUWpc5LQE7x/hmYjg
n03mm3vdAoW0+MlhgKQLeZEkg2POUFFJjpV6/yer7PT7VZWEwqrVir2boWGWwUuTRjFVzkg+3+8b
TR1hN4lXnPw5eWSejWqiHv9qxaGP8wXNbOc90rTQQOCdy8LzI7DrEAT+uv8ASZYsnaLXxRlqjiA7
CGU+LLvfMULs3dLpyyULX79+sB63/G1ObpxNN+CLTEDzeWQrGdR+bJqo0zYLBqGGBE1j3Nl4msKf
wkXDSZuJxn1EBDfJ7EEWN2yeGAhakiWLZ76QZJ9ssKlBlMzqtMBnulrjJEIlkOQ95krW19I1ktG6
iN0DHnTCrNHGmWmsNGi4XA8vDqZfgsW19FeNKEw00k4HAtJPuL+osAoKVfdN0RaiIP2WxVhVTK+y
JWcYZmPUDZHMm+NqFFBkTAUeKmjPI8dLCt5UbPU7HRR9v+EKXVsuy49mbPXHKih8t3Dyy+iyUKdj
SF3M6UPaUL8oZl1qxeSN29a6UgdmR+tMspxtL1hm+iuC/UkAv6ipIDr3vdq2oBLbCqKDiLuaTBBF
8pqJ3VixHktyo4lHLKj+zvr5YhkjY6qpMJLpdrminqIFkfkY/MR6xUP0HSasi81z6fAgvAXVsfAx
Yg7hdldw2lDavFc8V4Xps1TGYZO7AenjWvp1zeg7wkE/efwJJ7zdPvTsINhc0QoPBEwUe9V8tlOS
GPfZY6ptBgm77pIPYXHEUR5Kc76X/ETAcc+rcdCyI4l0X2c5ayrQM+EyxKftmqFS29ChAY1fCJBA
rZtLSteyluqq2mvXhGrUPk6T2S+PHzde+97+Pzwv8hEz25LxwT7rz6LI86rtcRSSGBuZl6IdiuPy
2p63o7DicHnIMP2J3rNA3CkLlktdQnBpCitIXy54FJRObo2lV0MZe3zZq4k2yC5X4VTe1QAiJkkn
9ApPElm75anNxR9tMZm6HkbcEczLYZIWr6y64pUmDLj5JDE4lhdDviWdaHMOZKdMY8UCZerzT9z2
lWX30xJCMa1yyMbacwP5T5uUX4Q4RD34rWdb5ylgE3KVQr/D7Ui1p86tiW6kgjAdJRPnvjuDpJbk
JUUJMX9swjYQaJ0FCXQzh6GQgb51Cl1vdjgTDrFlbzRN2kkBfhIbLK4uzrbv4bDfS9mbmdjTAyrt
jTtvueNQdKUScMQz5UsIpQTbI0gQ9QbnTix3XiRr3Kla0BrKPvFVhWyrYmPaR2SvwAkDJwDChGoQ
cGND/9o65qZekdaHYORu6gCi/5ysRshCDI0/YAXAdE4U18JtMhqfGp6uveg0Yc6JNXxA0XeKXPfE
MaZtaq63Meva4QKSFwwLsEXZ6ywarRaWIG2mqVW4X27YrejyikfSTwuO9yscSIUdbcKZfiPf2aRi
8U8//0OMjuL44nGbvIZfd6CXcTc0w0wz6zRiMpx1wB3Lt/Y5qiLlN1bSw3NWQTYL3JqkiMGkbyI7
rM/vmHMwVg+GquRU9EqxCTRRMSrhrQpZCzu2li1z6YtV7s7OihfC7dFLuhSIRruz3HxKfaDJWXiJ
Rmq4eZU4iW2RZaJLnN89XvWhr7rnduL0xp4qYJV9M0b/ONS+XRW546DRbxcw0ag+YiZqYWp357Zh
7BndLwvyOdunZhWK+vU8BsFcPqwnOsmYJYZ7eTKJrYorBx1Le+V2mPFPW4a9rgYp3/0sCSIgiJGV
RwBoRBzjTdkBmM+9OS/1obMXDI0V8Euqs8Xrn/UzmsiMaAN7v6dF/xj2So8FN7QiSQHtOwcEHgvW
MlHOnQrlHemEgC2E9cNmlFa1m3NTOfRtThd7uhPpbe9rTJC/bVB5vwXUPOCg5QTL4l1IJj17/Q/M
COjr1g647uPT+Fm4lMkMjty1ASKZDbRGtrnobA0z8e6CMFWYsZzoNRpg5QbujwJnvFV2AMXnHkc8
9hdHM6srn5+3HWFHzfvBOsZoz7m1Pzwv2MIGUfyqd8EeIjA50VDdRpA22GJkFdwEsMVAKGxMArYd
6q4BhwnowQs13tVqCMEVoBvUL/2O8uBLpgUx3TR34I1FII2e/Bi1xdNQweolyS0c41Hlc10+BYE7
wQUmYBJVkJHJH8icWUeXry87IAYiFWSofW38Nj/cbwqCY9IeaqKB1SWjZM1LFFovanvz9977hsiA
vw5FZgOQBBdUKxDr4aDPevyzFxOwRyhQNfbTgzRYAHrnv+HZLfz8uwq9paSzeBaIM3Ugx5O7/c4o
+xGhqD5YIxCtY4MiJSlW1ElIag4Be/cU8epFY36NdFBZiepSac7RPDTV6p5tPfhldgoWVJoQ0pgT
iwJ5Fh4BA3yIuEVvjYIpAqHd+qoXC4ArQtzwLtsMf/L9cOlZehXHueB2gpS6wK3qiMxr3SJqLKXO
1LELA73VJEarE4pnzQAJJZDD7QpTaIw40hmg7SeBVkVeU7Poc4R1hspgai1vRPvHWEek6Xt9COOt
yzjynrRqhDfy8BNNiYuLeDv7O3Im1oYqsCxXVWiSTvxdrF6r9Fidd8vpSAuCOfFN9eWcteURl9b2
BrbMnpZOm9Ra050mTq2nLkCY3XzPp9uunn50otpw74FaxA3/+xODRDNEvURgmSngAs3l6V3clnmR
+xGtSHpm5wyNHikwSfcaYQGd9GZxKyVu7tIqNBCLseNCsMMlGYq6g2gr2I5G2H70pEAXkUiu/ned
sV9oxNxKDoRyKe4xhLmtDCn96fxqg7SwPXMGvEqHXXsMP1tzK5YipBJ/tWeNy3wVs7+++JxXOVf1
dokNsj1wprqiAPYh2j5LKnvASWJw2ezSi+MembsPRccAJgTiUXv4ApZPax42oShIJeoPT8ztvCY0
m1TbgI2DqppfJSNsZ/tioDX67ROFCYWPE2M0jLZLpqNPXvsEPr/WPGW/xM1zBU9xNvHIrxZEX2ty
5ESeZO3doi1IZM30/vjn5o5hbKqmwI5vNbdcIXz/RkW83/vXLCG81WEnQaP3zp/aIOibn0Xy+br7
Vum4dxM6y8BfsGQGT1NhWok90I7vENzFOSv2cZAi2g4kPeqkGxGixRGFJ4gTEVARBSUgsto84v8r
q+scEnPy5K/qllDnpImdufJMgtDjVpOaWMWSkFCJIKfSSVGrFBR6YpYMQGZeqwtrV3T4VKEotkE4
Z/h5kBrqKT80iy44C7+oa8SHr5HV0pu/Lc2YjgAD6gdUflu4Z1oVLzyWrP24ztmSgR4JS6tnUn8T
/EIMWQoveX30CGqUMK3iN3AdGLoZZte7lXWTMcV4x2+BjHVtck2MCiG6D0duSFyGSqF5ImLq/QLn
OWXfbdnPZgxGVQXhlDlwBXyM0AclZkYZFCou3t3QUxBKKuTmDHwXYP+Qa25Z7ZOXfna6jMqhUNa+
gCs4863UMBJFNkojnAnLWWYsP4z07BInx3ZarTXl7DzfpnVg1g3WUPapyzGgc3DW0YUlYG60773o
/misWCJixo0QCIOedf+ut7MKUaURaNdg9L2Q39sh5ftHN92MWHXUipu7MZz2vfh4YKbCx3VUc4Sa
Oe0jKeaCi1S75p4bqVAqg0SSEMHy3EfevKUiP532N9/OYA+Z3i7F3QywVKSIFjhxq8NT/UOAfRNT
XeL54UZxo6jsRXXF3wy3JZplYSBrDuNY1XvXX4sRG3p3T8ZhE/RBitx6C8i12GVG83ob0sdPlSYP
kuTCME7HU+Txj6W20ZP454PukKcQJoiw6Xar0P0oqEY8ifJZwqLJ3xbqJI5p0M7J9CQLXK5OsK9y
ok4kEsyQLdPRaAndtV99NLDqHGXtfYAPOoauzbLCd+VyFsyu10VRazzn/wqSBkAg8CREKOPQFd3o
U1eLrliUXHPHXzqzEHLzUcR+cow+0S2xwl4i9zItd4C7Hl9d1LMKKQwdFhlIp0a1SyCK1f7/70uE
6gaILT99aXSJPhibFwcBi6YMo3EUeroPVEDy4QRr/2OKoidWesrReTM78Aa+ZZCDYLu8LGzbYG/C
utNGmu3bTdUPaPPj6ujCFm/GKjKx/0AZQp4tJqAmEyXP+B0o1bVIpI4aD8YsKJ+USheQHfUjWVAw
MXVmmjXqAwlm/KN6QDcoEO1WXMtnChQMGRGFtGyptnbDT+GXluBeBj7D8cQ3F2LVP0+kenokQVq6
wlBoGQa5qE7BMtDOxA+TeGdAd27umdA1P3o3by61HfdlHxBKRCUjM6ysYRAC5cWj3TnD1X158ttb
YAs588JBhRTYaUcNngbKuL1n/LYCAyZ7AK2h3TDR544gikStPp845T661SbEekpbKfUSfGW68tpW
gQ50M1LJmWf9IJ5e1EeNwsHnspWbh+lgfLv0Y11bmviFb7UYu5s4eOkYjMI6y3+vsULMYSCsek/o
dQNYZ/EPMY8TRUdecKeB6Ho4Rv2vCJPI4+ntyk+6Gokd79Tn0sqRoAd4DOv/v+zz/KH+5EGAjMTZ
cn44wXhXo8YnBzRDXzhkFF8QdQkcnEWxlSdE1vmfYQL0tjN8j9n6UQe2dFUZ1ENS9k6ETIUZprea
e3fuc7O+S2vdkPG+EdlwptDI5hfLHhHM87VrITVfm4iLgUMlMMykUkuMal9vLtMJhPJKFPfT9oWX
ypn5hTxjYk323J37hR0SNSc2ThbvDPmPjiKnIS+XW/ByAtHZF+TjNK4onDwi2US+5AGvgxfK6QGb
olYH2tKy/MWdcSt2qvjTYOXm2OOkR7zHcF0gareC9y3pSW6SBuGRVcQA1ywm2ch+/db6VrHbSFp+
RT1QQFeshAwPWAoEkwdcM32Mouev9MyFcaowPLymHrzudbDq4wfssq89dJkWlNIPjct0YDChSYiS
d1Orowgybk6n1EkCJ4AMZ58om/Yp1FAdq6jlxcd0oWc6p+eDlaWL+ujz/Aht8p6b59fl+/RPAtZn
P7C0VTlEnaXwiYeZ41YxtcHJDKghgEdWM+kfKlKJ3wWjU92Gv6U1ERpezzcikg3jqDnc5Rvd75In
AY2IFv6thkbi2ls/dAyOyLf6zUjsFuYHKSXioP1Q21sBuoKTzv8bPXGnuSPkGpp4RtKAc8Y6irBv
DR+KdFxTKlzPq0HhZrhChIgr/KvtqqvGyk3IKsxiztAtd1Zy9eXaG76k0Z5am4CDuActivjEPkK5
J6rw7sv86ZH9K5LLQh4xrIOM8oT+wKGGbLMpdoLDOUwbFw0NLTlu06WcnaLGZdBOjPTDRBi5Vxk0
RpN1PQa4EOb30d0gUSR8MUQMQrTjeUKi1+/aVlQ9pxTjXivaDhU5KpSQaYvG+biZc00ZQVcsdVyg
BIL2ayajEZuXHE4t1MRxbXKrS3wWLNzl1Ma7kXlTyPHQ1axrAbzuuQwg1ezpa21iOb2h88pENF4L
l80W6ALNKZT+/gmxPs46RX8N5f4eZ6uUuymRoq3hlwm/b3cbiXJ/Ujk9MZKE1sEZOgzNzfRrgq3E
/r4yDm4HqwJ6SNzX0tg+JK/06gyvarDLYQinKLnhvOxCEh/LjPVyQ+Zmve5mJhiWTqGxWdBJ2hLk
n6O9y4k0xGScqSlBSMBhPmF+8bVKetfFqwSS1nBplIEf4mAQsFkng6YHfSNLOk30KkcHzku3AN3/
kvMnY5GXjBcwbhldK7IWFzjbjcOFOo5SlF9bIh2ZHLfQ3vsypRZgaNn7JscbLr2byKtO+9IhTMQr
EcIb2WtftX6MaCFIbI4n0PWbyyg6YuNVBeQVGHuSM9DiUZyvbbjV5KLgm3rJrSrC14/seXJwEOnp
2BEhNx8KsZyMeXRswzgfkR5+7t4Yd1jJPojIhZjLH4I+nhoB3sHQJHlxCLMuvKDoOK10W7LC/hBe
wvI1gKkyHmT/8Ro9GV+3piTDzirppr24kxRAOe3yKt7A1h67ogAa7iQfdV3DzRmN3qcK9DkzbqYd
dWyMILs8BH7avMfgrHZLrSG66vWqm/MC3We87L66ZzjC+86NYh+JMY0KCyrO8oRhy1zQsay1+or3
nby2lfMjxkS97t9+awrhg8hdI4mWKpNVyYBD98PzlN00nX6w6KEGvKA3Q0azVp+telqTEHvGIsdp
c2RUP3vJcNnCoecGrNbZsiM5pQEQJxInXr2mwnqmachOIx0GdtMC6j/BbLZbNmDUfRJdxW5YAqz2
ytGRoh1XYQ/m+tqFd0ClLGYqG/EImmhPxmBZN3UMW9vJp76leMpKza3gGxXSQyLtw7iWMYB5WP8V
FihDjIqVr0IFHheITdqZh5lqPDVEiG/niw7RYe/djEoH5e13CDue+KpsEdMzhaaQTQGdl+i4lAPN
U4APbZ67weXgt/xt+nJ1ZMPPYhGSbLDU8VB7piOtj67DiQaiepbmRx+fH/86OSgCT6XQVOXn8gsB
LseHjlQxUHWG6yEC5BSigiawfU4CkXy1nnArCqIHFJoCxXiAU5I0/AwlIeEOHvkdnDvp+iPQz3Ux
oqsKd+FWLseAXqVaWEfBZouZl6kiBGuaTleJ9bKGtlnk0sGhXYQL+h+jgJBWgZqhXNlwFTj/2dVu
tlPXj6vPDz2P9MC4Twwvyk7qvLxJxvmcSgDYG38KPGScjbL2cfinpceTnioKS3R9OXWyL58UQJck
QDMxmlcpAJLkXRgb0og4F2ZHtCH6IBzC3RArLd7hJ8sxrtTZpZJabEXa5FSEMEMyeHe1rGKqQR++
f5XZ9hyIJsiQqkYLSN+wTczDEoKo/weeXwHqFmZpWYb4u/lStZZme8unnZWcnKdfbs8dbTWj2hMk
J/SWVVIO0yCKIWX/lBVATvUDCFvLOcL+BvslVrqdZXTHrQ9IzxKR8Q9RVJkQuTYSz9GrXcs5ai9V
K08Ek43O5mb0rZx4QtpRAd1EHH1vjLtuDRlSuzGvp3S3lof+6lJ+WOqqle9ejwU67C5wipy+bCrI
nfuBkHA8qfECGc/yN8nac0dbeCbl5lFTsnVtXavQtykenc3FWM34e0DO8E5wep7KBZQYFc7XzOf6
rKnSekKXjYFDRmbeYRbywcJbmj6izerNxqn3LRefq3AmUgDaObbsYmrYubd2bzEMdr/uV3Zie6CX
fOSAxHJflQvCeyWZ9DSmezVV/ijoCLZFIqdfhhEF6J1dmWp6plBHGMcINbdU1Z4J1Zq+aoS2tZL+
MxROn/kYoLgAHwdwsWGv7EP+DuXkVQcC1QGMEYXEerMjy5rgifPI4PE9bps1LpcbnpX7Zh4PZLTb
0tmYanWX5IgZ/x+m22ki7D2aSUh3v51sGAjw7g5aGZprLBGT0Cj40QOmkAD29v7ct4ItocCuFzPh
nLZmVZTST1nsxEsFS94lN45Mi5ugZzSETcVx2SwyDyaLLMoLRuB3xH3y9GKK1TbMV4Zccrw29+lw
kqt2YY5ceWncfOwzVvuIdlosDl/w6S/Hg6qavx8sMuHu2ASh1iQNCA/qtwsAve8doyGYjUC0UvLQ
kc20YndhSMHQghHKnMzOn+ZgHdpmEb2ghNCaPxKEppYkIs9CQWMzo+Y7F/n1Zt2whhRG0BFJsVy7
HJiIppPxxDOexuZ50cl+LTXKf35mT2VS5OMszIF6OBuWNbJfvyLyPW3kCp4WFUFAhaN7i87PXuh8
X9e4WYJ0KnhCF06xRNf7uqt08fePRVPwyBH6YuHxxRYajv21VGSQ3vxyLlPuW0AtV2PuPTf/5oBa
YmgP7PVUcAKaRg+WBkaCi8g7lhynEUE0YCDvz7tvWQhQzj9vlbGijHsbwlIoEVtGN6XDUmQYNnNT
34G9+HuVSbKJeDPDda0Fxb4BMPlWg25pVJMxjdIOUs7L+GkEf4h6S3Tq2padxVTSyEDFpUrKyyDi
RNCOBabowBbxrzsSd7DG5P4KAGp1G4z/inFIq8fT8urrNBa3wxfT06GCAiTSXMgn+SfaI3iKglRF
v48Tv2H98GnkFikYXIpnSCdWyAcX6ACz+aSzUK+Nuai1wllfimZnkZTm4Uj/+p7yCr5X6UQzSyXI
auxg7D/KMp1pqS6YGZhoE8s8OKA8QyZ52btOQrmj+SHCmktYEWfJLV3soEBkKUfOi/PGWarUjxu0
HozyVVd1qme2g4NUdKBaV6U8KS2dRCNb4cXAWmZ3DRmTLOVJgbkjcyiGgxomQHK5+nUhPBEG6KUm
p8q77wEITXpIYLohzGg2EMTzkzDY4xcO78m3PZAQtrbI03dXLL2BGbVLKHrzIj3catDJmQn0rBxW
CN3izny4evK4qD521bSVeX1n9h07YRzLR6awBaJQDMyykA3kvlVdd/0NVN4eI65Dp+afyWP2UXYC
h8joB6hFPDVzVjMWMdTmRPsaP6Pfgw7LA8r7/A7Qh7lYo5Op5ugLRt6q58G8/P6ovqD/h+n473Zh
sAFvLZwxFWioqyhKZU5xC2SsRKZ7zeNDhjjmqBBA64gJj4GkwFj8IZbJiSmLb/NOFyrHC+Q82GHQ
fSqvg389WsVu9Qp4+hfLuKo6qDXqsetKX9mFxaDOBap2OOZZSmOnXLTkHtYIs7JM5ER2u88cQDWX
M5NQN1TwfAU/ZbfP3rI0S0iIBsv8B0+djiSj7hsj+iJ8P8xHOKAup+PvPV7LXsGHNnvNdy/FKWic
A3Ibb3tCtJXwvExN/xhBZ5UiTTnrKH4Sd2deQPhH2JM5dXDIsq4hn2da3XAwySuCpul0ihZwyMaQ
XNbP7u4LkNfFjn59dECozFDZzRGb4JMFKTb3pvS5+9vBrzWfhHX7nM/14MXr32LBeIFge6wv5br/
G/Onw7EQl5LeW+BQGbPnUOx6donyBwyeIel+livtCbhEdbgXTzolqgJE4Rksxb4aadSNTHUnwI9K
fOLi1s0b2XTsy/aOav4uRntQcxOsLwuDv/aOkCzntUa26bVsNzo8bT0pT83IW5nEGP9ziZ2u7R1x
CHIIfz8lf8ONWux0f1n8xOuNl63fCCj+WiG6hQd/ogFtLaUiczJ27DD+OVf64BtE0RrPvatx/n1Q
/KlQxb7NngfVeZyqZ3532v2WDowpWQAaGzZXXBsItrc/Hv0dycLygBNV/CMaKtXSLr3EUQl7PKjF
P0vxQM7GywaWlcALzp6dMxxZV9u/TfsESjXc+eGbeTuy3P3LeCIPRw9m5aFMwy3CYO6T+NtC8dpI
nqZtDD5iN5kkQOz3y7ne9RyOoM3Cv5nxOXXvtvLpDcjSnOWd2NPWeMRhGEnJaU2JhpzUTLwgu9B2
f9zKgIsPbvfwELIYuVWoUB4zDY9IvhXVe+XeRbJSueJ5glO7dvCQYwkg32iWRrut0/wLicmAtsv7
v3b6lMoDpFGhJmyNc6rodED/g3qZ/JS19Kj6oFtV6RWMTV8AUs/UbJFtyeuL76S2b5xahGu03mXV
nvInYidFWkBahHPig8fkFMmoS8266GJYGzvRUeTFZ6f1KlAPxjACxrZJHe2+SYuG5R7Dl3JlQy5v
vUFKrLsArksYhjI1u47195UuSvvMyp82dbaewYtnS/tuJ2VeO1D2dnGaDC3i83ln0a5ANv863Pu5
DW7QNCm52ScE+NfGLFZ0rPbX0TTGxjd4lexz6bohcaSHAGx0iNDc3LrrQMd5rz4PF/8pI5O8KkvN
xj1T6IeOHQSzrFNZWstKL/5qPPqC5vfqcnjK0MDdtm/bMyB6aQr3wqAA721UKeyXLGktO/fOrzks
ptm9+vlcJrm/nbCic7ss1etrguY5BqXb8dM5bMiK07fbKIeeLlzN7T+0NzejoeBmqr37TLvjzcQn
8yZotMgb0Huf44+Y3rXbs0OsrzlK8rFvC7uoaQdd7jhi1001wOEsnzNAvuiTe3bmqHGc92ZXinpm
8h5fMk1n+KBlz0CPz33uTWXlniqERXaD+3jcaCkXqfArS2xWKTtLreok6Wmzs2tlR5mvkr1LZ7UR
rnirK5VXiN46v0ZDModA5RAdPik26DbkCrjasj0ZSgy65V44ZGG7I/pbSpIVH9VesOXoHPAlLBXk
zYbDE1p7kvxhMbYcYq6eu0mFrn9vXt9jNFdNMQxmALZZsxpnGu/fDiBYiJci23IZBnIuM9VVo+zD
OMZ61bsNOC91cHvCoiqngVjcvnMcmkWmMO0pADFOb4ykmFgeLNeZwJaLuqmsGCzOzIl24X7C5uqK
ELvSqFstkvEXvTK+AWwPnmYQmwJAIWkVPWgHiUVJrKLWgGHQEq5OK58rGI0qb+ywmuQ2sXLyw+qj
HNG4+uEjAsZoUZuC8N6IEuCegqBoBWPi1TbJ/eYuf8/Ew+Ldd8VuqCmF6r6yf6A4fcevuns3q2IU
vFCqoTSVDHYkdRZMpRikxC15xTil2krzgtpsThxNp3eWEH4n6zpn30fDsMtn7kuigsRRDESnyz7S
85wjxydrQEh1RXoDR7N4P+mzzBQ1RHmhExrfzSIfmXtUXI2tg9iWS/5YlOAUqQg//xrQRORCBpmH
EwT0nKOUb61G1kD6jqbKLQsChpEKVI0/tOEkjguZbEqU87HyCG69FYGB/zSrA9c2yv+idRT0FXuE
pc+RNoUymLL4TDV7qLhi+jrtgE/WCPBhcQx4h8+D1ODD5oGOhpky5eE/IXUBiz96v5pahfQtaFvC
KyiHqpLwNHh83p2DtQunc/aen79vDd86dve898gfX73X7NpoJbwsLNViZy3y7y6Sm3ONj4QllPgn
TfPIrB/wqWr0qMXflrsNZDF0N5IQyu3OAwwWIpByh0T8LmE6fvhLavjsj5ezvpcpzvw8CCdOc+vX
mSjSy13tiKEKe2yV6YknFQ32FxbYw6gIc5groXY+Vx0GFNdEcoBKC8ThTJXnIdHIxJftGasagRPZ
U5Bupnk8zNMzoV+Iv0LCvJXL6bRIf752Ck6T/H3MC0AQGAgEU19RDc0ltUQ6KPli4gArg46A2kVi
huLt9b6obeNXyESVROW481G52/UGbAsvgtU5wRnPZqUNMY/Q9rYg4QYysv+1N3JMRHVIFf5advpo
6JTV3NXQoRz7Fh7GKKAFkTJKKMfq2mrT7lcMuPR8gPZl6iTyJpYTMryVygxDyig8lHGlOILUtXXP
nwWODLai8WuC1VWUcboXfQ8KTRAAHQwbLRwr4xWPRzBbwfJMuR9REpjI2vZ2kvHhwzX3maBItj/6
JLr24kgDkGrJYUZVUMUctvaWd99HRAi69IZD0kHOa439rhwAmW6yk58hgpWUbblTvsNH9l/EF/7W
acp9shUXo50LCNR6DkXXrGpLrNB+ckwA9tRqEraPDdFXILJYGRODvFWgKgVDLYXZDgwwyAw3S3xB
EBL9Er0CV6aXxU915s5uRRZF2zOnFk+ElEM/epRtcUJvkEZtu0KaD3l+9jfv3CrX3BEasa0/M/kj
B0lkSHFu2azj4agUcuf2BGV2mT8a6gvBeEt3PM9pdKYCAxgN0RJggPPIuWmlqPqMddN3JrmYgacA
4WHzDrEle+LfP9drjmsDxlcPgeSi5DGUp6+A2j/F6Yw/JDooUvMH71epWMnfFIQSQq2gpr6uOC2C
dReizydjqE4Yuv9U/jKY9nkA4lYR46Hli0xMV8KJk6KYbogEVc4kyR0oOCkm05BRcvEDBt8zqnBQ
LD0jusvC0TdZWz0nBDBXLxcZITLE0qoxb2KVAQQygME4uqE/ggg38LAhtnjuMOBwgDbzc9JW1Os0
aiq/ncBujtznLT2vPahuqZ5iBjWXoCelXKgIM5cZFVG0T6/5fs0eL1WeiLMfQD0jXzHbdFmVw1w7
t1iMWI1sWM8bP2xFvo6ht8tWFGW0Wc+4ZSqpZx6oTEM+H8hPaTT9YzDHg1zPdOnBDu9QzKZDaHCz
udAhM391rwqriG1j0D+Hy5ACzgLfk8Y1VNuuve9Ank0THwV32vMTxSVijKH3E/DkAYaodvvOCXAs
H227LdtRR2B5ZElX8PvjkXRaFxk0sbyNktv2Q2lz7ji7VOT2dUqsoULw6IN92rUsmUOYMEmBvufE
PZT850nAV10ZVXFrGdfkARPqEfDEQg5QYZEQsrl0H0uye4Jemd6GZQ4rkVY+Xjk4gZn0p0rNFb1c
l0ZkY6th2UwMGmu2h++rt0XD8mBHExJKeaQTeEOXpni/Yg14lvSxngFz2lF9g9QGgy7/WxuKE6vJ
5+8GBASWESKyYFScpoflLLn0OkpaR98OvNnExcweOxC9RoUa0wykUdMucTGB9YVKdEWCF1W2aUGG
u4taPKRYVl2VGPDrtZipndjeM3Cdwm35Qn9vf46zw+pjuGlDHsTTq+U6ITFGD1Ef70VB/ttqmndy
xH7pDI4XmwGQRsqF1c3J7c75GAZxBE+l7RetqgrUhnb4/atJ0flPhYFlDre7WXhQ4JUFNyuyOc7k
GDH8iLZADhRZCC5eyGr+EQWdbN/by2OYN7BvrnsquUYZVs0JFMNKcjUlSKgRb96nphT/VWwtqams
SSug6ncFMZNHlKewu/q1PyJHjepla1+bua6Yg947XE2tG64jQ4s7NPa66TkaaQ045tWJQCO7LBAj
lussIIP/ogF21Dpq8SOayoT8QAjZkirnAENhzZAfHMZaQmCSvCQ/5OeCsVYu+5nnSr134bf51qJC
b2Efrdv8ldmxzzC22/UJJfPieN0UKrtsn9CB6gtEoqq/5AUce6Xm5+rI/rwrlEONOx0ohbPRZgTT
l4s/88i5WAxprYrfyg1INho7zYKnyKkv2CMzoTFDZr/sU4/XaWxcePFyT0DRVq/GGk8YqDYlEcsn
jxU0NSWSTqk4KQPfLgd43zhLSlWz8T/Khne6DRQWkg28xFe8Pnuo4LYbfakueph+YNqiTy88kdEP
9RzCm7hVifmKCCKoB/PRAj3ODNObKj2lAjujM0RC0hqyrUGag4+StkC6jHelpGRJ0kqZNXeTeGo0
qyViMmrJLDOdV8FWPnPojdUfnY03JzDGwsTBIzBT40HqNa3IJgZ29C1/Gidh8/R3OAFIPDoqEYo1
Y4k+zlO//z6Sjer9HfOck1RKXfMLdxJLPPtdvM6BF9azcuPKrYL3ERxCtwRDS4RLeL+DfGFT0gg6
FTfi3uS+jsUlapx2G1liOkEs/Zo1ArDNw8RrGfouupVYe8KvpuEIji8fQVGcyvw+Qy+ohoi+P4ji
nxA/2YxGwDZPxwKi64QbiXX8sKlYy4/38g9E2aTl5bNqULhf6/eJhWtQxa17Fs6MnIWS90dA0zHG
VMvSbE/532b3VKeRAxXANynrZNAZObLGiwlzGPuhqZaBefkwk+A4D41pG9trTs/3t1jqcP0Bma3l
Z9sa42S/KKW1nzhw3Wu4VniiUCULZWbjl0JaZPxPZ+IZ/t1Xz4ZBrGi1Ttthl1spaFKw+lWWZqoH
zTtCm0QU0hv5GJ8YslvdzkDPqnLyLPyspbyooijK46V3Qp4FZKgSL38Zxmmlagpnsx50kwV/U89e
pDOrBSSovpoe1YEMLmoIcDTaBU9E6C3xKOZASlcS8XO7D5TNcmgAJABOxKjzmBq6Pdsz+0VP56W7
hlrtDWNpmubjzW5wE/hg4EFC7XZESue+shghNHBjo33YbD1MEcNyu42EtQrEc/7KZ0/z9Dfqou3D
iwwPHk9Zx/wigOmbJ8F2mw0nlg1VkvDXLTQUq2pnYGSm7gHSDcvt90QX/DDhoAKMxvHMTy5YsIuN
y3jSJVagIRy5u7dw6KAQjty1RW4nAxts8CwrwNVrt4sEVCmX1OLp8T/IYDw0s4USrCvr+2HoW+go
yvEqd+/IAXLWMk+LLbOLv40kxVKzLbHDt98xx7Le5IZuDn6B5f2Ohc/efT/IltEQmGYye3evUzqX
Gmi7JRyG6a9NYvq/e6AdJ+Erfm3cEsfL/lxYH4BQUOUEr+S22XCAKhGnVgNUsixIZ/FN0Tu0poOP
45Kbgf7Okcg7MHSaErCV6XppE6ODOBmzDb5ubmUJ7mvci+2+T/OqXDimLj5qhVCSu6CavkXdb1XC
eqNqYOMmhErBSIGSmEis/aOonX8/Mz8H3Mdg3cNpdT6eKA93jblDg/9JGEFz3Tdpg7ZVdVLIUpwp
3YxfNkA1snCQ4AYIBOeoR6UiFcjSqNzz6OQ9Ec7Q06ZJ+Il94hQDYkeY/8wKJu37K1OG96f/+4WB
nyHNTQbp/2psabzxnGeMdqPjUSGtj74n7erZOZhsFoXIKSJSpjuvXMJdeFb8Ve9ACrKlXbqCWIA6
i8Itq2x9HcSeU7qrDzUOSqt74mddq9veMT7jxUMJhj/tXghu852zdZblWBjSa2YKn0DnTVy4YOH8
KyzWVqInCnhGTSwzICEwwKyCu8FePhsUdQwrDpoBYC5BDzOrz0I+B67myFPCa53ueZC804iNQ3zW
hkw/DYDU9xGq262Ak5Zj8eqGueFMSLSdOK7oXu9nNmEQISUtp35qhFbFSddiYvtYdGxJz5EUjne/
0Vj4Xx/4weFjbpHxm7MELXtttml0ind9rK5tDTjVBO6NdX/NARUs8Yjqk2+gs6LGafKyGNmAqvom
IPgJnauvkMQDRQ1xT5ntu61vatIKX62fyDsi8BIbszXHZtqJkVq7bETSNLT0uH20ZYVR40643tl5
9jW4e4okKmwburA0pmDNyARJVIGxWLY8r26CUjtK30W5f23/f9TdJgcKUgp/naisvSBbjpLJSbXP
t0mEonbj8N1QI7HwVrSKSnQljoaIiEb5V08khaCCOOXonqyvVrJt1cUXbAAAh/42twDKBFQswej8
wAL6zvQwAeQJfN1ScToDYeX7QwIXTm6ZbnMLbRrKZhqYl21Ag23gt3/3OPtldS4sB9Y18azd3eyV
K4byOf/MEJshvOZVe0VxNlsSglKpduRn+g+1ILgVHrwRIN9Jv7vSQV07wNjhOru4q8CkmqnyE9QJ
fogSyxmMup7JoD+sjCke/nFfkFK61IkzRbBiueC2sRIXNqGup75WAzUoT54fg/iMrwc/tcFI96N5
YV338jUmoF3LwkpCRRTT7aOFVSB2lv5S5bWHnvyEya4QrAI5w+ve0lTgilgoTtdcH0D0ytalGa00
t1PrTi80Z2sNyy0JSL6P1SPplz7c3kzSsCIV6qwV6PkFoJoCkJ4zM2lfxrQpVRL2zfEaWjsaBMZ6
2CJas8+dYtTeAKqBr4l/nPkd95S/yBUp5FiMa2MjRqE+/4Hr3Lupmu8fuAmJatrEcZNfLnQlgiZO
1AQvi7MuYxIYMFDMWjZ7A/EMN8XZy4CUqbopCCq7DozNzvxBDQJ8juAJNFo5laiD5OWtpo7ox1If
jCgODtoIdeP3XPpKpM4NtpnvWTdhY0hrS1V2EtM2PUkh0Y9cfoOVdkqRzUJKGcnzGrctCY7Bpc+4
4MKcpDc0S0KuIKSNP1zG3pt9I5hvTzHDN0sM+bJK9l9Xt87drnHR3mpgA0ugzk4mGfYEoqcmyBii
Bb79bQFN7Y6Li80VnIXXJ3ZKF13vEknH8TIW/FGN4Lwcl3A4qZKTsKP6izURgSMVdUQLfsCxxuCU
i5870d4wXClx51rf8YPlivrIvn9LrjdEQmUYO74ZGuQz4trYvFI164WOoDnnExihKaIbiHbDZ7bN
Lf7sZb51T3X5l8revrGVWoWpR2i+6OEm/Kx8rE9PJ67u0WoAXPEbHzksU5vvKNDlIZ1kfcZx8ylW
Ws6dz6jTB+g6PbBvpn/g60NdaRzpOZH3cuhvgE8iBI9mHuruBGFWIGpaq8aUudisC6HKqH8nv9EK
JXbL2hCUFMj4ZIsC2JimINmg3borXlxFH+1ra06RbhMA1ZlT1D2mi/HS6gXum+OmroyY64rkIaFb
rhtLDcfv8DIpzQ1zKWJE4n5apkqLLkOyHtnf8b7YXWfBO+dWcp+ftkvKzP1P4BoC6fpt+D93fesC
dBgsfPMamxCLTmjyJUF6B79S9lgj+YTP1lZb5xN90wR+Fx/st9iocFrrvgl/AfAShmhYo/qrmnsH
HeVIwZuBxyQP1k8AVKVML06Ct6JkFx5uliCECrAxjqed8XQIhWSzYuoQHtkEEItwgczDKG+b7WoS
JwyPnCNni7X0yvQMlcMeyt/gkYLyHy+WDFulurZL33FW0OX20bOAHVdqXThZTJsGj2+h8LynONOB
svxNYXfszahrDAEYRZXiWoFVF6BOeYoyvp3NrhW2HNYsIGHdGA10m59FDKRkeoGigu/aBIijsXdI
XQGT1Bb0O3jtOBz62bJWqbd+qdLhDcO+hF2Nsuto8mAgOhqJaCWHpRqavizu2MNB2eyxmpLzUC+i
1+DEOJ7jXQhhCX2aR/uARDM1tfgH1k304eRBXBR6n1WbFAOBfiqmDMKygKDGc9xg80FBTuOc2PPo
kdQwVVzzbpsKKAkQjacYB86djHvrATtE0m4f3xmCXW1yCi+10Aw8EUv5DXWIt3K6rMSTz2JKSRYX
Fkvgy39t7ZK2oGB61zrl4gzj5SHfP6CKVw0Q3JpJFXy83rDbNxdhawZwlIKjaNTijox/ze4wO99A
zu9b+VR0xloqW52FxZrwBW6lk21ysl22mq2kLz7Cnafk0zNCtcgb8T6eoReAt762XjNXx1i1jM8i
NkQST50N1u6AN7rztFsXclcdSkmrOCtG2PpZv9PN2FAEO4z9RJ+AizWG0hge2dlXz+pVkpsTKN5s
FKQB61WMr+PHglG3ofvEH27wtgSReP69aUZ6trJ1sSgwUmkBYs7CudCsfAl+ctMCTHy/FnL74njq
13wB4NNVkKpK00O8JDud46RKlBdH575i6Wf+Z7pv8vN1f1G2M/kJdCqlVimPOsEYC5PMU68xsoju
jUDamzV31ig/dHh7trAkHo7jM5JI77jG+hSEeaqQnvYV5NyuOy2xZ5oNeDT1ZXiXZ3VT+OfZwNsN
ye+2V6J+zjFJUzrty1X44jQwKWgYDuPqGoIOavnTkEOfb+E0udl53h2W2AM9TBhlPFd32WO7f7mi
fROorab448zqa7k4/YariwkWwq1BJX/WevLFm9Wmrn5zhY6cS5Y0zYb9vf3W+VMYyKkwxplFAemr
Qtl/DwRuFZ6n/AmvkPBqO6jO6ylFgpzdYT59JClBJeW/Wyq0ZSy1gxDzfgkmwZWbTDHYpfRDwWJ3
DQWHvM8tuPUgHaC43TUWHUloIoaSfgdUG47y35cdY1wbwKDqXylZncaEG5+pAZPyO7mn1uYwwpK6
/VOaIEoSosz5fS/cVaKS3RSM6tsFr7LzdJUkuq8uNFxMqo1PrfkrbDf4mZXBWhTa+CItygWgursJ
mx+UZS5YuTYM2eetpJWtCcUYaOYjv0N7DuerBjUeMleNdS+6AU/b6LFWY5EJL/BrbWHpjhl/FL1J
T4+Qj+nuEOBPd4vmg16a2lFOdxxxq+NKDOHZ91DDEFVrZYxetIFig4bE3V6bb6Te4Skzt9uK8luJ
/qKSG0I8gmFsnESQQYUA3FfWl/p7YsyPRbTZxDPwMI5A9+b744Kc9+urKkx76nuv4eXJ5kYke7s2
U7f8Dp/uttoUUJ+Ah7c1rhjhI8McPwc84XEDYHQALDEzhLU/QLaX5K/JSPZnrCTE4zmisOl/KOex
XIqE1gVOQaK/lThiuN7wmPWz5BQsv05M2Kj7pdINzC+qfd3PSyIbgqgh2ubA5YftvGacMSSiGqmz
Udxs/i+nBtFj/pmkrf1vfAeV4yaVAbfMMttWzgXVPGLNyD9IIDt4POHBTFjRwIHRA2ILvKVTDnp8
YIK2k1TTvMPfC2UVIg+j1C3o9MDPy4h8LtrTnwS786QjfOYec/Eoa8bokGxZFllW4EirardQTqYS
WIS0BNLXqcK/9DWRuGoKlUoOX8eHB2QfEmtD2laN/KRzj8v987AeCjujYJt+3jVThqEE1Y7MPyDF
/FZQYQiUPp0X/U1MeJ3GSekBIUT2Enp/SfOIRb3eQvYbbLy3eWTNgpGWfSswxOZ8LF5SuPeTXZDq
PRIBbdZhi5bEBzuVrA59EBBBeQPi6HsA2/SnOUbQHE+s+DYc6qZDXX0gIL797wKWhspWqX5OQLHj
PgdH8J/97/8q6SACCqTuCX+TWaS61V1qGXAIuWQ5jti4pTc9/Ga6gZwTjnN/8O4lfmLecxGipU4k
MuLtAdbLJuNThmqja0ZwYmd3zqBSTHktGGaMRpBCMn6gkXphDtmz5+Z3CzxZfDPeF4KrON9kgiIR
E1X+xL3l4TOpNsKHanBIDuTy1QhvYLJvcvbkAlaHCjQ84vRg0f9pQyXS/lr2DkBfSBOMeAhGL7lw
+Vny3rvRtdbW9NFP6w8yWeRZkFJgEFdFsbAiDp+MozdIeBEmV0NRz/BT8w8051D4WgWejF9n2SZK
cw4G75ifEe8cviKpfZaBB/bWbWIzQIxQAdTE1xRiewI5Mplo4dMTG8ft58J1ZyQkFsWgqhGDZ09S
5lRvMkjW2dMSyqHAo2+scJez3WHn5/AJ3KpuGNMBsNK2SnA3BGldteAKAA2ZWErhe4X45/PPQ+g6
ZeQyDy1UIlabLlB/kwIWH7yrM75qOFraExTx3EJoiATnJjGXb94HfgiS9n9zmYyQZVXO9nOg4y6Y
mdf8/Yt3gYyZhtsjI6RbDYavBoKy58DTU/2cnSA9sRqOYBynJhR/+uyl/cKol/krM/pWrgW1lW6V
tIatXLdQzaOGnlVbSx0HuA7kXKoAG9ib2Mo5L6tr0c3bHyVKPH7pUZRueaEdmwYjSVcWPNt+6k3r
aL1icbOoy8w6num5H85X/3IiJ9osmFlByOq/cJaSK1CQWeVLrF8f9aXBU3GyRsQAYvneotEmIuf+
5D5SDiuqrbv4JibLTeMSx7YqnTOJO8W7K5/4+TcbXlqiih+Wsof7izI74K3ZwSMdMKNBr8bLdNCf
EJJ1TL3KvigxdEGSkQm2Y9UBM2C8vnyjk/bC0VmCSF4eAP2hJuGQ8gLk5VxJ7vRIcDIGUCpwNnLV
p6k/B6BAW+jcc/5ey+mg9ooXXUphvD4ocbpuqCSho63wnypVwQjodEUT+sT9PoADUajqvHQmTfcc
QpGqnoEwo+wNeC2hyutEJUpRrhsgoinLA5fdYdhCgdYITBbxTXiq/OT657MEHUqa+5PHoApLqGLG
UbpivzeKBJzjo20viZQSrnV7y5mKvFYhH9YBP+qju0TJeqC6GkXagc6xVSnGZL5pjBe2gjISGK/M
KbcZ0O0tEH2Y5uhX/DvEWJETwwc0aGwfJEMSa+cUdD8zvD8ghRcHRi0Lfwua7DgPJMUD+W3Cb+9O
H3NsQCNtmfdswJq3F39zNbxqIQdMWaCy4pmh4MfvOkFnIXRQneBVM/FkX1fLsVT8E1rKbXfwv5qb
0nPWVKQO3/9AD7LFsbynoE5iT/v5Xmha0mZjaP7x/JkVTqyXJtMA3uO30QE84yPnSqV/J+pBtkJ1
fDfD+mJkMHqoJrCgwCTBh6beJxKU+pkyUZL8qFpkBTt1vYgvpbDsFCJXvZbLy/3Reo49OJwa+IEi
AdlG0GW/d+5ESNed0DzJM3blW56SBwDyuRWTSbqrAoXFjAsFh07K4B7YO6/IIMiFnf8ItvMBR0Ys
CcT3IuaA82kVb6Pm3fjTx6NL6gR9+9EvrGGADDugYRNqp5x2OrxVwGbCpw3ZBx03YcRxQNQyqYbF
HgtLvJ+MiZnCV+hV/4LigG9r7OEcqUTnhY4oFTQ412qz7+Ns/iXvKxZfK8wN/Oo2fdjhNcP7vIWg
Liq/m5u6supPfjqluZerHnroDp0zbM/xuagypPJnCRW6GoKa3ZV3OVSws5GHdcP6vWe2pDU8fmMG
jHpYyS9yc6Q+Y5ficPYwteD9uHexoZlGl+NJKOidOhUW4oFybKkJBXq9qQ520nFHdehDj9pt9qeG
RI+2DynggnyG3CaykK58/poGRunseGl8G9SxeCgl2FZ+N1WZGG3CYCkzF8OK/Cw8VcOTnvXaF7J4
of5DBhqM7DWs+qun60wF0D1OTPpYemQBF21oF0GMYauaIoKm7qjC/e6mdMbySLGdDCChYqNgSeXG
FWgwrfXhDm4yolBoqVh4m+U0NmFD6TKgkEyZ9GIOH8oR2ppetnsUgOQNwkMONvqfiErOT2vihY+/
TvZzJlhEXs2VPP1k25VLJdTTt0E1ITQ4XsBRAQxwODJebHNY90TQ581SbSrrbQe/yJGo8PKHw2bY
m9b/pWln4ge1TfvCUB/gZ51ACIgWclhRft6sUkWK2eA5r0Of27twToa3Bcfao/A6yxGshHSUUFyR
5hm/jT4mQAddypxPIzimKJjXEyMsOoE5Xq/g5Ygik6jCLgQEEwIAva91OqJ3A4EEV5UQuSI+vZPb
qMHnh+7zgaeBgwzdO6zPwREEKi/OTgp0oy8Ty3ZLQ9o2zK7gpsWOwRiHvyMvKLIHkfcjzPXkET63
4iKmS2WL7qrvDQxBjSrEvKzwTILndieZc0ISu+C14fBiCJkNtL7MPQfmx00ceEd0hR8Bc3WTpREW
QsQs7PlFzoeR1H3At0bRbMaSUZctTTm+zvQp4Lsen/q4/7/Fi5x0Vm25d/SgZAI0WaOnJCCkpcDf
Pb8E5edoc34YJzIo8edz1kFagoUboF3OhGkdvB7Q1mkKm6seS5PvUZKVVDEWsYWbZclD749obk9K
OhjR/rzmzGI8fHdwz4hZemaWTdDJqBD6pNZz81REuuLIHguyipaIJtcJsmIeNZswGck7POtbnwHu
SYRB9siEOXnJJejq+M+qCLj5978yCPOqKFZCZWwRI0QLTIf6aEQ7aZR9toVh9eSbc8pavJn81top
vpXRLMme7rrZ2GucoT9jcBFKIR5Fyd2hngYwqZodNDYhJ4aXcvPY4ekEZz32Hl2S9CHVlEfiCBIN
tdbrJYUh+Qx/eDysJLsyvsQN8n1aJ4SHXUXrluOFKiZdFG7Xve46zTkmx2kCSrI8O31OVSQAHaDy
tsVoC0z3kGNOu7H5dmdnLVa82toGHCtCEj7YYinycDMIuMTT36tu7NQsNzTO1N2oUgQz+NDw7oSW
BBooJ9533Y/KBUuwLxnQpouIornFcdNdJEMr8gFyS8dKU3yyWMQC/4qc+a7hAfn96V0f3uvavucb
w7UCi9slnHagg7BgPNYb1XECGwZvUTuL8qourorl97x8qdgYkhqD0SuuMUCQqgNBtpRakXtC74wv
FkZO/c+S4dvNdqgofxjgYGcGXT+OKKguhNSQcI1IBMBIBwMb0eiN5OC25ti8Ea/NvjvBTFUkgcq4
Iav0wje71tqhmzsinTzs5Mnc/934eym7RiMg2TByAMUViWje+NoY0Aj651KG7t4cqo9lBF8Wawfk
dyzUuPvlBsAD/F3y0MMA+Ge/6NmMCaGrW4cGMBQx1YkLNcGZlCW2nPLClZBYt6uZIDJCdB/RFQrm
IgLaWcSMtFoeUAvxDEWU3SE9tNYjztVkdBfp3Fziiktw0Vj7lE7lww9rRvBT+tvSWh9kW3O1LtbI
q50VO93NnQBW/rOEfMbH7m40/zjSDPvmQFQSHuqlPwBGHKZTO5mkzTmT9wgMm4wezg2zN0pnc87K
Ytfkj2F8aD1W94CAeK58koZn/RZO8RoT4nQNCsvBSJ4r5XYPN2GueaF7gnbdhkSaGF5A/IOcRAgo
+JWuiaIYZWOgNQHmjKcb/WGyUslni+P0C38ffO8l9UTjm8RfTC64fMEMISx/JiscYxaekAV/CPGi
GwjRR2i9hJ/AKXY0gsKEBNZzsMLj2z7pbh9dmSMH747ruGifaBRpdaFP5njAv7V2FwiHir2G4IRM
6cLPnub4+RiZltge3TarGrExESbAb3M+/MX0einFxS5OcVP/wMAOX58HTD6Mlg8ITSx8+4eviSvN
jhs2DVjFhnk48O9fbkOvdRHP59i0V8sD+5zHz7rdoKO+qBPe1BxVH+kQcqxOZBgZRMaWGti1/R1V
LlQImZNquC2l9SQfax50SwcbbzKb+4tvE2aTBd2FwxH6zcdF6KsdacAOFOFNFfJRQnOrE5fucFDJ
SmPPVRIYgSkrHOcdTjNUf/qV0iyx7mHXBMLQiO2cWKJa6P4K8iH80wogJQ5TNpodPBcxXYtfcICc
+Qa7sP55zo/WGUJIPGWVyOWFJom2TJRjY5IMTCvSUfgUBrRg0RqFGlsI/ArDaMAC7/2hB7To27MC
XO3HeqIJ99Mylt5MeY5DFCBDcRywvBSNGVF2ntwUCFGpbFaXp9Z4WjAr2Q0YdAeQcc4GdicypjxE
sQ0olRam2c7JPqFCvnOHwXGUSEm/BS2RmW8A3xYxajyodA64ltQqKV6miIKhVvKAo26FJc8x1MGu
7SRNjBakCcHfZv61UssV1A9qI97hxoAvuU+WK1eBrg1xlICKyLrqPOBVtjBuYj0cAhY0UWbN4HHj
4WvMOD6YjnpxRvzooN8Gf9u+hzq3XjrvzFqZqt9n/ZE2WSQoXOCHnKBd6iyka24+Vq7VlfXw9La7
ObW0cyZjAoBthJfWPbjCIAb9jUbFRWOgedJjrOzHHq1HwytkriQra+kPj9k7uWPo79Nyz8n6A/1c
oBqDJnv0xT6ti9c+IqGKpBx2dVFFt+8pLq1fvv5Nw77nor+dG4DLdFSLQJfpWoAlmQJc4qImAGGy
ffROCNsjetoS+Y8+CTTZq/pPN+Y0/6mtHO9+NOrVvNrVuhi9SLsAQq4Xzsw+RkadLYY8RRqbbjX6
qAt9Ju8bysxaLYu6O2kd5PsThlAauAgzTdm0GLWdQxBMlzwXZ6WfXosSJMed6apfesuTDgH0uqbk
1oxE6TaUXNzkNbTl2JaMImwGofC+RWuoH3m3YHzoDw80axW04vLqjT9o0+GqsQK4z0o2OBkB1xkU
XlQdwhpRfGDlqgI2EEO9lBiW5fP692KF5n4zGKGXzGHGmzUxLWyHIM6/RyqWOkYgOg4VBimTgJ7x
rxJXZ4aXewnumGhTPq1Q8qtz5w06D6Bdc2pkHN07+mzXIV34tgj/mmXB2DrrvAcZwfew/4OxcqXt
ZaS/rq64a5ISzmnemd2OxQAyQODT/LF1oHbSR5tobY7V8cRMShITeYD0SgzCAANADF4NhDnSAxsw
xwcISvSYYGttyUJpsfDt5D7clBPaplISMCqKV/Qw/AQBsvYxmNCuTu2LvQjRpgUZYN9vgDeIC3io
42eKhBg7fXb7uyYEnR21ksfJNCt1JqDkoSebGprHdh1uCbwj2UZBM+CQ/zJXPPenkoXK6xE0qHpO
u6f49nui4Wq4VJGno7djy0HAUTy6qvMNuqFp0w9Jd0lbf+ulFG0sKNV2pnXeOPvEY9WAk6yqc9Ni
+/zfbbkIwsNYsktxB+y9dFqwqH8U7Rysz87KJrnPGoCwhHWhENUq2N8LM+F+lvCdR3rqAYo6w+Gv
Hs6Y0BK0SB7xwqzjiSvymu4Qc/XKxZXpswJ/XcTQ5gi2mE/bArTzUbqZ9/ibuSC9KjjEY0QFB4zS
e3jywi+tSD4revkoRnJ4kZBehDD2nxvDSM8jEoACZD2/wEbUbqkSeoPyVZbRjDWhK5I0/TZXJSoi
dRGgGxE5OQb27SijM356vPmJ5bZFJVjXj6DzascFjQOpHBYEjxO6duLZIHdpDUgMOK+Ff9cFacV4
lPGKvrwY1AhVZrEMD8wsqwb2dMwgMmEwCueVM+aKrX2FbcPr2+ZuSXYVW6IOBXVi1BdN2sF6C+JL
pUCUUCeo9EgtgtfYjuNG4ldOweaAC4to/k1UmXpv3LP7qc5CHLHM1k75LjSr/DH/MhQ3MoG4Nip1
gZhLMdXYAFJ+8Y0/qJNlgqsYpYACdfXtsvSganjym4/NubF2lcvcEytLU4aEx2+y5XxdN1yt5Anp
7xvGOKOt5ZilfacaFGNoqjQ4t84e4njQmd1rBokNurWD2I2bkR8JBkjKVntDt6XK4fveZCfCV7n+
NTl0RBsBDILG6fhDogEcP8dYTheFu0Ugi+SwSEXBGaLV5i0S35cOlUPUzyTV2B7cpySwnTIF7ux6
AiI3mi3CITY9PJwWzUAlfNZinVqcvKu1hiDqdThYrq0BgCaRkIqtvqrp17XrHZzR+w6riG5Om2lJ
wURPUlOQvuFTzXWmn4WUe6pukBQ8DtM6ZXhNnT4TqeNnyeXfdnJSzbUns92yWlbk2hq2Qqa2z50S
9sD7/us7dbJjCm2uVKA58y1YjDK92DRObPtSXXhRuS5rp308nD4nVdCSZJXV2wQ7cYzqLFT2s37Y
jT5hqwEmL2IRf42XAXrfSnaG+Ecv+v4nV2Pw19YyavGV8WRYxHN8X3noo/15Jb8Qcam6v0R+YzrC
B24XWIkXJhp8lOZN2r6m1SzhPiu0UCeeRiQpjuUQWTvtjMd6Sf6M2UqZ2z28mry4faQ4UMVIAruY
dUBsj+Gj4iyEDtQAYb1Rvt3U2TOCqZVyVMalcsD4dMELrc4NzNzFWFm4hyMJ6VAakMTWhADMZ3hv
DmLd1WTQCAfvnoTxixKRxZqCbdnzIiSdBONtEOrXVM4lyxCqHtbvZfyoHGBOLwrEkV3aUF1haMEd
4dCNnEPFIqatkLY6R+0AdmXI8qGa4WJ/DIJSecTxE7XKiYecPuDRIy3v1TsiItwfEoD/LjuUWBfu
cT2X4IOyl63Gow7CgTFwSM3JNCp1MdxQokXxgGmj4bgSGkR4owzaLRZ5at3GCCNo2KkEtB0pJMiL
aHwJNqdUVmK1/ZkK2izs2NFiW4PJ5u85MlDrMOjn+1byGeEmN1wZqJiC5h2UF3End7ILlfSDp/pO
T7IF+vIpfxvk9AmB2otoC4x4Vmg5Rhq2boJ/xCY3gvDLO5Qr0wysRE4Gsn8pb4P0zemtLl5PJag8
s18x8Ipfp5XXwq+bGq97iIU42M30h8TAx7RhXsIvHaKVhBlsv+xjcs9O6K+NRSc+4+OUS76cn5SE
p+dh0ubS5ABgkYxljFn8R0fa4ZV/B6luwAYi3yenYR2a6QMBy800fKCdsPHMxmdUYPzQkp9cuBN6
wiDi5wmxZt/HurTZ/2T0H8HeCyHa8XjqM5iY27gYMvL5eLvHpvqBAn5WhauaJ7/gTPYkPrgLsw8b
wGOxYDZVURZI8V6iLH7T9pTP+GWvnRn4IWHh5BFj9slDNHsNKOIu9cniuV4xjF4BKBTaRXfO4p7a
BzizekTOo9+46hkEFHSVkxdMzL+BsD1pAJIeiCySPm6GHBMthRt5nQEx4C8+cXSfuJ5Pwlp+PySj
fkaaM1GloDplStRMC1qe0XMdzg7HYIWeQ9y4rov2q0FUDHG0kkQNXO5LFhIiGerLCEYjEcOFzgsa
sfIT5c/W/fM7F/FJvisOPwNXWis8WRr55SV14otnemr0FbGl3GPm77pXA88RQQivOtFFOH8EA5+z
iiBsEfFugczpESjodhqj9O44un27om76EBaRdTKS2JeqJCJoHSsgPO5TpRSTPJp9Ad6eoWNbuZE1
qFf56n4dLpS1v+MT6ZQJBCob3PvW9vyAwibkkktwNfYFLhGzVIlyv0yqSwyi1Jk84zgoTGr/c0k0
xtgYj1h0Bzv1xmk99zXFVDDLfEFal1YYTe6VGWfPkSQ+f0pT7K3MW17TPfXyeUgvWMo3y5ZFDo02
IMlmgDV/JFV//7RssOXjUR9uI20pCfaHN/8G5XKy1xwXgDC4LOAzam6qrfBGLh4lUVVOG5bLBxuV
mnxbizxppInymRNQ8TwITjnbmAQIx3yDDQB0+7fLk1hTqQBk5A3SgbOQ3C8lKXCJwO9vZ7HBUzMA
7l+jquU76SpIRQ33cLvCAOGt7PdWTnxq+z57KHYSqLrOw9K7GVmiHfMNUuQbUklKSKY6GRGIAAzr
ztL4p9ok+zvHgD7umy/bgwUHaOQ56igGPmr1nv/vTF8gQ2BqqYfyCPKaTZbDBIXPHeSrgopGWBk6
rxO3/iMhHfi5oa8EcCAN0+pCk4hJi/kT3Aj3VQpezU29Msgs5pIP4tieGi5i5nGiAzQWHHajqP3j
F0E/CI6XXfTMa/2mYAc6PZryMEHMxmpicxNdTpxNmnvB9l0bTV61T3rFlC1r+vQsMNFMf2xbpUQv
w6VYJZCrFkmZESf1jZyst/SHrTd34FrbNeqkD6Un1wJ4aptSuJwlQoa49JVktzAaQiTq0ucm9tXL
I8fNNtj+YwQu6O3fqXKLEJqBJY1IxdwvQJ3M2If1JSSQLtZxWisgHQfoMnj5zRH+sAdeQ26PX4Ga
/fBHQuh7P7BM9xnfdxGPBnRzSz8j/Ah+YvurniL9CxcyXJKDF+qJswkq+imCWpO7fQ/bVU5S1Umw
+8vuR4+2RA/8R0u1IJKini0VK9sn9KSg+4sQKXN1g7corKfo5+pN9dx+TJ9URSs5YX9tP5vZZZ7g
6TAHG68SAKxnY9jOYjJVd+3oD2vZs0pL2tZ97b4R8b+/K4Czal6WNbLPj2g2T0dpA42QcnDuSNP6
5Pu1XWiKZ7XYrvTvF+ECt90Mwg8B3dxkd2pA1OrkCDvcEZJK/QneRi4VYn0/SbVLz/fE/KGIncVA
EjuysWe46SRU89uL4+v+Hw9LR0Tzck3ThjyEanlp5fcBX4X7n8bTUSBQLvsAugkf5w1qsmipbXs2
Vb9dBHVx8QPEEOTOzLlofZLQ4K8zkNlI6+M02FA7phi1XiMpjGAlQV7Emot8dSEGCQ/svRDYtpEE
ulwYr83aZ+LaYWQObUCCNOw1DJ59BOJiexalzsEWVN8pLkwneRVHAUneXGctjynjNWAgaMYfQ123
xU2nH55bRuhIULu1OrBhvN8uI9SqNwbPsKUPcv3rXxfBlbfGHxsaPm6sCRFTw6xhzF4hKTAXtsQC
HJXTnmQMPYsobiNuaYef8I2AL9PGGPztqoe33Q+XHBJAN4QF/3P0iUVQgMcRSIveDYXY6/Etkuc+
oOlI0K6Q4t8l3SCjHJSKqsxL+neskxmTvbFh6/q9zoyDCc4J7bk7jp1U9QfoGMRlA4fQvqS+ojxP
euJjeRoKfHa7kgpcd178rhFameembsGPuOs69SuXlJ4Dcww7aPo3A46kp0/matUmvzme9keo0FTN
XTotfiy4OAwVExYpWUKd3Wy1I1VCyOgn83uEwusVy3iycCW50/+ChVlqH34RybRKkZL4HdW9akxM
xPx4j1XFJfKZHcvYH0EX/Y4ETzLN6cVjwEES7OP5tR6+SGTEUhXemz2mp2spknS51eIi1USt4gTC
K1NEvhMhn3isRf3RDSAC62mKCRY4WQQykEWwMoQT+5vbvSC36E9LApmKPaYzA89dyuK9AB4OFqsw
w9JGmblCmNnBaAyRLFmntohv8C6Wq4YfkUHh8BroQyV2LKSkKhxvxqsB1UIvC/datR3vAD+gcDkZ
wRm5qVDbdAIfSPIWUO2nMKWUd9TepxlPNprEparaFflNq8z/H9ijDUGGXA4B/MtHJU4aSLmJMXTr
0XIGHwXaW+hvK5nRmpA354lgUbkXl1q4YqLW8VD8Qc4BZwaF4gAWplLIwn2ZV9JlLv+SOpwpsZXE
w1i8nWt7T8vXRTIfZxXWUraTpVDM7LZ+jJm7FzGUhUHss17moSOpjQ1X4x4pye7u/xXRxQ/LW+WU
UkvzPgM2WOU8k+8VsxAKln2jda6n2bN+pPKhB7nMY7ZjLbe7OwC0Qu8swd+zA+kr6kthUJK4xxBF
myPDIMLSCbhdxHro55EMW4tSMyzPQwgeoWTbBAmY/+2rls0TGcczE2hpcfsdRt2sjugPZSn33h5Z
H+ZyDylzxIB6zRqA/DYOb9lBjda8TgGB5izJacO5v9JbbM0I3OW3Rrr2vvWIQb5QF2pnETcgDE61
NOWqJey1yqNdzPkfUIdqZYQkb47s4l0ASf8Yb3la7g4Zvk/Z2DZA+LhPmkshSgfj8UDRgFcTdREN
jSTIEitu3WNTScsz13Zx+ksUQSWEiWcD1oLo8RynTU2sx0EmSwlFUx/LHsGCw4A9sWRnK+KxKyz7
mrD+jmvAssi59IXixKXH3OmDOy2TJHVsRS+9LQyTtUqMDneRhTlvYiEctw9b0XCr2LGh3OztLK4w
0z42ifvGv9EDH1P30KhsUsiTm0K+VIktR7MbcP0NypY/Gl7bNhxoivfGybm8sruJf5JvSOMp1ctm
+AoD11vAjHUTz8KI7Ugn1CQ9iyM7VnI6D7Cd1SDKCmrQtxQ/lICF/LnuL5++EzoH5O6duHF7/cYa
utS9hG8tSpwP+LdebUvP3ELmjYnIba5UMqo0bDCy6/Dvow6z0sGRrayGD1+dF+lEhCeQcnEjIowu
IKbrKcuhxKiW6hHA/XjhmRkOsg/LUtf+9um3k2AziHhTYDaiYkft6YKgS10O2WnWHtRLedRZi8CJ
DnhYWtdqn+t0uJG5BqzeAw1LGATFOJGFKpfaC4VgiZIZuT+fKi67CYv8GincIFlCFEsUiKCRwRuh
lFd19YzGxK8s/PswF82A+47YPmCBZFVe3q+jjWV+NmWhNlRRKhKp35d9TeOS6vDfAffjbNUi12T1
GlsX0sXXzY+HrS26meqoivH/rOC+B9nK/8dVphMTj7wx+gXsIu3LSWvrjrq72+LqiN2o3+7UOLWz
4CDEihCFs8FAJnSc+ldSyufJJELHr5i4EHikzmdzYTgGyrAdXVBdpUsrDbpMwzUCSH8/ewSAF6Wo
Uk7DPLYxeyrFGertg4exgEBD2/jc3n81F5kGz57sWEB50x8q4rvpKDM5GgCLo8FZ6Vkie6SpEalC
eALL/+QF2WRxTmf2Nlryv4CObv/6EbNmDBoDmd46qhk6PfmZALKYO2+ifvTf9bPJ8BBQatGrRKbC
inrUbk+ia/KUwSD29J9B5PJ7y6XniLpBQyPmztVBFHp5DHDKY7A+WG2n98quhsjFrtP3JwBA368n
lI1lRWWr4ocaFYn0zVjjt7v1rOLiLyiYmoslYkVaCe/myw8VyCNnbvnDIlGZcZejKsr1nFRGubJz
uweXdKqH9jW2mq3d2VQx0alaMRkcSDlLGmM9dUsmbx6WyAL3w22rkO2Vt7Hw25rjfULCCDh0R4Td
uVr2uoAorkYBYQBFBXIUysqzkfs6DBsGAnrnQ3DMrqDYxiPrr1daFek0WJXi02rT51+PzJY1Jbdp
WpUnyBILzwRqHPBoGGXSTJPNaNniyEXcapOQcUaI0klGmu3h+QfgVCwQ3hVjqZdyGga+5EowRCqV
kA3ilc2l26vujO0iR2byzsrdTtQ9sdScy4CmAjp92EWp0teXdHdJ0/pliGOliAqUx1u8IvCWZuvE
JhgSqIkwUzjiceERT935ScbwIr5F5Tik9CAGSciSDW4yjjWnkofWb5ux9VCmbRLyCc2PUmyJKUcr
zL5ulJUepzYCnSpvd86HeTExHbASr82E1+2uCINeV/DEXHYkX18tqNAVRICPULUoPAYn1e6A7z7a
41QniC2vf/RTkmpgc6IxszUtPxZ6YJwIWDUzbpOxXEFyKHSn6BF+T/UBB6ImFtQWmWKCtzQDMDUV
EzOxiayPFegm/fcIgbu/j/QOfTh3AJ6JoLIt975EceR7FVd5Xp3JlzojNAir1BOF7WYEF2xwLHo+
gy/roBnsimcCI4Is07Q1bCsa6uHFEKGzekAsORMsaeR3PpZxVMPRxsbfNyDRKdLHvbuWbQyKZAKP
0naUEx3L0qDjLdSqnrG8Oj01uauOpyTEx9MNGVyUU+9HPHwgV38FUCo3IEvlI06bDC5VFG+TuB55
kzZSKZircViw/kORWm3/IAnP1/PFHvUUaTXBUrK6d37dHM8uqcHQmFvQo2qgo5OY9kXIrWj6Phbb
B/wDJxLCWSA1p7VRhgujvhZa6lRz8ek30PV3z1x6XlgMM0FiPoNTvw4SiH4BsJX6Kx3C/Bofvb8v
GSY+xvcQDwujx2Qk/ktAQs0YOh1Mbs3A+BhY6ZQDa4frKQRKutDAdU2QjlBB9yImM+7xcNXrJL63
HFM/sfgoid6V8/B0PM8LWVECTc0nZHsGIgKUjee3jYLlmuLkT1o3GcwzCk6ASDosBJCn0gAryZYB
kRoe5HvXT2pxiAxtDH6sETZh2uAT4Nd579Z/WulLnctZMkzVV45QqcJWPAnTYRY6vLJRGV8yzCAi
CdJ0B99veLLufeYcgT9LP/9h4A2t3foTb3120SAcI9aImBea+hCeLlmjAWZNp2VtQwIqGAxHyBd5
Q71djvPu5IVBE9iVmPGHgGf0un7Kspb8i5orSKphq7ofmHwkDIRjF3GT9GgpO8YZX9Rg8t2Z+CCY
1gx9dv/lhJ639w99/IMIOFi/lap4nMwMX9VF6DInJwmGO+O3WK+dxCiwZ/fJu6xBjPLk0yvf/Opb
xdKC/XjSPOr8tCiPL5ar4U2fssOasUHNdy6GaF4Q4gGuJo2XlKyyrr4dbR8xonBr++cziNbadraI
zgsgLsigNT68Xj9jr7Rj+GATy7wGw88lt/+DzhKTsJHZS8D0Rvkd+6iAuPoXMQW+RcBn873lZqsR
kIMydp2mBjXBqsMxAGn73T8kC5eWJS9A1Hmfbz0a8+Zh8I+XpeE0VN9ZfeKRBMYbrd1je4VA+mbL
ASvampR9+PcjKcb5KVM+DYZ+Dp24mZuLFRU1HQ5cAP/CoRbquxkS9JonV5fbiWo3H5r7dfc89g3l
eltgQmWdeTYEchjgZz58IZHZMFEovgxtPYNVLK9ecjmgzoPrM2Ki+cFLcWycNPRF0FdVcpnX7P8o
eMcUlxqzDw/lmBThcy+FIRMK3OQkV5i920HNGOEMCO8siC3wGLPd8pKL8WTDi1ldGE3SkLyU9in0
ZGEBP3UPdYDTwLarw0vTJnbjjopGbaX45F8OGby3SM6/8ZHNmUoPxvxPEq2K/eWPOK3nnmrtV0zX
rUt0+UTIGG9eEvTDMpv4ma29SZHDE0e/cd8hnP2dc9ThDszoEHM980FBA5Pu660771gndgg3oxOG
lZruMY5sIGCup3NjDezoXE1ALIe2swgrUnDLftXv3ekRjC1bZYFkOy4jbb4/ZVDfzDHeD0j76CRD
hd3g+/kp+yTbJh14dGIM+sgxQJgNKBVXYf5Knitg6wJ+BLiUN4IBEvCDbHXnFRXxHjhbJYeDzWK+
8hL1pFluo1ilGUkGovnleSnhzPEXu3X1yfFwlV5hnWgzsm9J1SL5tUs0oJAkh5kVITGK4icJszLb
tcOoMRpMYnfxiwWuDipbM8TjQkUMIfzDB+HBVXDxnOOcsCJrZbASKYVV8cydr/MsJpS0ghYR69/r
isU0r5bZhGFHcLiqOfODUkNTxUP56s1QBSMDsQS2ql80B/B3+yBJC7/gMGAdPmVWVVJVU1csXBSd
foCwj6Kh7XNGMmF0ZB2Mo6K4/xicJYkchhv6ylnevcXuqIN37rrzye49Y+PArU3Jwlonz6JnqIz2
JP8mN+BQI2cWNOj/46NJYMSCyeGquybpksBtGdb0iugH11OeP3vs0wKiY7V2o2OeErPg6eQdN4on
3BYUN6avpnBvOZ63S67Kx4PyxKzsF1ew2ytIepgC92VdkNGBprKr1U9beIXTEVaEJ7Nxf+WJlx3l
kgF0d1iLxIXpmxcmvUfgQWsHfbzlWnoGCyj1aTi4GTP6oj+X97hV0+7FuY5uQo75urcTr68Xs4mN
2cZd3ILkBQ2RM0srvDFq6n1gUNfW8tFojjrl6aLQjqh4PZ2OWZxEeWK5lA/HodX/uAon9CHqQiqb
NOXAn0fOY1iPgsC4D0YZSe/pFkdCk7+Q1uRmovKiqGZOwLjy6mQq2pZJI0OPItgSJBVDpJxxbZU+
TCija2lGboj7bm3GRXjED43TeqycIVD3orD+Ov8QKfPOsceApkl5r8eYC2i+b06AnpxreHxve3/w
Plwgi2IHo6jYGb9sLs87lR1JLUhyhnvUda0jSjQZMvJhhw8qWXhW2/KHQQgw7fWTo7YvIoJlknOs
KDZozICoseu+pdH5nfeCdIk24SJELwfue+zR5tJNapfvBwAysoi+omcJeL2xzg9K+9J/ZcdteP5g
XlnpyqJ0uIkri22mFXgTU6gyhMJFe1f7CaVJbbMVCZ6XtBUouDLbCLJCbLuwXCAkB/xYWLAJ98/W
4pyKJzsz+h8mknk0TW+k9IvrOcUZTOmFplGFJUNkUrhjlBkcqiFzo8xsSQyAzlQm2QlSqBB0iiwq
DwXHEH2U3QAr9T3UxXnZiKTLNCjWZMMo/IxKdEM0skWc3TLIeKULBd6u5DwumOWhQhdWOYqX+0Fr
944UsfJvWC+kYs3UDLk6++oAvgLl362AgT+jKPgTm4lfAXtmDFKQsFkakowebvo0GMxE3HKnmUfp
5Aq2T/5cDkG6DA9dmSmbHEt4JWNzXVbeFewfWBlt1pG4rOGerYYsuh/4+UWs7mUHFcOQlskMoMPV
zeqgxPfeCgMFBKdNUUpe9KLBoloGZA+VehBk3J7wtLszuYjj8K8eFUAuLhCQbj+qn51ES0cfrfcQ
CVpaE8xBPyXzJDy/qVrP3gLQYY4sJwvDy2a/DUURF3h7YKRVyOwuqyVqfuD0QSZwlo7nyET9M7PB
pQIlJXk6MXrc3bCS3RpEgkYEXPC5HgMWFjI0F/7s++dciZioD+WQmqUTRhUdHkS8p5HbRydDyK31
c5egnvmWWpKSpS3GmHYXUdoy3IMOvkmOPAWLtZpAKLgU/0rBzlKDJVLio+VJzNUNUq8GgWK+8jPu
131s+Bck34UG42S6EmI4eNtY9vJQydTb6f7sWMpD23gFQQZKxgvH6/I4pLjMWiqukJNs5SZ9lSvl
yDnhS0iM7Xa0mr+Yjt0Ydzl/lYKKEXI9JxjS1UBY0KqdbVe0xqNw1IdCHb1RH2BN6mBB0N1EBkJ7
8tf7eEj5kE7ZgNaRAmcPLIRvZEXlZGyl+OzT04vmyvzTGijWBYD8FZLONGrhp6OBRm5vp0H4/3/s
DW+9U9r8pPKyuRu10hfD386OpdegUVadljpVvghGET2kjDkN+mesdIqiqk+5z7Dsd4pBlevtxkxI
0vr6aiXNzddiMn6fUh7O0l8JCREEW2USpFQjT8jM6Ds68xtbzCi24VxNlCfJkG0KmNy9M4GXLN4t
YD4rbJBtmDiLuB1VweKmq2ACGma02O+SBBjAY4RwLsS4NRHdswJ87N+IPn49Vucxi5cOp6U9wL0H
S13SgBFCKnOl509+tu3zgXtxD6spbvIh3FNUucZ9rcsqSzb7vszk4NYkJG5CyE+0mSsY+Sn0PVVM
RUhdHJ4ve9zJdv0METMVjohsyyUTbxTVmtNBpg4LwZ0rAqE4ptdQcDVqHSV4RAhAJJ85Qx4woxg+
b/Td+p9TTyUN36Q1j1DGmP+h6t6VOT7ZgD8nct88LaRJjeVeb5dZgdhjQwtIQsWd/y3O4e8eEJQa
M+loaPNrNLw1W+oQtv507gcgMYigIIfx8kvMPn1LCASTzoNoJlZCaz1d/dafrLJJ8e84l4KsSf9C
xlOsKcZbJ8msjxfRtnlOAdvO34KKw6rfar+jK5kTvB0Bl902VT10xmWt7AkQj3w8+NNIOxImy9nY
1RJOP9aVN96mUwn6LdNj7zNNnTW7KUHfXRJ47e+9xsW4a6u+/0vvKcA6h2ZyhWZIYs7AscxPnzQ5
XpQZzo9CgHJdXNYmAfX3iyaOuiV+uZFix4pBT766g7/brCT4oNWn9Y8nhDw/3vU+6TdNlvZWuoQb
pVJdi17vNSASOkXHQhgwEw3MGg7a9POW+/GGIKNs8ImZe+y3Fd4KBLX19fHcRNaLdzoUAhclNX14
OLfbRfaGosxrO5YgMJKM0UYaF0XFcGcXUdD9ybczT60oTZoPyQJ8NQsbbxQ/DjqwHkqb0V/hXm7u
AC5/r0xD90csKo6/TlySkGcxh6KWEBNSom/u1p085gy3wceHzF6AgvRc7J0ijSlM381uOVSaWu/f
G4YawS/rWpK3aeCzD24lvQ1oZiblxieGSzVSf9e0kmgrFy44n3IRXzMo/SmFCLuoHzPjxD5NsTmi
MEFgqQrWZaLjzpWg5sRgHXzBWpaoh1UQcxqJ5M6idr7ht59/bgp2sxUlG/HjEQE2z2Xo7FEFGqbE
bIZykB3shbvl9aVyFDxVamphYfmIwX4y3AT3eOsnOOQwK8Y3r4jBwChbZveZB07t48582eHztyuw
NOSDz2ET2ulDzH3HT4/WSqC7d3h5tLUevIAvFuGfLGPKzvVoHCSfJqupfsxwe+VADk50c4IcQU92
5TVWSAXNYHxxvvIQB6lyUoZi/lKfDRBc+b9KowDTHDaRCLmi9Dt7UqEvihiD9leVyrgJlN8rl42W
gEIPkZznNzHgvB1PCZ5GFx/bonWFCJ4aNbqkyyO3FGmcDw4zEFUpZKjaJzEWyzhmiFvGBef3Qhpw
84P+HLeItl349dlzg9+Gq8JYHl/Xa9lqy9qhq9dWBwU17WchCz/J/jZqu9zj7fxV/PaFfitxBbla
PaqlqmC4h2jbGeaVsEPX2ecvzVsWo1Oa8qi1TzWFwzxboxT36KiWlLeFse3nHrfviPSvjJEsmcw7
LfNshms59YEpdojhayq0RvrWHD5USvBTyaYwXj9uC1WAYGtrsoUSnIHfon3avIryROws3F0rIDJr
J9L0NO0pR50nTwoJWVu7oX7YheASTsHZYHoPr3Da0txmDXQ/B+rAcrzSzK3IlyNEidO3BH2N2T8I
vekevso9YTTIt5Oh6HJEYV93PlgSr2r2YfAHvwYveJf0d/Tby8tcPfgTUIAVM10/HSgFbK9gKlfY
Un6suUhibwDgj8uUxpyWhyghWA4pu90CFFof+bbLZISRVWsZSDOvbAb7aQLNF22zHaFqFA24Lllx
iJljCdLJe4kcaE0/JICeEZlV6F6uvdX5683sDXWIEiZkkYQaGWflIceYjlS32+pKneWfFtK2iXY0
fo+v6N27C3GP9aHX7WjIs9RLWy+A9xfzh/BW6akbGvsZGVQMOmGNF0E/isU184irhx0vOgdXKeU+
a3tgHm1NSGfnRYg2vl0oaCakOOV+q7xOLpxMJRbT80DTmz1Jrknad57ltn2YDQdMPXg2VGOysoCg
rm1+5DuhXQW95AT1J3Bid07IlMrm2414tIMLJTcm1duv7IRSUXGXXKvgP3lkFxgknqivwoQEXA8p
9z/+wkABjzwKuD9P2a9ZjJI9M/e9fF6xU21r4Ovx1iJ0KuY/dNr9ai54Aj4j1F3g4d2XQGWQIisA
+O8HshfAAsizTA7Myu5mM6JM3YP5+Rc6LN7waWTye4AS85+QJMmMtrvzR27OWHyCWLC1kQVgUkog
LzIwD6DZBF2MWyK+iN2TW1xhabJaBP99GCPTIYZoXPZx0GRLRHdwgvEXj6R2+ZKmoyg9tnmijczS
BbO+TsEacE9fGUuIsD8EI4bvpeK13eawioqc/Vc6sBYPNbb1ZvIiv9uCeFVRR+AbE6Bo7NwMyhcd
4yUX+IIfFiRJwxLRWySKEC9CF7vIsLmhjJaHxcWZEeAPo6J74/x93scTAmz8RKy+Nmnll0cUpBSf
4kyZhYiyMmTF3Tsan0uhSx6giblzs+BeY9OO9Hnis6VxEP8ZhZa2phNeEwt157fZ0ymbCOvxAzCi
fvTvRFfi6skoOiSWcfU8uiy87CChwz00Nu0z3smgq5W5VkFFF1NV+wXyfp0N7nA2RqHdaFcf5zZ+
cLgjz+p241kdvTuWNVhJaS2+PM9JEcWLpbQxiB/Q55ARRoTLeurBdVY0vXX9xDYa/NQ64Nrr+hNa
PlE4uGAOj0n8a9NOfZ+t2mGjgK1eQDRfTuFqqVphyVdEaHbJUO77aV0xDrp5jU4u8SlYz8O829IH
GAPxyoK+U/rQyE3DCNkMrRzVQN4OBgfzSJ/2s6WTj3vZ1xeJyMPVzr+BRH2mqVpkWQdsUZw0eSWT
cIWIY5IYNA3Gv6SDl89ZzRh+M7OXLPtGS7fvO1UQ6sxFSpwWXHN6phXVJcbcSZefdYtJlLqouifA
Z+dA4DffQ/7evOcZp3QVlr0wMGKpwB16E9bznf81fh93gw0SIdf82OK6YO2xi/ZKd3ejvjzENBcm
P76lNZS/qPKxddRyIYXZFyc8/Iosh7iIAKYPdpc5AUw1ktA7eTi3jxyB1UgX6I9yJxcRlySLYs2C
GLBMHsutYcCiPhVW5G87Udp3mEda/k7PqfCMw0NaMoEmfMd7j2T/fB/QH9erLrjdxZnSqC4/hUqh
ESqUGEFngiN10jpUOj214T0WceDRePDudTI2Kw83hdK9YarxYdD9Bs57vFXBnVX4Sa2puG1/3yW1
b51oAq4Q79BU6uD9uAs9ylI6YjI6PxaKKoxKA7c143+Zv1gYxLtdOUWV6U7WMc0n5Q2mdzIaTTkZ
TSAF2NqCUhHJtiExU0Lvhzzv9+7sboAFyfS2Z96Wg/3Ka9DoWGxr0syOPd8CgTQ9M0uKDbqSqaD9
zNfQsb14wXCZKKe34o7uBP7oBr8HLIUPvPBqEbhr8ksVEG6uu5nzgSsg3Dq9qowq+fFE+NxSpClc
7jHRTT6T3G8l0EdBrpFUTO9gbiYLDdlqhuysiLOPUcw6FXBlrfDDqKb8/JFweNMWZJWY+Qv+ESbM
Pxi4CzVfmAFTFiUWziq4TaBpM1iHmTRrnozlDyLa+/zQyh4REvmTTIwgcuNKdaFEr82R5JndauiY
LRXNO4pofHTBfF6AKfj43WOevTvKWRw8hDJknVKB9egSEsPu6OrNHZXZ9v/JLF677TuIwtwNXUBg
VywA7nOZi4kFMth6hkslymygKyIin50MtCvIv4SH1vXMPQscSwMG3IQNahhMVMG6Ra5VjW2FGDjk
P6rxdAsulsTf2sNU1RfkbEeZwL7m+8YU28NITi6d9JAMGzPaIgnZuGtRfMNTOvtbCryDnsKHo5EG
I3sF5PJAtJYD3KMZl+Qzl8aHtCKKt+KPxYMyg5mBEcWQqhBSazne/Zpxu+pWbmiyhBwXwKKPnKVO
pTGddJNwkYPrQjSeWL3KWc3KIKYLdpqLHUccZmKH+lOjYUA0DLg36KkUa0Y5iI+QkZIALWuxiGDU
ZvmMy1RMEIGqD8HopZhNURvcpTVakRnhnKqDMfkpY2qqwodqT01CsV2TafKPKqLy9Jw0mFLlq5a6
1DrQu3x9+sxrS++aUMNobvt8Rd7BSqur1tTubqbQUWxiv1O3DcOk49oiTzjhItZ72wzr6yE/Ctjd
KZv8A/qErEnmax4724D7LcEI/VsrS9PwCoBpESUwhc7jmZH6o2Xywka7K8Y3ojioZisyiY3X6181
Zzj06X2q8ME3O2cc7cR0E45TC4xOuwO/hj33IArYXnz7IXCFJDcoERnI6DaeimcrJyE/KUuHryhv
D2IkR7RDWY1NXwJXbjWOeH4Gxq+hx/0k8iieXyM66iV3ixhlxVVdDJ3xLb8nuoKbz+67jIjlbvZf
oQNxZ95DiOwOU2rUQacEtvxmnQOj0qppUBPyI/jSJg9Vqh6ZdNDgB1Z9Pz2Egt4oC6Eo2vPiA53y
40LUW9h38Ksv2fuO3iMtmKlhjH7Kx77veQXT23ynnFOpy3SkNbtMJriaMhGSMD4ldUyciJ5y2p8A
s2KGju17TK75Lj6Zqd/WsvxqCwJHVEYB55Vqbp4TfeHq/fxuIwJxySmLcHLmznP2pOirEO3s1KfT
jaccLIwRdVVdUReewNNLjMtlHBMC1JI4ZHpXPRTuCC9vvR9iRxJvQfvhuPzWXtc546BrhQMOFpw4
T3FYau9UZTRFlF2hcnUMCids2T4YwEQitDP6E+8m2FtVja5OI+5PByj2NBbq4wH7XdJW40QEWqfQ
DuQPEDQ9Hqu3K0koqHv03dI8j32csPRfDFT3gIfLSzFePIfF5MeDvR/70QTUXCRUys8ht0/8wURn
pkz0bwWnhIzDa9IvCIphPNq76xveL+EbAErnMgmCqvXCYh9sYkV8xaMXXnRD+nywkRU6UqxEVsDu
Wtt6PSc38UJ9doTyNjNdRiIW+7PR1pSYTk7f7J44qWyuBF4l62CoTXO+WwbbOXu0vNECJAoYEMhA
pmBWna19MZdA9FaXOBeRvnRVhX+8ROxxu5MJl2KpG8ZsTvFyG+ns63VuSPI11D46LcvUApox7TYR
gERETWvi4z7K/jbvANIIptYEC5lLzPT1h8nyPDJeSii4EP/85YaF0CkQuXPMkCDaJCGtraxYZtGY
OVK7MC2YBqfwPC4nsiVUhLmtHL+3SyaCTd9ufng+EFLMUvMsraEbB1C1QNecEDnolhoOwZV6TS0O
it09czcWzM9e0sG51NARZZnVnG2h51LRm4FA0FV4ufJrH+bzvhwp7KU2L0DT5nLaFvHOs3UtZNuX
D8a/X/eLwHF4kEtLpgOtmV7mkYBd5NsLsNuKdgnkGvSMIWJnORHE85PsvYM3MctXOqSE74yqvMD2
2uBbOTXG9cI+sjhNdn9nMHGrItZuOX153mhuVDKD9QxM2O5ZicmKuv37GL8M8D7BcRYYCI9GYXsv
msDXVsKJEQWdM6TPOtO5Tn70DDW0mIb88C1bK1N+oeSKoVBKP93skE8lXo4mr7iVRW4hC+hkxYoG
v5DT3iM4C7pffcSiBwsFxH7RTDfpQFpPN5nbbW4c7MwnKkABlROalta/CanALIJo/qpliRvN3Q5M
9Pe/NzCIs2thh3GEJYOcU+y2MUfkj9Ux4n0UUsAyJ/25LSgCIoewF86CrjbLiSZyTXbFs2hXbFQD
4IUCeVFv0BnD8NN0D0RPXUxqU/99nh4wHPJdwjDOlfoe8UtJfNQV5yN9+Bin0DIp1rVnFHc7lL4g
PGYY547NPEExhbfuLN7aAWIwNQEVMbExyT9VvIWcjNB7jYNyq0kF0hHrgZ49yAJWZoHAXJsUShKk
VkaXibJyvcP4VQyIqBt+wrYUdU6wAGguKZBAx4ZpE3GFERB8vgfL8NBjWK7bI7HJnzBi309v2IbO
HaVX1xZ1iVgYlULslSmdYYBO6+AxGRUNifXfjAjHH3w3MIjmbkINeILllrfel2rebQbLuOzTk/Gz
C0xg8AVj1/hsIsjK7rGl706E05KNEactyxFeHOkV2ECe++qazz0dKP6bT8d6lnC1Ot1LD+v+TKxX
ifU+EaYWifviqoozXx/OoUb8gOpGHDILIwvO9obvSSx/f8tZ9fEwhPcybxXi7PRa71MblTphVr8E
d09zZIwvAz65pkTGaDWf7/EO1Gyr+FTY70wnAcQxPEKi6gPmd0gOp+E5K4e7xn3xtNqzkWP0V1wu
2nSRScz2i7Y+49/glTbXfXKPxjYEmq5mam7uKnrZZB8W6l05NI+Riqnsfo+ioz87pkHEjkxtsAXg
r53YSKM/P+ul5CckFIEHcc5V7mRYHkJCRrqdiJ4ESayp8bfsdKbGfvfXEbKq6RHaxTwOfXSJMtBF
/FgXu6w4ReEl5hpaiXYoeQFzaBG2bEZhyCZKba++QmtSgA8/594hDPykNLs7n38EFZbMKbBRImIm
rBPUXQPAwaY+3sj9Qsu1l8ga6KusJ8JrkwakRZz1Fn+XnN08zgDfF+f8MIc+0kyv8ioYQOyKhkx3
QKwo5SAmnAVAMsZabsuu64ZNIapdERwRFTJF9qJqCv+SfzZxduDj2ayhNYlWoZDMSjExAzZkGR0D
a251mi+gH2MZ7Gf80RsGJwbwjAFgThuJ9N/Wb+De/5omuoyRHaxYSpU/PUsy/l7l+DuLpqMSqmyI
EY9cwiE5OpuVv7hq3OSAvpzK4N2Cy2ijUMAmkwZdmybC/bVM0MWddhyQHnRui7zWefSo4/Y0poWS
0vR+aF3QfDGL3eOV3KZufgHHGWxgUhMuz1DCO5uhFjHJfpKXxdiJPna0V8ZU5BPvkUWbVigUnnXk
E23gHbWuRRll71iH3a017NIYMfZRDnd7iJjCQ7P7anxy8pByzEZhqXp+HTiqZa7nlfjOLm3NwALS
daMmZBh4X9CpX1elzaSnwyeLhEpodJK8xa0X74KFs8GG6i8DhHBOWlF45tCDKgwwj0M1/ntqcl8w
MK8Rd/9evq+YfoL+QmH2kT7H6PwOsdox/gMvP39daC5aK5UP6sbRdnqQJaWC1BN0l92sqdyYJ41W
7e9ACW8a4jv/MjzM5dkpHvg2xVFhjBjpiWKnXI7Dax9Obb/y2SQzrJalVjTZRobvQFu0DoHvLGvR
JgwMC7lZHnNXJnrbR404/r42zYw5teN+IBnhsK01p/S2KNeqJBMrtHDeVwZbrbQYJGSX0ISNPGsF
FeTfFua8j7VtqCNEGF0GawfBfuzE2hMo80KJJrm3ToJZ8XdD3G8izqSE1W38TGXT8o4Cfb++o0+J
LgCAq/bYdEe1bPJowx5RBKpQk5rn12XBjAPX7mvn+eB1oulF4wgZ8oc7tXXIQNcWMAoDorNXUGg9
Nb49h1EP+eA1VNZh5NePdB0SDSVfwnNQopqlJu+JCZOJMSRR8eoHXs+dUvbRM4IoC/7dq428A8tL
q2p0s/FnTsX5GmyDswGq/FvbvxpMLijg+Ee95/pBeC6WFO3hJraJnK9zR2pA2zFz/4QW1/pepL59
IlstFi4HfRdvGxNiT1B2RpscJku2mC9ES1EQCmJH+xVogezpKuxX6xyUdhf/WsRbZnQRym2Xzbxy
xwPhJQZQVKQ6QrENBELiEkJbLpHicuOeCoXIbjN+72mIgSOrpE9abKLFCntx9tCy578n/wI7JUvs
0iod78ahBlA09h99s5ue6Z4TYjNDx8wnCRz/Ifi8LF6rJsZq0B82caKNkdAjVONIBBobx5JauKQ2
MmUuWkQfVW67uJ1VbhyYyQ6DotbjdffhY5C1D3kK6XebBhXOh7kEaqIu5Ahvsq6iq3h0QyNe8Y4C
yXPARUEBW5a0yVppWNhKPhusKWM0KbEFEOvz88812XTfUTmL7fp2iIuOCnYdZO1dYVsoPyZjqMGf
6+EncYIgdTtLKFUVmjL+w2CrCUNIjl7jo2ezX6tVpXgeT4v8lgnmuLRVhfS5Wg6mhNED37NWGyOZ
mZVF9p82L8I3DOyq7QT+v8GrFxHHxId6qicGRbE+WR62Idrli/5SBi7VCfVQy1mdHYeXGiO0VsLv
0VAHIjrhjItzlakRndZOJZvgXYbLsRPKRiCziktGSc1T84WcoZ/haocCJYBDEQufvFmTqvFi7WOf
XvWKdVrQbGeXQuteyE20Yi1MtbDEYhYyCj9RGdV0Ny4EzjS4rll3HC8dt2AqbQ+xCU8+QTMj1jLz
VGfKs7gmGVKzIZnocAB47E7nkITl8bsXN4A6BIyClFSNZftAXJqo0gOaljVPxWqOBYNG3cnBNfAK
ns6owyo37XmzlcIN/crnoguvJOm4141tzyx4UINzbho9AHSA+ex67hY24MHZQoXu+JrSd0vxKEkx
x98oONabjwziDwmNEP6woErTYyY9TdnyFBtvzC0+oYjexgHS1XmL170PPeJVTTSNcZ39gjNk1Np9
rE0cs+u/VsIZ94KX5Yxo6rWT7sVRhnKv/bDjwgvHEj04/yn0PTIjrHnT19yzo05p77Ln5pNd/xiH
+sE+ghqQzFdxvxkjjfOkxXNO36RjB2x8ZR86oNj7p7PjDD7c3YHfP91MT5lBh0YS7c0x++Sgeyt4
ZY3nRcaq5zZc+a/JIDW73yWrFgz9MDvD1jg9mSzGFxG07i06tBhnZ1bVchxOXwwNPrTNZZDgZmyY
vAv4MW1yEgW3l1WBwDt/M0ZStT4+7Zcfk9SZg82dLH4enQv1KIujjTosb6Rrk3hNjdyaGwlXOFBJ
Rj1LXv8mN/ezaDQwJvusk3w+VEHnbrNqKT5y1YfIDXn67m6BUewvHbRLESLC1d6/UyAWwm5lAxt4
fUotGpIGFA2tXNvP280PyGbOPPwxf4m7koBIUN9zQ/LnDkpmRcOVnnwalsoqFEIc8hToKyAhV2vf
WB2H+nz8Rw4JikTFatZ7u3Tv/WhDMjtWupTgCUweAenaD72+1f4YnZrvAdksp4Bg0JrBYXsceBpL
DsoUrLPmXcnHLZB3pBoDis0zU8xh92YIMTN/su7MK174rqyIpvHwTkAOexN3B4mHAPaTOBHaLB6i
do4y6mq36bwXKEB12LbPXtHVP6YBuvu3tZclLi75ZGJ/b1zUE7EiivAAaGYm2DGZufqvf4NcYLSs
U3KBWd5J5lU1LjrqaAgDDIMlADecMzxz+t0rQE/1Vyz1M0zb6cSwNXEYRo9JBbSIx96/6E4LRYG/
4NEpwdZRWnVX+HcHVdj+WTlQSHMcIkgBfrCroOWpFNBprKxgjSyN42QhuZva+HxApM9qSpANhC/m
e4PxalrtW0lvZCxiKLgEbZzgDu63tWDNC7h8IMKWSOWmqFvqo7B5ESGQYTHEGP5upjXMLsCB6Bp6
hEo9H6srUfXWaOjEheq8hv5x0vKXO+Z3Zku16ZnLb1XKrSzet2mYDiXO+CoipLt3yi6jsKBP0rNx
P4XEUVj6ZolXrzyfKulvMVCGNvntPfn4s0MsnTZKN4MohJMlepJCPxZAU8RKSyG5ubeOONnWcW7H
qJg/DzrbIrAbSIv5D5gY0mjQjLowctdayLWo9lA4Y6WPk602xWBmhPb8tE41O9VyYlxT/MDX3fvZ
Dmh2N2zhImnjssTxrXbqWtKEEcecYeNjp470xn8OSZAGdkdVj0OynahEzQCx+SHoyIO+7W4M5dpG
YLgfcAUN4zH1wmhiIN9YRVLCvhM7B/qUqcEFQ8Vguowzla3KKbzYrZ2d1YROErx1Z0q9ohU3jAm1
r36f7gvx+0BWr8/QfXwYTNOjhBmgx4ZAZs0ZhRBitNrDCwWXTieGXjZ3vMuAyqlPrG9n1U7w1yFX
nLtSdc6VUuoddUzZbZC9dJu0Ba5RoKNqA5RZ0LRcReU+PASGWRAkG8+PNUMhGf5VZa6tKOKEsWNQ
j0qO1KAkndZIB4ypkDl2TAmgZhiI+a8CoH34IcC3sluVTxeotb/JvErbvr8jfyGjDJYhFbZfe9Km
g84iqCDTWF0DYxOViTczVgnTVIpk9iyySfseO/XtNonPeTUqZnNTWOAF+kBln0yFCGeaZcl93/qs
wiEnumfd/RvNaXMeuA33rTULk6vYVXfsC6LRWxgrz0leR3RP6rOkO1Uh5wl4Mcu2lMp4VCmVIpez
D/mqc1XfSFzaALl2I5XWq8tCrOJkrqfMMIHWR1lzwO6figlKwtCE1ZB9OonaJTJHjv65sZ4sSuVB
senvOwNy7ZByg+Wm9HLi+/mToeQ7ZOIwU1PxdqZ4MvvRuIe+jCmNr4UeFQ0qPbN7mw/qZgs67/Em
H/5pm16nj/4PNqHJVPWZ4/W3UECp87sml1LEJpeT/2Qv5j1k5JNirPmSwEF8dgrZWWV5z4e0URDB
uYGPaqwowv0urn6kbd+Ay4K8PNRCnEy7rlb1cG2LjZ6ReccKk3WyOJvNLXc14226hQSkReSEx+8r
PlFg9f/E3vFxQRJd5lMzCI48Y2NW1ytdlx8G/9VgZYq4RBBf+PfxfXSCCgCDjHECuzcAqGvov1vw
9l9o6HQt2Jg/acjS4F/Dxi7YDi4XyDYD77mtiM3T7qWwBUS8Tk1knrTineC2trlS25YRSHlsXGEa
Udo+E++HV+eOyavoAuFffHhYmzt8kq2w/72viqyTHyf6Gi8Flxom7RZdhjWoih/p86VPiE+Uu5c8
YLPWGCQ0bI4zR/I2dulc3G2ViUfbhfIkJOHlJvgItmgcZ6ggFnHrmfMzmBz5kXfMik4+zusHJgJK
8ODJm1s/JPYLTbRsBK4P38Pc2Me46Tgrdik6wGT7EhcIf7s9qnZkQClsMGUqpiWdICuLUs09OZGI
74CR2f0nnuplvm8/UNOkPzVtElVMXPPMZ2EuFb0k69lwqCLMNC935xpPQAoIHmI03nFNS4hYRPab
gx409i/3FrqCfsvr+eU5ZFFg9xwMZNs7AEQr+yVxPXFmRIC01PbSKE/GKPqxuH9U7TTGhQAxu01B
QHuJ3uu4TDDxYtJSeh84RLYPhqGOIDlWDqqbJHY8oFInXASkOMrkE6mBxhT9TDn7ZYCQzIj2CIku
/oWoabz99qHzuCGNwQIw1KhrCN+lmQhrHIzRYHZMP/E8AFOTmGhkzA5xNk/CpuWKNNcyyevTvA4z
shaqrOcYfnpWCjaSt7mgJ4D5T03GibPiDCGInxxt7i6CSvm7ZjfH8iafF7HN9T7KZNhFpOiekAsT
pZP+31KYM3W+DxL/eP9EpCIEn6dbsnSiPNWdgwKfTkACeZMso4D+5PX1R+NCyY4RCiFbKlqBC4lf
31NPBhI3Z+nLIy66ZkK/orWSgBTgDXvdWAM/lGxenqgn3v+J5XDiobrpv2+iv8wEwqE8CJF9tVoW
qkepL27JnJ6Pa5RzX7+4iMPZs42mRcbFvx4LDk/V6vXoIpZwcdrBPM0U6SExc4ux/+UK3Rf/JCRH
zMf6yXS4XqMRy+uTjaXEDdrOHBJYYyKHq+XZaREDXM2Vdy9LmCIUa0CtaY2W7AbcAQypCLZo4CEs
FN5ZGgLSXJ/UBorjbaZGaprP9yW7vzwtXLIr4cdw29oCicf7kdBaYfAeQXymBujFBGwIgoltj7le
gNIzVcpdCETXLpiPJ5g+xq2BNK6NEZNVSETnRzumcysgbIlqReaDl2Luux3t9OdZKMJGKH8MXRq1
Bc+IDkOQMZQxlxy0g8Jdm1o1PORWOmTfV2slHJwu1mNZz+0E+cDM84aE3s/RID+Umj+/uj53Oyk+
fbef6i3MyozhBVCN4Pa37rGdiA4PazZ+Y/GA9RDNjtDmRF1hkYhMgN/mp37iPKUr7Oh8geUSag2z
F/0pBK9400s/wMG3SQTCbvMAIFrkqXRlBQyn6VLVkNkaXOdPegmISL51i6vK4ybNCxBYTWKaFCgy
5Xx18ch2H3k0zKrql/gMfT6f8RTvZh7IeZTmgeR0Eb1RBi6CyRfRYf6OUxDUgQ7ETQTInMFtEN8P
ZsQammt7GjXv2A6l2tpwOPdZM1t5AdcyP09zLd5kqhBAG3RnGk9chmU5QU7QtDWono3x0atVGa7b
rjSD/SIqAzGhM5vjF4l3kgod8azvcoowaapBT/vKguuKO9BwKS/6Ry3n/16HkXmCN5Uk56INvfFX
DwdjhJXTpUZaHi3JgWz8rV3FRuPEzNEHLbYcvy6z59/4oU4vD+tj/k9RhcBcorTVxirfmjdwlRlp
2tt0BP4kouRXQS1dW3xbhtl13KChHPSIqjvef4TAWtCq8G2f8DfDveHCx4eGkjw7LTualkKn8mtm
MJTqBd7Ey5GjG+OpKXFsMI3FhLCDR8VCTNUrS9937xP4B25wr6s9K+kRjx8SW5BrZTBHJJvzAq0D
T5UqwNR4CjGNFBtFWzSNDrSi+dv3PcaTIsM3kKIgenpGPTWb9+iZLVyCwzvjz8v7tYsCxWoxcuRp
fw5qUkUyoXp7zadc1Rkm42soh5hMCibTPok65yDXYrt37z5Iyqm4pxKuOvFXp1jkWy9JPTZBTAGb
iqaJ8OufKBoMAhqN56azZ/XJPjZk6PVPSqDoCwUvSXr7eQpaz5Y10q4MDpGAsXPgIt7+ixgRl4ok
G3wnvurrZOAVgataiVAIDjcUTvsEbFKl3czjdqdDO2IAxp7v7bda8jJqag3TMf9rKVhegPR1+4kz
zBbEwwPzculR8/zhK8eB96pD8VVrCIy5BZ8272AsPMLO/vj/oZQEOLK1/Z6EiWi1Bp9qKn5Tm0qa
UvV8/2rd7fUfsFWo6s+qGQDKARlCzc2ZgmmkstHkriCzFaVsUlk1JuGxnML87eqs/reOhOpu+HX1
SWI6tTDXh3ReB+LjMFKRtZ85Qdjw24HqyvVhkMju2V/WaxCv4z7YxRaQU0ut2dQBSh+DrOVbOBxK
zEnGjmmVIic3AdaBfwYj2hADULBM0eu9pRJWLpl98nJCSLO6iOXeTihMOt6+CMxwoThKWiFBrwZJ
zFg2m5GTrrBdRU6frl2Eivu6BVA8LB+ERJSYhtx1a6tHujANfB/H+gu38FA5bg+0/GVY5dlQ+faz
PX8PFc8JeypQbiR3PXY9ZVOKKTkuxmvluH10qHgszu13p5sw8Y5ruqXYkI/9IqratY1wvxNEXbxf
oyUHaMoGLNl0yHjC4+Yp3ciB3C3BBveTGK4jNrr/W09m6oubhyFthCBWF/omD/WfWGX2Pyiju0gd
Hdeuo0ypt3eTm9xSOfc7wlJYoas+zLW419+9LujSmbUQCfdvYthl/vKfTjfKgTRjUDE9VPDYJMrq
gSYLopTXBB8dnAQUaqapyDbLtWxsu5siFfO5gUre3jNX7pme/VNc+VNqLxhg2Wls4q3Rfp0Zrlcr
gkEpPYh0hjfhSLsRX/eSHwIl2DDlXAf3t8QrvdmZkrQvYLGr+wMqCHQ3jFKmeOcqJuZgkjUu0LI1
xMJRb8B3y1zoaLlRlWLZfhw9JWVKLpNiFG93+/Qa+S8BI2TlLQtLQrh9Le/zJgz5nt6dXHqd1HQG
SFZEne5lYEjg7T0jG8J6Fen4D5FV/SPF3ZU508IORqmwJ8c5VCQAHZCpwcv99lydMGYtuf4m8hhJ
XU3r2iW3E/D1DTrve/4zXH1lP4ndtOa8l9Fl2ZsPyS6fZBSG+1WbMUGh668hLm41cLdJ7/d0L/+L
iBhWse+LC+5uAmZtEI2ycCzIzVus/KyYhThMeRYmTTyYvHhnUvXv7XGowYNaPccnj9Mh95dS348Z
5QZp50FvY1AOnfER/58DP7Pgzixtt6R8P/SFuYFfYxCdrt6GM2eCJDmEphIyObGeMuOVuAcjJt7t
RbRJQfRLidp2BFUI6xt6gcMtWFNB8ot5S9DWgDWwwAqrFHip6F4m6U9trqhP+FExOW0gAR75pikn
wGCtumLABcwBOGbExOeTUwkcd/2Er77j7JSqGV/gIyBEXQV8QaLmyqWyw56h4BiPKeOpuhe6b06H
9otQ2RKyPJzeHOtupRWxnSLx7P9Xtsl123zebP8JOhUMI4M+ypWvzDC+/NTR7URTQaVZCXOnM2hW
aaL9rFIEnsjBjrSE1H6+SDI50lEsZD79fdZuaG5ARHMJMgIsvpfhG9VX2inN6SbOfHVE6ayg6Amg
dTR8fryOBmxKxJZYvnZu8mf2EffhtWRxJv/jK2AikmoDm/DPAEQTu4cziz6AJdgKqj7nk9z5ITbW
Q6HxFV3qM2mxQOETDDjmJ3yddNvlY6AiB+FlhekmtA8ZhxfuzW+Is0UUzlmBpA0hJ+3S8kojwMlV
ABzkoD0H4jb1TQQkdH4ZE5t8lR75c8Frzkgqeu0EKlc4cRMVSeMTFdh6DzupI3FjeTyqNrvojKVV
wTJQfBvL/X7fJIilI1Do6l2OQJ3xkDt0q0/5Lcs5K+bmDGlp015dJ4lQFRk1cXkJTUJsB9vgXwJ4
PtHKjxtnjfCs32wS8SGKP3Mc8XlWE4FxrighaGrfG21+ozbbanujEaSAPJ/UhePRdPpTLByqyBh7
rJyEArcgoZhe/+PN8i/XQ0ojFclSrLnv8zoMGTIDZzEwi8fSOOE3hNWlmvK3non71vU4hb+I6EHI
cNuVykDDTsw4rN+rXnfIPgBJ1iiIiv/3uTboGxPFc7LOuTIXAZuV6EPg3kyVy5cJpeNPx0pNssHa
D8N0flJNVVNszHKJOy2opw4obCK+Rj0ikrix6y2wGMIDGqc7OFxqmzdxR3GPuprPaVSZ6CKzDIds
fQHfdba+EyamxtA9FhBiv8dG0BmWHmwKhU//SQKEekoDYEfkYzukdRiZNE3nfi65Sl+pAQOI2d9L
orjU+pNuOcnmKHnWHFI9DJoyAE/B804MkIsUOrnmvCkjmokd9gOki2SIG68ICT5AyjUGeAdzo9l7
Uur9OcmlZ/oVyhD2QO+n90+o/14xg2ZsbOzFtn2kwIfP4XZEDLe/JNTDioQY/In32f53+UAd5xBe
F9AB1bfUvAm5OcB+GljeztJbEC+jlEOGzfxSDcLtMV9kS0qNwLt7AYWjdzirZ4yeD8RYnHDKxm/I
nMnhSQkg05qdLSGHtLuj4OxO0Ud6FpJ65OJSu6EC5qEMSZ5+qcAbI8pRaKDN7sAlWJ3XHG60fDwD
MdWV3jozidFNObkLw8dEkrKOX71AONw9aSXoKfB0R8GlY4+sEIfHAUu1WhDmYff7RIf+zP/t1Udk
f8H9WYw8eXOJ3WfEzs4ms+SvcKJ1xl8JOQKAOF086H9WuberI/OuiBngOsLJt8BQQHDJkGH7xCNd
+D/JLYYh893LyRH6wGiMa/274IYT/Ob+6rRS/+jlG7m3g5ICEXu+wWg6cPcaZY98fszjcemS6RoP
OYVH5Df+sFsvbwbnDlQizJwjXchxmptA0uMuoCstKbDbCZ/EOKBjO38Kxc5fnLs4V1mjB5m6XTUk
WXf403pkTl96FEbI+hAduCPjVmFcEax8I8jzVU58fvt94DaphB577IABag90DFxym1ludBLgPmWR
3D5JD0rYlhWSK5s92JJRdWp8x/7D+WPDXz0J7rMooArqFqN3mSWFStKJU9qfjOm9kInwRkk/uuOk
XKx+bAxipeyrl1SwzFYGNG/Fl0EnQ5f516Kfpulw6DOsrD0fWx6Qla16DsmObv4GHe/dWp90UqJ7
L4s1/alLKSoCIRKDNybbOeytIOZoNsM9hdeetK+GqZ4ZvYgtYlgHV5QvxsFxFtuF4+y1l/YtFp+0
6y9EobtBzPoX1ydiuDR8T4wAey0tqyb27OY5XmAgUFLAwJOxzm2cFaHQZIRhzr28NzWdbox1lFUt
yYH56CA26EuLvQYn3TedkaD8TeHs+YPYIA5eglnF/UK86GBoLmYw7C2W7yekNyPcfETHZcObRY0G
wxsRX2RYZ6jHTCl0Wq1IiHft1pMsgdmGATcvvdwAcsalHXeseBxYA8vNpcrju7jzT44g6nigtC0a
dRdq4Edi3ZmsCF/MX59SHHWfpuEAJYWdffJMRtpQ7k8qQryNdj3SMQzgMcnSQychDijGk4Tx6fYA
Xrd/QT2CsmhDsWv3BVrA8GcjVUL9VByH2rYZUWrNmzt1CLqPCqZp4uk276MdcR3kDELLvmJdBdDN
zKgucUpclLBBciiztmYsFPfQlb64L3ekJVI+F7FxQaeFXpkAEJg+dRJnoNL/91sNQPDS6mOjRyXd
rCr1s60Bz4BeLYGYAS43ZaJzfzzImyvox2u9nd4RTZbF1XwFjHvWSzllbPHX/ZsQjXyUoLPEaSwM
yBfYxi9zuyeW60GqjmNdrpPVXa7/D+JbyiBTkdE2wsW+38NHBCX5L1b19RSOI+bO4HYEPfvJKwbh
NtiOSwUFjaFUlMYpX10ZFvIZa8rGS3o+kNqxHMBBA3k7MFW4QWz/LUA1L7VOHWWBvIvZvYXm49uK
AL9JUwVBTLljhoJPX3EA2JNM5DujEkbbuczqvb6UxIUQ4n2Wj9yDkVFUDr/qtzWd0y/fcGCITxVC
GDSlk2ZA2Csy3dsWJ/bXeSKkXsrVLL3EsvnePkSAYsMDK5/vg+iLQWqIHkbOfsCFGilAv8OnsSxu
Cqy0u0/sLHFcetyWxAt+2XjOV2OM22RZ44dVkZWjx0+FDvEOMJBmASHo3+c3YvrhuNDAwRUr4JvQ
V3iF0xKRn02tcmnV/XGNZv30rEJAGCjxa0m5nwN9k3qZxO9SVu5m5a210U6i7+nj8UEwyXf4gBLy
hol1v/NaQFesif3upPW2BZYrEW+vFfkJBkLXOcWXeQIumUN9vSHn3t6kFID2cgi5tLS1gyky8/Kn
wsezudT16CCoEgWhLEgaHZGx3fpywYDaM5KdkBNbTCnOPDSoYrKfMvp09hIeYGVuIqu+W3YaeMsu
MI6TnQG9W8ljsx2qa5fIuU4DzDdN1Om9nIMoGLNIFEcNtzqPqb+6qPZAESmB8iI1PVMB8MnOhbGt
DTbHlTs6Xx5MHvdDeVHdekiZ1t79vCod+RqwbuIhEXZFy8MdtxazbgDWsTHa7KA13CtgU+v0HQ+7
wBhxKJA8i1Djs53qaQQuppKpL96XMpiOkfxa0vUA4d5FsvUrcszm9v8zE2PUtgkQX9bt2s3tcN88
hM9ZMIFcCw2LY70XoAS985Y+JuqXYde+kKVAjp8jkgaf48j2mqbuSbXPBWQieSMlSpXIPe/s2iCL
UTch0aCxIk36Z5mc7CIEAcx/vTfd9dpN27nFpKX3kNWbjeJOHFnzvmFZD9Pbc1cLUH3qGeB6DHzM
Hhs/5tO6SMtMQS4Qj3rSjpHPfrbualiZGRx2m3j/vt/Tl000Q/vL0+E29wiA11lWp3RfaiZzUZhv
fKzcPc9iQREqP5NqVmJEfBcd+ObUf+xvrtsXE3D9JESVCoHQAR8e33S3Q+hHpeq/ICw2MSzoUaoB
XptOcyz0Ty/5Y5n/zyUTSQ8t5taU/ariq7tmrIUOMfGCgTyg78Ic1/pZpwqf+6MXvHFrg0rzkXER
rHOHdi+WS3EyK+cYvD/yLwPfvnGCKuuZDHkYT0YVyUtk2PFrS4dVOleAJXpEN3ZSIAR5J2+hyg50
x0QhPOT/eVeT6q4iu75CONUsoW2X6jrxNL9a2kUs8L16bQUDfWe6Z8Oy+co6xrMFbz83Q3trKJqI
jHbpnaoJ/5TWuH0HIGOI+kKBqy9wi8ZTC9e0g00IuyqiGVdms8wY1hAD/ynnF6u+fExMyb8fS0VJ
NLt6eszA7YtlXu9M+eZyKSxSeOOm6lJy68WILtZnnMD/9TFvByRZbkDF2JF8rgPuDnUbszzVPjl6
EsuZbaNpjuo+iv6Vy/mW/1QjEplJI/H3DwmUa1/J0twvY2UdyurzlwFzHLVAEIZ7XkX0IdyqSxiQ
7Ylkw99hxGn4XPeWEerEMnBEJYMaVFdCaQbo+EFytfdeL1oObPugdT9CcA1J/HR0Vlu28fDjRg5F
eC2MgQ32g0NNrd/fnL0gCRIDB/IfG9firIIhX+5SxfEpox7BtLCurRdIrk3g91HoNlyqUVQG2zgg
nuCt23fF+wdaOYZXOwdoIe89FI978BQbArJGYJTGYGsNMNuVSdljeHk71XWcz4HVSfrYfDDBlhW5
ytWJp/PiijaSAQqQokSqVKU5e3vBsXbJ6fjyo7rflftdiLQgyveLthsrhvYAtcYJs0tNdLO6a+cE
d5iC4lXuecpPC25VkZE3Y/wWB/hB/aR8pgnS6gHRzDT9Q5VoBE6wRnCV0s2ntdy5WwOE1k+1m5Xo
pdhCp1fenk6xFux081TEmE/4hagOwjaXpapVtZ7JXkhBvlAffD7UNHiG63GNBmueVZt0Ry8cV9Qt
FXjPO4zlK0R+Ob/Pvh8WZfQWnFwe61Itd4pBXYtcE4MyKNXydbDZf4RnHiYqaSnB+jh2zoaQ6Uaz
A/4v/4LUnXsa4JyLlLqigxI7kPOGMy4DWmV4f48lHNcESWVQ7IWEwGE6ThdlVEpvkT2GkF+wCuaS
wbY05E0O//k6Vai4kmBdPzeZd0tu7JQFUiZBXuetuaPrw1HYuG94akBxy1lQbBO8JkhZLTcoYIO4
lmtuZRMq7n+Y47oU1J3IJKBQOrnhfMsWx5XesInNTJybynUlmRopT5jJjLIE/T7fLW0nar8bbPuI
depmnSaLOg3O4h6ITMhUqsbyYqbVXbkThKqHUM+Zfh7B6CLjA4FgV8EWa9Jo1pGVD3IywXWFkNm1
x2MzLZHrBuSWysU3RovbCeq13SghclcS8YJyqabsohfLBMpItEm5ylxhdgmwEhCVoXj2J5rtZEXo
eYIymNHm+ZCFB/boq7jCh4dj4eoZdZGiFGrkxigM6RGVAOz7vhAegLExUuXZSfDQy7oaBoauHvKh
4OCmlLRvJ9+I1ybjhfnlgCxpRT9aJmlqamZb0QaIGYxWg7uJY9I+pb6aRnLiFHcozD8Lv92OjT7l
QYgb/dKXVMi4dYrk2Gfp6HMiKQcquOcKShe378vDlQaU8IBBDJu6pMi0TIAmCsEYejuFmNPbOqUI
oetCzEGJZ3pV3b4u3genmnvrKSQgUnJnRXpkN6bucMrqUgMKAw6u8p29n5dyJTTOWUUO8aQF5xvK
Z1IRx+TVriOyG/CCI9W9gmZxFxogMb0g3HdnmJv3JwUx0nDSpaR/jcI7gsg3XJJIKk5Ps6UVniOy
ErsuE6ZK7XppLRkm08aH3zeOdyj2xTuZZ08v3VTieWb44tUD+bO+j+2lMl8Cd1LPA4xNbnFIat26
sUbM26+/fZW1Sb7nekwX8FkKhbH5qyf7B+sBXk2r0UDa+6FqEzBweiLCAwVzVu9aI5gjKhR2Z/dj
IxFJMTb+3eQ7CTAZrXV1gWJYfwkw+kOf+jUrBHvO0rb3Z2I9Ym9SBs0sXjsTEsKGjIphVV9ueN09
fIrqO+JHWZhBJaAbgBJCtqK5mh6DQ+TK9p/8gRNYMSABriDv/7PDkyt7qlhRQIxlIJWSp+W+OUQ8
5sCPnE35+gdOf2f48HqSSCDgr+7FUvm7hs25uunEW/TecCaJGIWeN2x7iv479C0eAGvIf4UCnDde
jGse66NKJm/VfRUewajrpjLWXQbXz7DGh+816aSaT6/dCgXvDkBbWDSEnCAQlTKpS0oGdnl30ZUe
k+GlAiSmvw5yNFgwKLbpTZNu0h+kcIYzB9Lqpv1Tlozefv1eBkfibnmLiaBc4oDkxsTdTXQBQdsG
2+DY6uDsGBlBncXihoJTZjPNmIymJz1R4cJh6oggdGkYOUS6Q6+DgK94lu6z4w3dSM8s8rGb/tiU
v48wBok1H4w+WClupfDp6bxHfT3P06RVjDUtOZOUseNFOarnnMcWHU+rJ3jKgQJBHnVfb390K1PB
HNu9hPphf9HCAiiQlXATTGfOsIDqKAiRlPOLRB+AOfJTKwmLSmnaX0S9Hb8zy9BXhHTSKwAG/fG6
bfiiFchtCqJ4w60iBcNBhQfunbMb3lMUQlwZOGoUjvIuC8flpRKOBQx03PQd2QV4UHNfGjo6IPWK
CnWnANZnl404QGmFjIOzGY+k4LwUXed9lG0K6hX0siqWg2PYBWFQZtB854t1ygnuX9nXGXuKLArC
BAj3IEMszGfgbgS9+yBPoKN8m2VsirO5YAy8D9OAmJE1nCZSIyJn2zOMj5QjIbC6ctT7IWh5UHrM
55QFo9laPJdNC73R7a/G5E01zK+famiXKY+kLon5+heFE4YRKhfk+I638AaP/R0SThRKtVNMG+bM
d3iAmMo53nu5ctzj8p7CwpueXRuWgDH0D/+9mp/u32oCUWW5WXJLZjaaKpYELCwfEFNT3/6k10gr
EFs1EvfWHh2GTRb7xmGt9BGHE8t66rtl0VPvM11UjJhQLkkk+VqdufZunJA7uHPCLL7EJROJ0sLk
wjPKih5BiBX3+5NOh80e357hpQ/rGEYfTLpD9MWYJjHSehdsUhJ/0YMzowQOXcOrstd7vUUJF9ej
iov5P0nLeuxVisZoM5RKojzcEWZK+BU5RS4GGqf1xvG26U3o4x2IInwWLiJ8cKivHzl6nGvZpyNP
sfOnvaf8T0SNJfyGOfjCZMKAGcdtzrq5QIJ3+xoiTdAl+R/YCBVlV3ayTqKFhK8/FIlS0NicMPhS
/KaGuQy9nHVup3L0ZZbX18Daez/VIjOJX9jIbD3FSaJ/35UgUL6NXXSP4Jq+nPQFeLMt3BH8FuPq
owLv1FBqJOD4+ilNhL/Hvf7pW2bO+sqwNmXUDaBlOlGlz7UJxCYwbIdWMkeil188bn/Grycq4Z/y
FRlO//U1V58sRvS7HSjugjIAx9kZXEHjtqyTHidSe9UjqL1deJlxHWKOnUdsRs+OmA6xebARD5T4
nWiT48LOZ+lG2jvdRxMYX/Ebx978Ffkbk9sYVhVKGaNTGQiLIDefbyHTU4hF3qc9lMg3+CJH9NOY
d5zSVGq9M6du53ENLCeWTVmVCv7eAl8w35xS2U9hvpvDMsy9ocaDicD9pRoiLp8IOiGzq34x0J0G
LBlUeLcdNGJanuonAUPavT+WIBA+yU9NUwDyMfJ8b1R+DgHJtw2uX9HBBb8k+TbzeXYPE7oTteAi
zNvp6K19VPrVeAwVQm4xGWHYC5Xxzn0j7cekr9cBGC5WNOpNwnHIOnrZPirdrEkSGXS9OBE+6oUt
nSPpi2yjaZ7Yk36uUN+yBqwWvJOLdhODhCr2F+PS9qkDgWMtWcDNfzxIp8wVAlAWp8DkOrg3NN/V
APnPDesyevTsr81cEE9cxO77L2ImUrGI+UMMd8KX6dmM3+z1ZjCSsrpv+vSRKjT86/mfDz9CcZ4z
kog3J45JdXS1Gz3Ac+XmtHQMBuECyHdOxjLnVEdmjcQ8TU2riqzAh7iEUZwncfdO7JLvMsb0+wz+
gliIozHWL7b/4bP9FX8ksA35u/dSrCSyrLSHuACX6B9E5xGByKuRNvFzwrbyYgmVhqv59+T4pDbt
dPQN43XOujhFVR/EQGGjAop7g7kOL5BqtvdSvcRg/DExoRow16TgmBRpsWWskBK8BrPsuuGsRcoT
cIWRJ/FtwJjSjkTvB74wt1DLn/k3R3lGMyoF/+aYgRyM/8T/uWwyFnuWG0i2uqhxIFfRFk7Yy2+C
5L/uMZar8NE3soKrnlhIFXIY+L/OpNKOADsn5/11QT8Uydv42P72Hd/Ceu3k8162MtRNCkRHBcHK
OFL/wdVmbT+US48ddVnQZ2Lj5LN+TF/m2o/seC52dhD5MKqnyFoNxc3UGdVBnhTfbVhLEWdJLDP2
fgiZEa3ymGJQ8v9tHiUehLeIEYxxwRUrn0bksAs1g3hKzcNGzQnTpHDAkIx8OukwRGTYKtpav4rm
5QxL7VDyTI1T1/dpxFA1iUopR1Th7JCd4wPDCW+OPJIkN7hxFLIXwGwvBBOqo7QKCYElhp/l8bFD
ksUnBm1dGanfYpk5j5BJiGNHwsp02o4hx5MS38cFKf4b/s5JITTywU79ZUOR9fawRsCryW8gUk/k
ncYgBWJf4zu+YyzN53DZV+/kYpTvOiuOXzwLFbUuJVsEmru6xRFrubCvEQ5fJi5xZXKsrbZe9BL/
tC6m/WYE4K5DhlEyL4dxw05dT95FMkTg7m6dEPGBCvwhd8d0d6u8QHVrziWseMHWheyfiRdERC+i
rZ74h/drSJn6mmosYZ7VEwFf21XPQtjpVWcF0dc3BQ1XU000ei1G+Xxv1ZQ7qcM81CqGeBMa/ev1
LaiUj/DT1bC/TZJsd59pzthPlXWTIt1qdh6DoBVaoeB02I5zr+/bUKsbkAaNKsDMzLv/pFNlPxBh
QRf2IpH5vdi808zap1aMmngZicYLXBaHNCQZ7Up1XSCBhREXLaxyOqhMaWMTn9cHG5CpUsVTXF9c
TocCxsuDeI7GiHTTQ5EP75tiFcErRekCFdqPp01rAOvJyUsZIxNQpyNE+Cq1/vIKKE45KbWHcOj1
c90RSyO+bjhr69QwKQ2IVbf38Te0xTutrYybWPIYU0n7/1ssuoXv+6T33CPcIHRsdsTa4t3YZBTw
J2CQHTLa6Fx33Zhy0B9ZWhZvH5Wqy4RivRFsJAvtTZb/Qfe0y+cdL49RcnFRAq9ZejOMtS55FuLS
IDabz4U3FQMfGR/3Y6gcMCRqutbyYfu6g0TXBAN7y8cl/Ml8HXKdHmBKaAjbmuXMyb74vQXOOUp6
n+G+y7jnmK3TCiAjenQcIo6l8LeWYytDPevZ++Oc3iwDVflif6nnGcT4Y1n47MViteoFPbZ7YGeg
ZjXAf4I4Dcvi2omGyjhzqiPEETuzYv458cAciVZkOrxXLF2Izm+uQ9PPEVwLxwpXLXOWer0jGWKz
NyCE0PwZGiCc5B+D3HvQdJishRfQyjTpQ7+Ka69FKdUf7T8kfa23x51HT6S56/l2REZIwKoxAM9r
UlSfkKBQ4M5aVkddWIv1BE1GGygd2HN62mvAEUXyq6eWgXk4iAeZHtX6G+WsKmCkzKCdlVBUJYtr
mCm3c/vMgT+PovIuBZsXZ5cwmPCDT/oaggKEWV9GJHa4I3ZL1lxGMBnXybwhWn8GVoUnaZ6EKUDl
qn+xcGGCRDjEzFppwXhQwDUDGRMIK3FIzkH2zV/ZMZTMTXmQBMNCfcKfeEmJbg23syXn4AgCOzB9
Cx6kXcHFq5bcgYh0blWHIT0daHALn5oPqH88/OIHdm4Uy9O2OfQn1h9rhZdP11t1vDmUFVm0wB1G
Mo3Cr9UT8eBx7d39c9pl/rzESXi8Q9lICFB5qR104HrQBchjo1IzEDSaT8T1xkspO3BIQ1KfUxWz
QKq+U3D+B6iZZb+Sx7TV3h92lJpJ+PN3ix+VDmWlvDIxBa/M6Q0qv4oLVMvuNpU+vekH7Ub+dMUT
Ge3Vd5T0DssfNWkQKlyIPc+A85GfzX7GONVsZPW97CaXSneN5WxhRCzxWRhP69xFsoYnJpaI1Mpt
ORBMFdMLjmeHUCjxZVZBh21J4rfJjaCNTlWG783Zjiv0vJ9I6hjs/H0YcAsjNcGtg2/igYAydmHv
snoi5K2h5/bHR+hl4S0nsAtaeU/Q8bFokVKjpoEO/Ea9/GpAbk0FIqYtnPsAfRTDHsX7S0TQ0U9A
tHorz4N58U7fjn+EOEfzMw9muwkKYYalZM/IxN+De5dgGnRDiC1vLhcNOrzyl3e02nAgo1gd6XFb
IyfLYPr4DlMczy4DlM9XipY6fKNDDLjgkkawG9uYkB6snRyBJEUiqZPXtWDyY6WoUjc2oq9tJxPg
al70mvTZgAy11OdVgxacw6ALSr/Xlay53rTVysjMj/GGI2R90aPrwLqr7rLmTja7qA3uMxhuISJZ
M7qTZvHigoX/gx/h+zjOS8YZtmYRQodUAl/K3eeJYctkrgKb4/B8fRGkTCIzepdR6BVGlpWVL46L
9sfQ5CQIBH3lDOWRiNnTqIeKW+eKl8qeywKcRUQ3flLtbJ1G2TEX/b4lgaNiUwScqNeqdY63nsyy
8FqG+mW6+05CGtiN9RgehLCDsuPXta4T09ZqwvutpOW+1nehklHQG9UVuO34NSgNRKSK0Yzrewlr
qxdIEDlYycOxdbt/QNCQYZ99To0G5oTy7s8KCjbrUQI5baI3lRm8x8qMJ4S9fGqwYklJgFkRqIl9
Xlx/LSoeS9fvxumqxgxN+SDhbsU78IfGpOwrELkTisgO8PoU1XJbW9eHD8hUf8hINk8+aVoZvXfS
HaTd1Af7C5c+HFzdHMzmQHKO1Le+rKR/pnK/L80Wk2QxX7zBsbR35MoYErfjtZ3Ee9CUlgcHfDAs
AvK7grlWqCo/QvPoLQPwWkYI+Z5L0el746mFpCkxAjlrxflZZtv7/tERDYvuBIJVVnVUBdPHdiao
z4gpJs3aBuvI62eM4U1gox7BFEk7Sh5ldpE1Ei69cfrXhVeytpyf7zocdoIJys7HRIPN92z4qXN4
m/ODCu0Y7aNq4KOtGXGBq1UnjACUHva7NxsPJGx9+SCYcj6K+1Nra4iJ9gOFccN6Q0YUB3GNn9q3
5GuhbdqQRBR1TXsYtTyy+Tsif7LTVZTixeayhQHXsyr+hpnU9/mRY7VagUAmGccrijCnyq0DGpnw
veJflMTSlbd5gNKeQC2rR08IydBWJUoyN9sYlx2jPqmkEu5h1nTqGs+erPH+NwTH93T42U5adwKf
g4fHC78zm1Syn8e6wbVn8awACBugGt/7fp/IR/zY818lh0aQHRfKV5zdIKIhlKfRe/3CKW8Eb+D7
PgMbsmaR4eNXgbVEShC6Ly12aKtjozWuT+Zm7yRwwXm6m7yaZZHIk+kjHVVtm2CvR8EXubMCv2ga
jmVBLe/w/LaeOKKMJCACaffBZWrE8kNZamO0MFDI175CeY+/54Dr5Z0mwZ93WPCt1fnYE4PodHle
F3y0jaHg95sSre9+hyOsqMi9PTLQUTurxdguPsWwNYKTU54dfLAg3bMB6MjhqsA03SLZvOkzD2jv
Mn8sZl6NE2jd8gQXEkIaHNyiqvKEeDsnnrrReaVPakiGNo6SmFRz3QVw/kz+mNB49mlcfS4ge5M2
G6NGDIrCe6FTigjgDC02wTnMKbcTPT2TCnyHQHxHpt688saj6YsLM84Z++mtflfaili5tx65VDfk
75q0kkyMK1a8XHSy6EWvVan3CoZSmG3mLdZAeV+vkl4yYbJDKGdecJLnsVqi9Ibnn2m4VFygkWDZ
fMPL49RBKPQLO5fTonJbCvq4jOogDQH3OcFVvTu8QLx8UWbbe07uwFsHSTZB97+wp0rzgLW/4f/9
+goZmSgKQlC1CFKH/vseSJeRwAO2G8NMpGMOCCycNXe1jQj/yyfKCNbkvcl6CJU/Xj2UpHvOCIwn
wSq4VJztvNhGonRzZo4oEXBNnwZSA6Y0vD2gXNNJzWP5XwwmMZEaUZ4GczUCn6qU7cuJYoI8E2yp
7osjr1ta0lQa2pXgRAq55EpMlVAd+WoudFFkZujd4IG3pEJgmGWmxB8zMmPLzZW3vkjI696BXuKk
ah8EH8IqFObONwgAYh5PInqU832H760NJ4VXocAKuv66gQU5HwoGA55E47lCGuIAUtikf31gG7mm
FrONLUnL4RRoaL4faiFfW5MXED55r0Wl7KxJZWsQ4HeNGvXs9471MC9St5G0qQNZL7yMtb5DXBBI
8gzsF54IYhrVwCx2DGSqQFQGTyvAxG67I6L4cosDH0IYbS4sg+EaoMpb9Zw618pmXkfbv7UvwXYs
HlIbRlvUfaikWWewtRNuYS7u+/hqtne84Keh3BLXgdmmjh/Typ9y2q4WSWabxxVbK8llgRDvcqZ4
QCofZDQJ6cdAqRmXMbVcThi1mdexj+bVE/YhMJa3yAe0C/xTxrrXRcdafHn3fthtu2HnQhjT1kof
lt9t1tj0jGGuyPgs9ervUUP+AcfjXz4R9vhBdUbJJBZDWIwvr7PunM9bVOEww8OVsQG4TiKT+vgR
jEuO5YeaJHjiq0JLUc8B5hzLzLqEgdrNcWS7XyWq/29IpdlrJLKJx+G/9HEEdskkMZoTpdYZjBgh
WeSPekkr4ckN3Utrvbf1nzIpRnlWLyGNDTsnCx3sW+pCngt7YiqQLjhHiMUfEP8fincKIICyKBxx
zmuLRlHPFjXXsJcv9MiqFQQtSBhGVDx0RwMjpP2qFXCjkS0t5Xl6Ulg6Xpb96oWX/vKIoBZ19JNq
uU6tOf5EYhUml+q3i64I2ek1kJu39HLw10aA+nejzS1DqNkoAtlGRo8QlcA0nXv5fCNSWytHVKLD
aF+HV7gu2XAuR3mphhbGUM5qFbPLzoZl4avkz3gEhnEwdW8fp6q0nHw8Am+lAnKnQQYkQvBpTZ6p
Vwpdh1MzyccE/J+Lj6UPed9prBihPiDL+9DLFuZNKp0e/SwdybjH/kE6l9iJuKFaeimAFqI6Y5c7
dlbA5m3T4i07HBTqYcJtw4OLidfAXuhQl77qZjgeadUTwoVpQmyBLo22ho/DB1T3Raq+Q77F/Zy9
5hd3llQpKcyp+CxyFk/tMjd40HYv5/hy85Wz7TehoiGLvMXcdr0Ff+LWVmPxGDFYyUiBU1iEYaBw
nQTOrIa1JKSJsYb2/pqpF/e4FQJ2sbUwEQxat03nHPpansEcCbcKGIRNEkc5pjsDd0uhPHn4/O4T
UASaZ5brxUYIQnxAFO9MNVeDEjsYQrbCYtdxQMfa9bXIDh0oOKaA91UMcSSjIbypVP0yt7EiWChd
Z1H6vIwPg7y/WGZ1LEbgFmoufBNlJ3/t0zMt0b66zPmUXm3d0Suwky009s412RiLX1Xd79fr/elo
IDC9oqu6QU7wexdmuOdrYXinyPtV/wbouxWVf57UddaS/Ul/A8lQto4jr7PKBztI5kaN37cx+YUS
r0UNk7bXExNZ5Mjj5Z0FRpoIUvwmyabQzzsE8jYAdqPdYe1fcY47xYUjlBthptqVUbKoVHcu5qT5
phkZsw+R8Kzx3Yqp4u65BwxFgOPdTwWjj36dNM7wqgd+rR4OfqHTJSP61aOu9Pc1aPKGQvllBWbP
3xNwoWNzFIVxs5Qla4qIMUv2SWh0F7ag5J6A04BJzMCwTDWBwtx0S7WNCyuLQLOWZt4uSNSOQl/Q
FQi32UXw+7fAxw9mlpE7asea3r82DH0k+UsClcybQFBGyrJ8YA1/lIAWIf89WwPRm0X2EGZJDfaX
cczAwe/PGHMRUSgR9Pa6U+mLaRVZN1XqQK0gVeVjmsujxBoluNLzdQcKT2a6VHMBcPe0wZwwkI4j
XGYXY/g/XE2ThNzsqUkiCzWqNC66twQBgCbGCX2euZpdHGlalyPabtTG6Zkpq/+p3U/WPlzBykuP
CuTlsq8OxIQ6ZqzeNGnX+TiNWEba5Njj8pQscafP+mYeF5MmBlkPBzZ2vAM9bdXOiAJhlOmwGgg3
BcCFFSB0MsSJGpIZYMqK9qMBQE9Hn3tgZkcWWLwhIolZESlTr9pTocUYGyrb4Uh/MdwApvMWlJnC
36FHlE8ybECv4c3brpI7yntiDMMbvaNE2tl+B6wQXCi2SPH+WDSyeP2Cd7PNOCyxUiBgVPtlDdfr
vcOCxpWcqWHYAUbjjf8RMkFpZcz7nkfoCti7reK21dNEQvHdWWX4l/D9u+VbCyUjn2LeMjCw2GFN
u2700zWYfYCwvmrmsSblXdv7rAZ4vJpqxTS+h32cGD3FwgMSdR2ucyY0CtfjVMX7S0SyWVu6tAis
FtiSpgAm8PM9It5rO80f9JcAi5eMghNH+ue/rAqNrsO03LJ4MaZjbwIoXnQVT4CKj9aqeWMAxK6U
ts/2q+GY/CP4xps4I91+yARhF/2qFwAf4puyxc/vc4KLh9pgJ/ZkAlupM+eIQxPI9KEgAfI1zSPO
mbRCB5jPFqW0xwYMa6w9eYLOWjw7wesyLHyimLADussqhQiuV3hM/cPtqriwIJGXu3RAe0E7O9Vi
BbpPgYDRsgcjq4wIvd3+pFjKgFvyp488a2+Z5xf9pxIxAZ/xW5kR3iAhBa2o+OkjyfKRRqSdUKh5
6ePzCwLBSQteftj1LFzjI7AUhd87CqzzC/MxR6liihwE4C88TLInx4Wd1KBDTwDlYimwjQtK+ElF
CgG2bW3HJKBLsG2yu3h2iPI1Ku1OTEuD+1/C5BcuHrMdICP3svtrASNKGnLESlm9XLyiGczCOavs
iBy0EE0F4xKNj98hykzBscUVjcGmeox0pSZNO1mlDDJrNMP7Vb3FiP75ra2ZfFVHsRvT1TjCAfX6
QXPx8pZymsCGB2W6vmhZhb3A3gdoLbYxtoMYHacngtwoV+hBB2Z94Fedxgp4YvCaXrigBBZZ8TzY
wohxY85uPSjYUvEj4cRq7jWcE3AZltWtjbGMIVXZsUeHwcCrxvHYElemMfn7gCmirdxifpHKrER2
l3U1m68QRIfHmDsynjXn1i6kPRfjfXAlP+WxaPfPRA4/7r4oo83ylkZnF5FLJVnLypNBLL8h4F/u
v4Tz1Nx7mgd2MZgHDcIOHivQQZ9TlZ84URewudIiT5hTLg7BnJYDwEphfqlH2YSQ9qxzZYE9lfM4
m7QCpjBCNXJBQHUT2jlvYy4zw9sVeIeopqwAKFHPhWCx7I37AGVm3fSNSZy4MmKU+VbayIdlsXZw
Ob2bjvRdvosai9She7hKeHuJ/TWW9Nf5AQS+TrVQsPYLWScwo3i1KO1vP/iqx/QdFSQjVtFqYGnH
PpCO2l654Ygr1kbbYZPv1CQllXHRPHQPcfsHDp4uqzq3W5bOrYirwXgogRsKCEG0/I3vWkiDEqNv
BphiKJPchgh6MnNVKqYCOvJipWpyrQ2VSzYxTVCcasfEn3B6Hjg3e3m5if/GOSXZCO+k9AEVr8Yt
+Y/vH2VtAXMrtwMjwgsPmUcH/xJCBO9JtJv2NwjTyC2h1c7UrKy0Wy5O+CLIaj/FTJE8opy2OtJQ
n9yvMxNGnXYK21XfK7Jk8zhcO0xFNgogF5PhnGsRUfivGKWsWpz9lVayPKZ1EeVbz1hJ1NHY/7Zc
Ra1DPLoAzPayuTxrJBLBw0lw7P6e9N/ur5HsWcMf5hGut94z0t+buSiPpfZy8k8EbnaQCg+KeMTb
XK+3b7DCkcx5PYEkCs8NeqAWQ7XOavujNXuR5ygQeg7USfhCYkqM+aCdkNINZsoL8/oLZS5Upmhs
zaZy+J/wXoQrdtLdohEFlqznpxfjmsWxcA6Ne54IrSvHJ0E+Y6ujDt9w0Luh+wFrjkn/nu6l8526
gNTMEOj38qtRF2lcSKyb2wwZxEXlZLNoylWUoiwF6af3Yg2nxVprauBy5DhNmjnEcLfE7sbs+u64
cLanqjoSiSUzDLVLs1Fw+0Rz3ZY9giZOie0w2L5o1Ufq5WOY9G/c9vteVPtIcj1ZVIw1x3gPj31k
AVGS60eC+lu2OnJkyjEDOMyZ26y+Mbj2qakNyaZlD/OhC6h7XaumXYKl3Wt9HYYp6tBwCg3gSW9M
IZcmregUUkRN+wJm6nXllVCgBfionzj1BYOrnHnIK0rLL3UQSMrY3A4WKlSprUFt1j980f+f8DDq
6jGH60MchyHWinhe7sBdz/dJp0K11yrC9GQ18ALDS+LsLy5BNm/7xZmr/XswP6kAQuXaqmApjRPj
gvQgGJgKwx2/vC4/txMLNFypLMD6cNbe2WyltVO9FhkVVgibE5m9wisASzbW9sStVt369G6q3YkL
AKCNViU59uVYNHtAAi40S8uES6OZnzO82rgWEhJUkrqdE102V7B9gvv+/0zMdbEzjE9OFI1ixCDy
BhlPxmgHVt2+DsOj6qWQ3lq8d9gMSLVWv/HnbCYrzVOJXa3GNnoP0uT5hD+uFceQ0tIa2QDfozrF
+oa4UyQRqnBcWZHCEzQN6cB9RBH6hdQWQeWua67yMjY/jtG1t+Lhhsgw9WtypkfhPC6WpT7yN94F
Amo8EmpIzQlHNnAhOJqBDdVAdO4d5I+PEQ0Eaa1hvwRhk/2k9k3sPetHeJp6I3FUUyGKQBYMZ0PO
HhBOspI3caSKFdKeVzzPsHnHELkRTgSFM5pkkPrQgRAA7uL64I/rx+WOCBQDQWXekL/VGNnlMsN1
fE9m4ZS8veQo0X/EHWPTtzE3roZhm+2C1HiL2LGVT/MvGZ6gxoxwq7Rw2cu7ZowMklwcZTqiKEvZ
GZPBV5/B112zTRdvYXbi79Ru1JxaU5cAUym6J/R4q9xMgfMAXALJyAqU5KYjowO4pATdh9BE80WS
WcKocl+mn6AkxPRvgc7bkHcjQ4OG+T3p1EoQOm30ac5sBAFfmRd+lxL3g4i+G8zYQJSjjMJJzchV
K9n6K6PAqhlUfzJ/PDo+IEIGJ6bdPVqlyyrl8ZVIjww0fXcjO4TDQjCfnCPn1umkwFZ0aL8qJWqd
rmMOYZ5Y/TFHHeqWWhsXIxFOqKeSQHwgZ6IpJbi8ptK+BNaDYd2liD5LVPf/yZ6QZYC7mYJdBLqi
xXNsASaAp9wy3nwqA1QWzFShauRyVPRjRH5O34lK4mjU1VksvCQVUGus2Ef+9MY5HlSQrEWxcXFz
8YVkCT4s+NA3eLRW8SPwtNcKvpQPX5wVGpZH26i5eryEjYOZchLo74Q+o82Z5qLMU/zqcrYPHKzb
oqo/a4W2fTZ9RSl3au/rMA9vzt5nJep12bI4QG/L276lw1HARYZSBmrURT423Ezdojs1Bg7m+CMk
f4zsiZWhplsWPKTPGbzCN6wppBQGz+ualZHWc3voU3sXN0a/5HAyGWW47WIsZHZzDu/O5gC4yRQO
WjMhBEj8+UrlcLovaZMHIRg6gLPvY/rvGUtePkbH7ToYYq49aPuNja7jJ1T5H1irktutU60CxIKN
AUO6fZMxw+XxkwN5AQubkOUg8kRSYoxvvObKZKyix2jpFvon5pthjRi3bZfVUUJkyXSrZbYed+IH
ExQgMRH9Dm1gbC76VoxbjAxNUbQO4F5eh9RNZ9JiZr68vc+saOtCF3GCs5H1jrRt+36JIp9doK3a
tICiq6UzyZpQY0A8e8h1zjM1lpBqpBanDVcVgpOF9QjnO9QyRcaMkHUwSm7AJ3ZNSrzlzkFJCiYV
0sko6Nceh5ls5UbU+I0GjlYh0io8N7CzGQv45ayIZ1w5K1/C0yKtFSP2ur+w9Z3X4tve+RaDnxYR
U6Yh+bdYqtIifi7aIyms9s4EPyyTbj/G8xjlNvoay0eHk3vdMQWZ+yq+dFwrK2oFfMezLvFGjPDs
9nWf3SmQjBixcU8g0vKJollqn39XjLvmwGZQM5bAOESqfsxDdQsgEtWnWjOaZlNjELm6/WGFHnch
HZLOKtrxDWdGN7rW3JlJm2ABR+nWKNWJRygE/HGctoakVBngDhR5iraFzPxW6pbto462TpeJ+J5V
wRgGXQtVoi8vH93ggx0LZIMxlOId/MRAEKB6HgSru26WJx2gUMEuWh/lmoFkFs/A8lltpte6OLQw
uyrBB5s1Job2Flc58aHOE9MUfoenn9/qyRIzYAdwRiKBTFQR0KyY1bIFBAchl18uuhEq589Einxv
YEg4NidXbhGcHXgO/Ar1zKD6LRI9Yj2/2mLGJsQaMJ5Cf8jY77uo7rJNwhkVRWYK0+8ZIRxO5pfN
c2Vqb4l2rL9EwjJ/3Lk9Kd5JnKobLeXGEYduPZDMY60Js7YqiodbUK0QvtZ2sszQSRfZFWzYPQCS
QMkjoYJcnYtw/tUzjdevy0QKZFRoHSFm8f4qOJfPuR9314LqORLm+dr4kMw9XAhJUCFl6319B9CU
x3WlpHLh9n4hgoywEvND8cuNIb3EVTAhRkNqjHdneCrcTJVdwc+masTD6oiGuHrGKAGne79Lm15L
Zt/5YQslkkl2Xn19BMJBU7vt36FheKLY1JW7yZ6C44bYXbGOQckPKljpj0kKKS7tDV7JAsgp/6mj
fCTa7WqMQ3zKM50pFAx8BF/DtsTw/2SGQaYap735egGWGa+7WYMJ8Lm9gKv8KiJIFtcjFmGOOVIV
8l+v4kMFc1WdiJFJ/Aai71KmtwwxQora3nRKKTwbwPBwk471JkFVoZSTKaOHfXyRpSFY63rALF8n
4xON4U9h1YZpAdMEwXVqRnFn2qWPRKPxS96DGX1TCLfFQxNdlfuGRhUd2AfrNEnhIpsDyZ9r4nkH
tiDFlS1JZ9bGLWbcwrxFJ3v/Dy1mNw3dR8nFPBWEGjVufqRcMYRhQTiZc58wJbfy3ghQ44nshrHH
6xPqj1fgY/YRknBMFpJaKpB+toldwDefREAVVec9Bl7stka73OhukQqdeGJlW3GbLQa39EkynvQC
0m0eKcVfFxp1YzYe3MfJqyOZz+++5wB9CbXnPuhkiyFgzJA5xBmCG5XaplZhc6GPwFP3agWZhNUF
2E469FVmLZq1bTuSv4gRolUaFqx/BB2b9vjPW6y9cJc74OWSVkoRSx5cgN4REdLjV2BDRbPlo66k
lKrwLsTtkhdYkz1RD6mWGJBl4En935Xqb2nMqxOJ+pINXRGgjLnJHzmX1zstaow4HWjC2JkcrSKB
JsiNuztBKpACheZtkOqwMIIrLPtKXVgHOLUcpFe6lJBKBZU48iCZ/u4qBzkGrClS2o7i+/uXECAV
jKr15gzn3uh8sl6Ga0/oCQDaEsnzMzl9W4uwVyKLCv6aSYVi+//NXdVL4ka2W3mKv7/o2ffyeiKN
2f73RjGu0QQKafngI+TIjPbRNQyVjsRadAA3htgEbZb49T+QUYoO2ptkuas3p5ZGNZYo5YZh6Iho
vadcjMzJOE2LeJ0JgQznfTzGv4cXdxJH06AiJOqx5JqIQ32dBGV3tkgYZdvmUKDa7tRehzZ6KsMw
0fby+bOSdnIQJGqCS9mgW/k3MYdJWGQvGCDMZ8a6jjfLRnZV+7DGKRt0KaTNO9EtgF9HtL43cTo/
IO9Fk3UtWQG1y4TTSSj4exnRjmCkz3/8uwxrm+Zuc+Lwk1GirWlPb2cKd7At96RQoaiD0A0xJk9L
EeTX4FYvW4BEknUugt8+ktiT62P1i28UxdlVReUQF18FRva1GZYcHDjQ1w8PHl+AeMjsoS5wkjj7
VEn9c/fbljvnZAUpJRtH/rzgYf8rZGcFvFeraaQrE2z1IKvdcNfxpFY+azBmXXxKwJhmBmbeHfAK
vreP7Am9KvRtIgDgFrPyMEVMe++4MyARttEhFvWhOQ0Z7FoI1HTanuApL2mwfzNMy8/5xa2gcXnJ
o4XZO5sPdFaAi2epepxf6To4j12McVMMrKH0tvIZgkUSWPe4GuWzPIB1TALkbnK3afpfY+L8Ac4H
MwboUEjES943E21K7Soia1BRttYVesAkRyF+NxbJQ6hKSpf2BjODud++gEpB7AxRUCpoCfmBU1DM
FHpQzz6KnekuEjOuSDELWHBzk5bA0vgUHvmFKzXxwgHckc5Y0mgUvLluLLVjc7xM5mk7y/s8CvH/
xcE/rxZNfvQE9LQwHrFvXS8KHtqMpgZOaoweadNnfHdeOUtIfsbibzFX6FE6KoNcuwfulKXnRwvt
u92kcybMp/sv946yOhnjOh8+4KQesxkBHMWO28mohwGWpziyEabF9oPkj6RpJ7KZaxh/ljlaN8v4
d5xF8ye5G6p6ycKLAZAXeLfkw0TMCgSY+pRZSU7TPCrMQAq3L5n72QxbUPiCvRl09lY4m4xFZwIl
ZwV8Q9nWhmNSqUproBq5taoMBylNrr9REM/o/k5Cs8iY8R3PZh9xB9+vtZMcxlubCddgcxK8Qapz
hOJHMdiTCOV1HUIeC7gDf15Wfh9euD0S2e+1SmW41TlVqVqSCGRDGVuDvM/N9OvikLNPYY18+t17
Uzs8fZj9HOS5/faa050WAxApxwAMcikpBWx/qWefxI/3AvBJcr8VKehNPtHQh8lL0oA5/GFdRbHE
YXbX5SWeEFGQMCObz7wwsWbhd/lW0r1pUYaV1dQ5IjfxQxrSKzTLPnXJDYWWh3rz2sNBJiDF/azH
kAPXVlPqpoN0ekEyg7ayrQLVwpeP7bAgh9b7CH6HkRAh2gIAt+F2OJjO+Jqi5adCUYuPyNrONMaw
Ddt9yH2uX+oGhT+a3YMqkCu0sgDdtzcFFGpccYd3pV4ylwgxNiFqhcbFd/KVzGMk+k4Q+C1YjYPJ
qyxMwzowfv/bTEegBJkt99s5VXK7DWk0uTDoHeLxOx2LJhj+Eo3cu4hz8cjlN1ezX1U20rnYgwNg
mK6XXyQu/fL5K1omqlyBJxGlv9aS0CAPHi7F6H1ZTLhsDdzvPyaiolAJln4Iuih+9Z33+SWNQ8IZ
qazWh9O5/QdFjIeHfckRbmWqmQtDbs4vKZ/REJA+mfecCS5w1LyO2omCo15OEVGf62nMoFSiF1aW
RgmfXUZcGYpip98bQX5LJ/nexjFTFuarfjjqcuvM7H5BTmP6Rcb0BbIZT34X9WVLZfvq4MYUu6dg
Url+NzZl41cCB9xeU3hyDoVyibrnMH3hMLohjuNdF5ioJGC0VnOmvL66pX5HgvPTpzHpauxpg6z4
87GUuSxNTdALfRngLTMvLnLhQuW5ld8TBflWNoS2nIcS64p0kSsxZQ6uOiFIrPsjQlmuDbB+/40W
1taullT+CfZYEqjuz9D+3wR51Y92tnkXWcelKRDiaIbB26Rb6qVa2J6YQuhQHt4WUXZZEOfFl3Ax
6cVnqtXzzmLzFfhQsTWR2xK30/NH0oejMSnlZs7UubCa4LrlGWja4uOfPsy2XPoPFiEHIbkK0jTC
YlQCo3kYBFo7uxWVg6WoxgJaUNaLwc7yduhF1HhdBUpUp2/vzDv4ckRpgypFIOhO7V1kQPVANR4+
/yIH+8VBFRxQ3WZUUICDu6nuHUbjS1Al37x+n6NCLBg45p9687p+nQNvpZMHXvzlCaqzAJTm0uj6
dWCq6efpt6hW9dKsxGaYJeN0GgK03DdUl8pUAxrxlbqNRr7j+kUEvg335U1i0NHMgmBOMuD4wjpt
QPMTX4QYoDB4TLlmpcaJOmYMEfcCUHeOgrolhv18DK7sIZ2lIHDBqnON9/lboG5mlHKuRDm1HFGT
lzKxjdbCBsHM/HRWfnVahm5zv6AyTLIjNFWsSS8wUnBBulwthPLAD5Jb6Na5w0eATptKPri+ZUtZ
Vjuh/RQ35yvVReQ/zN6bMych1uLMS1qj5r4zaUa3pdECyetwZ401oafsD+8rnHOyM04dXXumOUIx
PtUkit/0YVm95r/wHX9HjL4bmj7d3SzvZugHjUZuzVGtaZ6e5JKuze0a6QbBawDYNq2C2BVa+Hgb
nNCh1kZgo2oJB4NOMC/DSF8lnY/4eP9+mi2utRQpjeDxyoKbZp/9plgAHYm8erKW8VGOyH5PAHpN
v916jN9+2PlF/YGPnv67Jll8ofG8fUXUb9E/01wJIdxFBMkRVVpCpsw8dKpUdHezAKiY4yyEqGEU
bN5y5kbcez0Xjl6XiQfsnRRpnCYUKhKmQJB2cLvBuBYoD+6W0lSA7tEvCw5Iyw2vHj1e0JAj73as
TvsJqEWpKI2LfMq3/IAh8UupHkH580X8Qu7ZNREnqCutqcvY+e7No/Pm03FdPJKDbZOJb+Cmx3a7
l8ki+nTBFQeY24Wu0bf77BklA7wUXyYLJHG0xKZ4iy1KyWcsKv1gNNUvwreE/5BID/TIH0VrhIFZ
LeSOcN5pwPfXvdinY00VPjrPpWspCDSoPveoqahFzGViqD4gP641+/H4bBz4nUPy6v5KeVY0wXsk
QJeNNV3uV36Mj+wK6yEbDw7t5IO956zaHPEw5bPY2TiYoPLCx0oonp0Cmqih7QW8UYLnZte6UZKa
Ag4uc/BZemz+tzZttMocnRbtQVVyhuzSgudhRYqzplXiIitY+D2qlAflUdxmXOuhdB8yb+9j4sl4
OIS4N4HwRplhxXjciJQSaCz0DWWrlQcQ2PduXJXG4HJF4CIKlP71F9rPB55kFukipRnoG31M2eLe
TlKj4U16IJqcjVsgO0sMwVkbJN6CTKUQ072/JoliEGrv8HiEOaxIcckiy1VBYKHjJMg/r9HjHuby
rkKic4t3A+jFBrhD6VDQHTaNpPJmvz31dACBh3hZh4mEDSBods7Mr/peNaO9Z10zoStbrARZNec0
SyNHCJP+mODt/sm4pyjBOQ86nsP3XFFEJiF6yFnCplJBTMen50X8YASUdw2ZkidEUFEMzhTEfNBv
A+1ZRfbKmaT7eDrLBULS3GK1ADgKg7mYRZGgEIjT0HGL0eqgKXQeA6NIzxeC5G+RR32IG8GLc8s5
2/l2yI32Ah5+dyeEOPCwmOJ5UAV7AVl1fjIKsH6FZ1vSJe7N872hoNBWG/x75ioTnV+k3EZWEQXz
xe10gZvZZoYgpYRH5iFGR84JdmGjSoyfXb+NfL0vq41l6yVY0DQMD2G1ba4kLhtjaQgatglcS98b
R3Z4HRHEr6DlUTv65j93g+E4SXdrlXZPse3MLpbjdGt2m5JQfxhfsnNBg8aoJJhgCV/Uq8UVQvJT
l8mxwxgBqbANOVY9eNr6KliEqO4I8i8hLrwQWw6ubJDf5BbgqqMJY1cQrfmn69BNqV7Dw9o0V5Ky
VHi+GZC/mn9qqSSWbDjy6cFG7ec+Y/L5hYEAgULu1DBi1FJhdz8QjyWaCGvpy6BHUfmfcIroF9hL
ajcMNAY+XsyPZYUo8stofVhvJfoalxc7NpIFutpHkePJp4WMExqQJXIVfg/PNz4SuotTQXdqr1K+
7X86r/b4yOq3dkv411g3rHVL1UeF7qdduuA6mxO7IGoljGnYYGWgXyNV5C6f9myJ+Ua1qNrsXUqx
nVJIggaocVfhYMccf0u4Z3EZST2eDtQnT5TvoNKl3xkIUO3MtpuYI3bqqpFiX7rKKDMLocYhs6+9
A42P0Yw8OVpTRU2j4+PtJgO24ym7nnOwjr4I1gI1KwJ20fEVbs5VFFlSTEprIihg2O1GQRmOVbMQ
MMomH1STw3SQEmNbS1CA4MXJDZrnwKHDKRY7+8FDrF7VSwva4/LOd6yi1EctRohZPd9EeiaSKUnk
AoI/9cKTqSi6jI93bwgyvP4A/bAWdw+Sbdlr9nZiMCYIHrxVF0pp2COLTPCm1kxcLtQXRrydykCK
y/+CMBo0HMsDK0A/xrcXnjW6OYZnRd5dM1zqxAMweQ0nVMyIPMqC7yWwtLqagTQ2ji52QeYE7gFR
mHPNsqjck7qUndAfGfUBmVlg7J7pG2XvKvs6JltgZE6Bh4G/36kgl7a7qLN9O1XNcJy6NkYOt9Hc
VvKACHnIFy4qRliyayBjv67H0HOApIibFYehjN+xuvlWtmHABtRSrZipp3KWi9qcfE0761AUwslV
5IQ+YPehqLRxoL1GtIketq0kx0nX2mhCIrhibELtxwaUYRkfae0M0zc38ZnItqsmcRYwOVsHTSGn
4F2tJaU46qqqphWHU6ytH4zLurQW6K+AFC1+tGpvHPj2vN/PL3SXpBpnuGH+VqYXDfFJm1jW2gPY
SaGOPCCJf5BGx35Df7Pkq1Svt/0wivzDai5VL6xB5Z1D7CisXdrFodbqBQtXtnMKLxkA7E1r25Qq
HEhQKjvyI2rno2KrnAhImGyQfuQG2Cxynfz5SYIIdPtOnydcKL7aDppOQl6GLRMIBB5VHHffJYaj
vddOSBAYUYgKtttTngTFGSbzSgTEB0dsXgFgo1MXA3Ono3xSo5DF6XrxXt7Dj7q5YUtJ486dlX9/
hmx3NJiRS5lqW1JmEDLT7ejlUQ9QKzbbspfbnHohboOEGT2PijLgw1tZ0hSTTz0jbBUWKOJB4r9m
ZXTd124Y9yIanmQP/fDliRNZniGVEodhTt+6hCUE7lG9nntsqPZueBlqQ8G9p/bhdVuDRdcuiSST
Nb7kPaiw9yuJKs1xO60AeHSRPOgFxyKXB7XHJaSFIpRmIjFfBrvISaT183+pTwpft7gYt7LcGx8e
sWFTnHitY4oRJvTLGt+PHTdYpQbQS6IMuDebUFZoCutBuhunv+vTV5rU3R66njFS3nAU+cIb8HU0
DGDG9mR1GTZlC/KW3QbQLbJgmBfAIIGwiCo+2A99DHHFt2DDltLHNKt45EohiCjhHIPjc30tZZgT
APGEtolC6ZHkJWFC+3lpjOTqBLvfEgfCsHJTb6btW01gS08rE8x+IXClyEMP6XtYmt5RV3WXbB3b
bSoayZjMqpR7AAC24TQC4uBbqChOXAj7B5idvCIuMcM1SwNJ5PPgJVwxv7IRL3xcoIEvJ+E0qA3E
ijk9w/FobMqAanOqGy3ifO5BpJZp720iqQDvV/pjmhxOzzJC6+qQUIkhbe9IGeL+jRU2PukIiBpa
xvT1z3RozLwDv/HP0xk38Ps1XbVhnc68SumEkYvL0rmzK/DveUvzkIvcoUgvoT/4K3SegCeWJcp9
SioMkxHG5plQdAJXDbZfCr5oVZBxA5uuePkXr41/BcLHYGCA0wLRFNQRXRQIHr4eDhx32Jqa8rWb
C0nqYyOrziR+BKRfBg6hrNLzlw7pK1OrtsEWMa8v8aMZ94YOqzFEysHh9pjrLqLAGSWUocT7dW8Q
XSbZEf05pHuyM/UNda7Yv1mDZVGtzKVKwGj6KF+gqitBoxCjy76uIgme/WoMVBzOupo/ZU/EwLF2
xGvpRZ/sPL2sqIeWe6VgtgvOVKuqFfXGTYzFFBkoY7yaij/iBAiEM7RRAuPIj8Iadjxz1g5U6i8c
OVD9wIUBoUbAStxIiNOf7m2NU2PApxoBErKgchS2P3y+LAcw7DiPf8bSMcq4OJgXWh1k0mhu6mZE
5J49qfll0Vs9WJj9tIpLWaFUgbZ3Q8LT4cjLhn5ppOMfQMVCRLIHScHD5ieRzMLo/jnPyDYx80PD
R6AOVMKRObedvsqwdP1xVRb4IZZMGqrmEMEfqVHfpXCkMIsDzu+hMxGHj7d8ZJrcIlOeTDc5QW/1
jYPFZeCKkTlhCLrd/9JMtviO6FtMl+bxawVeoi7+EKDSh9CHIvGbgX+iw96VFybudkmsIKMDG6Je
0bNEfJ/o//2DdgQYmP55WcEoCRO5uqG5MaI+EQJrONjkorwwI3G8FktlYZwAaouLeLPm39B4aU4g
mJA2hq0HQpNyBUbjubIOQiV181EL5mUQq4iQcLNjWROJ/GlZNlagSsIL+Eot5/h60qoE0l3+KsFB
sf9IGL/x+AC0OsMyardk42wjpdZrf/5+fv7J5ScU4ycRkDDaANXNIw/GWtUc/WqkWlxFZRzziHSx
YxuUpCARqn0EtILxNAdi0Rveh4fV+xRd2yzMdyn9D56MKK1z2FiHmGzoQBZt1fknKRyuoX+cvVVM
OnIYtu2/Bgjn1Z+SgcMwB111mnlvbKq+gs29qPDnO7n2v800ve8MbivkQXQMLICOf4/sJz27t0iu
VlxTMNr2IS0F8wGASy59iZpprCi3VbqQhbsd+T9ZNrEBKg3shfeNZYFhXmVSxRlwRCWipZxUceus
qXKPUmB6wik86cku9vx9Rlo6bLC5fyW5WS8FubnWc7pPVedK7O/ZcHlycSjfeW8djJrApffYjPBF
GqEWGUCaMDR+jwaVWKaXbiXbWUdRCvpgDF0YoMMoh+ac4W/EvRHz4jD6AsXI2iXIcWJ4M7wmIRF8
8Oga0P24MzNpJLNS+G7sM42GM2ZKMWGez4fJayV+4iRU/oOCFiVnVUCkkDrez+92W9SHPdKyPCij
u7CVu9clXq8ynxl6u48OCNeZWQ0xGUMQOLmcIDrL+E88jchchlDJEIerkWwpBSg9B0gFQc+jhjru
3t1XgAOXt6ipwySDBRtqDUqJ9UTVi+5jHJqMNfaA6bdZJ5zWWLtXtEe/XTamsKTECneOHi1yzyNe
I33mxXm2LRivKFmDkqCEFCmt7LS2C4x/zAih6kOVM5C1ebviqhf9auJPw4JoT/c1KWXsnIQuXnGY
raMuN7OYxXVI8CK50LRI00uwtCI6E4oNuT+YtkR6Ptyer9khCYqu4wgjkIbqLF1/j1LfT4KVfnJg
tJKe3nU3elIMQmb3+XoY5uS1hE0Akzc0iTjxwzah4T2y6UvbIKQ+6LPpwwGlseaMP/Y502FEvzeO
1J2FCX3lgQu4phatxVoXiXVuMlZocVLuEj31IA5Q/tDejiydS3/LIPzIQrmYgZXN4rPIQa7ykPjc
/QhEaZKAVbjHCF15O8jzAybkU2Pv7Sbtg5X04CWn5hd+VxVe9sLzWTjjPthAZIfDqTRfXcLOOndC
a6XwhAGVMttpoC96G4nLsVLDB1THwPl+hzRqxTRSSgY1vCpaGNXD/5xKwxzYB8LGtphZSwUGlA87
/MM1aZfDR9HbwrL4cTRvOB03r2WPY1wAhYAwPJJSWVxBXTWKBSqos8qwJzUoyHGVL98oJ/vmsfjV
kpGrsL6narXfTD2RWZX9eW7KVdl0OfQ3pn0e07pFXj17L/j1HxomkVu7q/gZj32qNQUlJg/FQoKr
UlFf7iHFDC8uN2acqdpz9F45+eHMoikLbekwz4KCe10ztdv7Yq924kbdofONQ2aA3aM/0SIn5m0c
aepIAiSXCKlzb22RhM6Ic7Egnp7CdVmw5dFTN6MDnvFghnej6YSBELiqSdYGCypE/uICbiE16ixA
KR/Ox++2Zl/YouN3oK6BmyTrSWjImeAcljjLoMx4HpZ0WB/PCIDiQWzsoEPJta9NvMRpx3+bBon0
X3lENdO0Rz/yopMBc7ih6KAAWKMyksSZK7B7Pq3G9yDsCUvZ3QvMNg9lemelVXk5qqsOo9/YHP/u
Y57C/joosAHkCEpKHTkU383l3Q25Jgrh+jrV40miMbNhONEznqdCHviPk/3R9VSgqhMD3wjmDpuJ
dzd93y+BUC3pkEKFJSNXUU/rSngEu4NOVLkaVErTMjcHXalSvfoVl3KjunvW2dkyv6DQa9f6gpAk
Hd6i3okjJvqW5/w+q5fbT6NWAY1oM/s0pGil9I1VPzghgucAOVCJcpoJhrH81P+vnGHQ9al5IeVR
k+H+ppFWQDYHzuUWv9DyJu0eoTedinCsBh+m+o4kMsBIhG6BOWQ7OWrHv+F2hi0+Gc9fNRlKo5Qx
fdgQPBfKcRfjGPcfqbQ53487Lvjfogy+yHBoheV7//uCuHS6KVoVGWb+qBqiqDlPr/x0vXQXw+bc
TDQ1okeHH2/ifaol1AqKpnYWTqoW0ebP9xDqRt6hwPiFytiL3h6imP0EpvmlO/flc22h30pNk4Qt
qeNUjfmESeg4TpG5dK7aL3fMQBZSPdcj72IzI39X2h/8x8FSu+wEve4LMA5kjBabkuE8SY2Ok0dQ
1QkHSqcYynzl/V8YIDSmhw8HoFQ168IW8IO2Ja0+dnb0rj5ezQZz2yOu2V9jsWTQu5pSZGNBDCuw
`pragma protect end_protected

// 
